
module IF_DEC_regFile ( clk, rst_n, flush, stallcache, stall_lw_use, 
        instruction_next, PCplus4, branchOffset, opcode, Rs, Rt, Rd, shamt, 
        funct, immediate, instruction_regI, PCplus4_regI );
  input [31:0] instruction_next;
  input [31:0] PCplus4;
  output [15:0] branchOffset;
  output [5:0] opcode;
  output [4:0] Rs;
  output [4:0] Rt;
  output [4:0] Rd;
  output [4:0] shamt;
  output [5:0] funct;
  output [15:0] immediate;
  output [31:0] instruction_regI;
  output [31:0] PCplus4_regI;
  input clk, rst_n, flush, stallcache, stall_lw_use;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n1, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148;

  DFFRX1 \PCplus4_regI_reg[31]  ( .D(n66), .CK(clk), .RN(n144), .Q(
        PCplus4_regI[31]) );
  DFFRX1 \PCplus4_regI_reg[30]  ( .D(n65), .CK(clk), .RN(n144), .Q(
        PCplus4_regI[30]) );
  DFFRX1 \PCplus4_regI_reg[29]  ( .D(n64), .CK(clk), .RN(n144), .Q(
        PCplus4_regI[29]) );
  DFFRX1 \PCplus4_regI_reg[28]  ( .D(n63), .CK(clk), .RN(n144), .Q(
        PCplus4_regI[28]) );
  DFFRX1 \PCplus4_regI_reg[27]  ( .D(n62), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[27]) );
  DFFRX1 \PCplus4_regI_reg[26]  ( .D(n61), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[26]) );
  DFFRX1 \PCplus4_regI_reg[25]  ( .D(n60), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[25]) );
  DFFRX1 \PCplus4_regI_reg[24]  ( .D(n59), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[24]) );
  DFFRX1 \PCplus4_regI_reg[23]  ( .D(n58), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[23]) );
  DFFRX1 \PCplus4_regI_reg[22]  ( .D(n57), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[22]) );
  DFFRX1 \PCplus4_regI_reg[21]  ( .D(n56), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[21]) );
  DFFRX1 \PCplus4_regI_reg[20]  ( .D(n55), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[20]) );
  DFFRX1 \PCplus4_regI_reg[19]  ( .D(n54), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[19]) );
  DFFRX1 \PCplus4_regI_reg[18]  ( .D(n53), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[18]) );
  DFFRX1 \PCplus4_regI_reg[17]  ( .D(n52), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[17]) );
  DFFRX1 \PCplus4_regI_reg[16]  ( .D(n51), .CK(clk), .RN(n143), .Q(
        PCplus4_regI[16]) );
  DFFRX1 \PCplus4_regI_reg[15]  ( .D(n50), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[15]) );
  DFFRX1 \PCplus4_regI_reg[14]  ( .D(n49), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[14]) );
  DFFRX1 \PCplus4_regI_reg[13]  ( .D(n48), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[13]) );
  DFFRX1 \PCplus4_regI_reg[12]  ( .D(n47), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[12]) );
  DFFRX1 \PCplus4_regI_reg[11]  ( .D(n46), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[11]) );
  DFFRX1 \PCplus4_regI_reg[10]  ( .D(n45), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[10]) );
  DFFRX1 \PCplus4_regI_reg[9]  ( .D(n44), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[9]) );
  DFFRX1 \PCplus4_regI_reg[8]  ( .D(n43), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[8]) );
  DFFRX1 \PCplus4_regI_reg[7]  ( .D(n42), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[7]) );
  DFFRX1 \PCplus4_regI_reg[6]  ( .D(n41), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[6]) );
  DFFRX1 \PCplus4_regI_reg[5]  ( .D(n40), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[5]) );
  DFFRX1 \PCplus4_regI_reg[4]  ( .D(n39), .CK(clk), .RN(n142), .Q(
        PCplus4_regI[4]) );
  DFFRX1 \PCplus4_regI_reg[3]  ( .D(n38), .CK(clk), .RN(n141), .Q(
        PCplus4_regI[3]) );
  DFFRX1 \PCplus4_regI_reg[2]  ( .D(n37), .CK(clk), .RN(n141), .Q(
        PCplus4_regI[2]) );
  DFFRX1 \PCplus4_regI_reg[1]  ( .D(n36), .CK(clk), .RN(n141), .Q(
        PCplus4_regI[1]) );
  DFFRX1 \PCplus4_regI_reg[0]  ( .D(n35), .CK(clk), .RN(n141), .Q(
        PCplus4_regI[0]) );
  DFFRX2 \instruction_regI_reg[3]  ( .D(n6), .CK(clk), .RN(n139), .Q(funct[3])
         );
  DFFRX2 \instruction_regI_reg[1]  ( .D(n4), .CK(clk), .RN(n139), .Q(funct[1])
         );
  DFFRX2 \instruction_regI_reg[26]  ( .D(n29), .CK(clk), .RN(n141), .Q(
        opcode[0]) );
  DFFRX1 \instruction_regI_reg[25]  ( .D(n28), .CK(clk), .RN(n141), .Q(Rs[4])
         );
  DFFRX1 \instruction_regI_reg[24]  ( .D(n27), .CK(clk), .RN(n141), .Q(Rs[3])
         );
  DFFRX1 \instruction_regI_reg[23]  ( .D(n26), .CK(clk), .RN(n140), .Q(Rs[2])
         );
  DFFRX1 \instruction_regI_reg[22]  ( .D(n25), .CK(clk), .RN(n140), .Q(Rs[1])
         );
  DFFRX1 \instruction_regI_reg[21]  ( .D(n24), .CK(clk), .RN(n140), .Q(Rs[0])
         );
  DFFRX1 \instruction_regI_reg[20]  ( .D(n23), .CK(clk), .RN(n140), .Q(Rt[4])
         );
  DFFRX1 \instruction_regI_reg[19]  ( .D(n22), .CK(clk), .RN(n140), .Q(Rt[3])
         );
  DFFRX1 \instruction_regI_reg[18]  ( .D(n21), .CK(clk), .RN(n140), .Q(Rt[2])
         );
  DFFRX1 \instruction_regI_reg[17]  ( .D(n20), .CK(clk), .RN(n140), .Q(Rt[1])
         );
  DFFRX1 \instruction_regI_reg[16]  ( .D(n19), .CK(clk), .RN(n140), .Q(Rt[0])
         );
  DFFRX1 \instruction_regI_reg[30]  ( .D(n33), .CK(clk), .RN(n141), .Q(
        opcode[4]) );
  DFFRX1 \instruction_regI_reg[31]  ( .D(n34), .CK(clk), .RN(n141), .Q(
        opcode[5]) );
  DFFRX2 \instruction_regI_reg[29]  ( .D(n32), .CK(clk), .RN(n141), .Q(
        opcode[3]) );
  DFFRX2 \instruction_regI_reg[28]  ( .D(n31), .CK(clk), .RN(n141), .Q(
        opcode[2]) );
  DFFRX2 \instruction_regI_reg[27]  ( .D(n30), .CK(clk), .RN(n141), .Q(
        opcode[1]) );
  DFFRX1 \instruction_regI_reg[2]  ( .D(n5), .CK(clk), .RN(n139), .Q(funct[2])
         );
  DFFRX1 \instruction_regI_reg[4]  ( .D(n7), .CK(clk), .RN(n139), .Q(funct[4])
         );
  DFFRX1 \instruction_regI_reg[5]  ( .D(n8), .CK(clk), .RN(n139), .Q(funct[5])
         );
  DFFRX1 \instruction_regI_reg[6]  ( .D(n9), .CK(clk), .RN(n139), .Q(shamt[0])
         );
  DFFRX1 \instruction_regI_reg[7]  ( .D(n10), .CK(clk), .RN(n139), .Q(shamt[1]) );
  DFFRX1 \instruction_regI_reg[8]  ( .D(n11), .CK(clk), .RN(n139), .Q(shamt[2]) );
  DFFRX1 \instruction_regI_reg[9]  ( .D(n12), .CK(clk), .RN(n139), .Q(shamt[3]) );
  DFFRX1 \instruction_regI_reg[10]  ( .D(n13), .CK(clk), .RN(n139), .Q(
        shamt[4]) );
  DFFRX1 \instruction_regI_reg[11]  ( .D(n14), .CK(clk), .RN(n139), .Q(Rd[0])
         );
  DFFRX1 \instruction_regI_reg[12]  ( .D(n15), .CK(clk), .RN(n140), .Q(Rd[1])
         );
  DFFRX1 \instruction_regI_reg[13]  ( .D(n16), .CK(clk), .RN(n140), .Q(Rd[2])
         );
  DFFRX1 \instruction_regI_reg[14]  ( .D(n17), .CK(clk), .RN(n140), .Q(Rd[3])
         );
  DFFRX1 \instruction_regI_reg[15]  ( .D(n18), .CK(clk), .RN(n140), .Q(Rd[4])
         );
  DFFRX1 \instruction_regI_reg[0]  ( .D(n3), .CK(clk), .RN(n139), .Q(funct[0])
         );
  CLKINVX4 U2 ( .A(flush), .Y(n146) );
  CLKAND2X2 U3 ( .A(n147), .B(n146), .Y(n1) );
  INVX4 U4 ( .A(n147), .Y(n148) );
  CLKBUFX3 U5 ( .A(n133), .Y(n137) );
  CLKBUFX3 U6 ( .A(n1), .Y(n130) );
  CLKBUFX3 U7 ( .A(opcode[5]), .Y(instruction_regI[31]) );
  CLKBUFX3 U8 ( .A(funct[3]), .Y(instruction_regI[3]) );
  CLKBUFX2 U9 ( .A(Rt[0]), .Y(instruction_regI[16]) );
  CLKBUFX2 U10 ( .A(Rt[1]), .Y(instruction_regI[17]) );
  CLKBUFX2 U11 ( .A(Rt[2]), .Y(instruction_regI[18]) );
  CLKBUFX2 U12 ( .A(Rt[3]), .Y(instruction_regI[19]) );
  CLKBUFX2 U13 ( .A(Rt[4]), .Y(instruction_regI[20]) );
  CLKBUFX2 U14 ( .A(Rs[0]), .Y(instruction_regI[21]) );
  CLKBUFX2 U15 ( .A(Rs[1]), .Y(instruction_regI[22]) );
  CLKBUFX2 U16 ( .A(Rs[2]), .Y(instruction_regI[23]) );
  CLKBUFX2 U17 ( .A(Rs[3]), .Y(instruction_regI[24]) );
  CLKBUFX2 U18 ( .A(Rs[4]), .Y(instruction_regI[25]) );
  CLKBUFX3 U19 ( .A(opcode[4]), .Y(instruction_regI[30]) );
  CLKBUFX3 U20 ( .A(opcode[0]), .Y(instruction_regI[26]) );
  CLKBUFX3 U21 ( .A(funct[1]), .Y(instruction_regI[1]) );
  CLKBUFX3 U22 ( .A(funct[4]), .Y(instruction_regI[4]) );
  CLKBUFX3 U23 ( .A(funct[2]), .Y(instruction_regI[2]) );
  CLKBUFX3 U24 ( .A(funct[5]), .Y(instruction_regI[5]) );
  CLKBUFX3 U25 ( .A(funct[0]), .Y(instruction_regI[0]) );
  CLKBUFX3 U26 ( .A(shamt[4]), .Y(instruction_regI[10]) );
  CLKBUFX3 U27 ( .A(Rd[0]), .Y(instruction_regI[11]) );
  CLKBUFX3 U28 ( .A(Rd[1]), .Y(instruction_regI[12]) );
  CLKBUFX3 U29 ( .A(Rd[2]), .Y(instruction_regI[13]) );
  CLKBUFX3 U30 ( .A(Rd[3]), .Y(instruction_regI[14]) );
  CLKBUFX3 U31 ( .A(Rd[4]), .Y(instruction_regI[15]) );
  CLKBUFX3 U32 ( .A(shamt[0]), .Y(instruction_regI[6]) );
  CLKBUFX3 U33 ( .A(shamt[1]), .Y(instruction_regI[7]) );
  CLKBUFX3 U34 ( .A(shamt[2]), .Y(instruction_regI[8]) );
  CLKBUFX3 U35 ( .A(shamt[3]), .Y(instruction_regI[9]) );
  CLKBUFX3 U36 ( .A(opcode[3]), .Y(instruction_regI[29]) );
  CLKBUFX3 U37 ( .A(opcode[2]), .Y(instruction_regI[28]) );
  CLKBUFX3 U38 ( .A(opcode[1]), .Y(instruction_regI[27]) );
  AO22X1 U39 ( .A0(PCplus4_regI[30]), .A1(n133), .B0(PCplus4[30]), .B1(n1), 
        .Y(n65) );
  AO22X1 U40 ( .A0(PCplus4_regI[29]), .A1(n133), .B0(PCplus4[29]), .B1(n1), 
        .Y(n64) );
  AO22X1 U41 ( .A0(PCplus4_regI[28]), .A1(n133), .B0(PCplus4[28]), .B1(n1), 
        .Y(n63) );
  AO22X1 U42 ( .A0(PCplus4_regI[27]), .A1(n137), .B0(PCplus4[27]), .B1(n1), 
        .Y(n62) );
  BUFX2 U43 ( .A(n148), .Y(n134) );
  CLKBUFX2 U44 ( .A(rst_n), .Y(n138) );
  CLKBUFX3 U45 ( .A(n148), .Y(n135) );
  CLKBUFX3 U46 ( .A(n148), .Y(n136) );
  CLKBUFX3 U47 ( .A(n1), .Y(n131) );
  CLKBUFX3 U48 ( .A(n1), .Y(n132) );
  CLKBUFX3 U49 ( .A(n138), .Y(n141) );
  CLKBUFX3 U50 ( .A(n145), .Y(n142) );
  CLKBUFX3 U51 ( .A(n138), .Y(n143) );
  CLKBUFX3 U52 ( .A(n145), .Y(n140) );
  CLKBUFX3 U53 ( .A(n145), .Y(n139) );
  CLKBUFX3 U54 ( .A(n138), .Y(n144) );
  CLKBUFX3 U55 ( .A(n148), .Y(n133) );
  CLKBUFX3 U56 ( .A(n138), .Y(n145) );
  OAI21XL U57 ( .A0(stall_lw_use), .A1(stallcache), .B0(n146), .Y(n147) );
  AO22X1 U58 ( .A0(opcode[1]), .A1(n133), .B0(instruction_next[27]), .B1(n131), 
        .Y(n30) );
  AO22X1 U59 ( .A0(opcode[3]), .A1(n135), .B0(instruction_next[29]), .B1(n132), 
        .Y(n32) );
  AO22X1 U60 ( .A0(funct[4]), .A1(n135), .B0(instruction_next[4]), .B1(n131), 
        .Y(n7) );
  AO22X1 U61 ( .A0(funct[2]), .A1(n135), .B0(instruction_next[2]), .B1(n131), 
        .Y(n5) );
  AO22X1 U62 ( .A0(funct[5]), .A1(n135), .B0(instruction_next[5]), .B1(n131), 
        .Y(n8) );
  AO22X1 U63 ( .A0(funct[1]), .A1(n134), .B0(instruction_next[1]), .B1(n130), 
        .Y(n4) );
  AO22X1 U64 ( .A0(PCplus4_regI[4]), .A1(n136), .B0(PCplus4[4]), .B1(n132), 
        .Y(n39) );
  AO22X1 U65 ( .A0(funct[3]), .A1(n135), .B0(instruction_next[3]), .B1(n131), 
        .Y(n6) );
  AO22X1 U66 ( .A0(shamt[4]), .A1(n135), .B0(instruction_next[10]), .B1(n131), 
        .Y(n13) );
  AO22X1 U67 ( .A0(funct[0]), .A1(n134), .B0(instruction_next[0]), .B1(n130), 
        .Y(n3) );
  AO22X1 U68 ( .A0(opcode[0]), .A1(n135), .B0(instruction_next[26]), .B1(n132), 
        .Y(n29) );
  AO22X1 U69 ( .A0(opcode[4]), .A1(n133), .B0(instruction_next[30]), .B1(n131), 
        .Y(n33) );
  AO22X1 U70 ( .A0(Rt[0]), .A1(n134), .B0(instruction_next[16]), .B1(n130), 
        .Y(n19) );
  AO22X1 U71 ( .A0(Rt[1]), .A1(n134), .B0(instruction_next[17]), .B1(n130), 
        .Y(n20) );
  AO22X1 U72 ( .A0(Rt[2]), .A1(n134), .B0(instruction_next[18]), .B1(n130), 
        .Y(n21) );
  AO22X1 U73 ( .A0(Rt[3]), .A1(n134), .B0(instruction_next[19]), .B1(n130), 
        .Y(n22) );
  AO22X1 U74 ( .A0(Rt[4]), .A1(n134), .B0(instruction_next[20]), .B1(n130), 
        .Y(n23) );
  AO22X1 U75 ( .A0(Rs[0]), .A1(n134), .B0(instruction_next[21]), .B1(n130), 
        .Y(n24) );
  AO22X1 U76 ( .A0(Rs[1]), .A1(n134), .B0(instruction_next[22]), .B1(n130), 
        .Y(n25) );
  AO22X1 U77 ( .A0(Rs[2]), .A1(n134), .B0(instruction_next[23]), .B1(n130), 
        .Y(n26) );
  AO22X1 U78 ( .A0(Rs[3]), .A1(n134), .B0(instruction_next[24]), .B1(n130), 
        .Y(n27) );
  AO22X1 U79 ( .A0(Rs[4]), .A1(n134), .B0(instruction_next[25]), .B1(n130), 
        .Y(n28) );
  AO22X1 U80 ( .A0(Rd[4]), .A1(n135), .B0(instruction_next[15]), .B1(n131), 
        .Y(n18) );
  AO22X1 U81 ( .A0(Rd[3]), .A1(n135), .B0(instruction_next[14]), .B1(n1), .Y(
        n17) );
  AO22X1 U82 ( .A0(Rd[2]), .A1(n135), .B0(instruction_next[13]), .B1(n131), 
        .Y(n16) );
  AO22X1 U83 ( .A0(Rd[1]), .A1(n135), .B0(instruction_next[12]), .B1(n131), 
        .Y(n15) );
  AO22X1 U84 ( .A0(Rd[0]), .A1(n135), .B0(instruction_next[11]), .B1(n131), 
        .Y(n14) );
  AO22X1 U85 ( .A0(shamt[3]), .A1(n135), .B0(instruction_next[9]), .B1(n131), 
        .Y(n12) );
  AO22X1 U86 ( .A0(shamt[2]), .A1(n135), .B0(instruction_next[8]), .B1(n131), 
        .Y(n11) );
  AO22X1 U87 ( .A0(shamt[0]), .A1(n135), .B0(instruction_next[6]), .B1(n131), 
        .Y(n9) );
  AO22X1 U88 ( .A0(shamt[1]), .A1(n135), .B0(instruction_next[7]), .B1(n131), 
        .Y(n10) );
  AO22X1 U89 ( .A0(PCplus4_regI[3]), .A1(n134), .B0(PCplus4[3]), .B1(n132), 
        .Y(n38) );
  AO22X1 U90 ( .A0(PCplus4_regI[10]), .A1(n136), .B0(PCplus4[10]), .B1(n132), 
        .Y(n45) );
  AO22X1 U91 ( .A0(PCplus4_regI[6]), .A1(n136), .B0(PCplus4[6]), .B1(n132), 
        .Y(n41) );
  AO22X1 U92 ( .A0(PCplus4_regI[11]), .A1(n136), .B0(PCplus4[11]), .B1(n132), 
        .Y(n46) );
  AO22X1 U93 ( .A0(PCplus4_regI[13]), .A1(n136), .B0(PCplus4[13]), .B1(n132), 
        .Y(n48) );
  AO22X1 U94 ( .A0(PCplus4_regI[7]), .A1(n136), .B0(PCplus4[7]), .B1(n132), 
        .Y(n42) );
  AO22X1 U95 ( .A0(PCplus4_regI[8]), .A1(n136), .B0(PCplus4[8]), .B1(n132), 
        .Y(n43) );
  AO22X1 U96 ( .A0(PCplus4_regI[9]), .A1(n136), .B0(PCplus4[9]), .B1(n132), 
        .Y(n44) );
  AO22X1 U97 ( .A0(PCplus4_regI[12]), .A1(n136), .B0(PCplus4[12]), .B1(n132), 
        .Y(n47) );
  AO22X1 U98 ( .A0(PCplus4_regI[14]), .A1(n136), .B0(PCplus4[14]), .B1(n132), 
        .Y(n49) );
  AO22X1 U99 ( .A0(PCplus4_regI[15]), .A1(n136), .B0(PCplus4[15]), .B1(n132), 
        .Y(n50) );
  AO22X1 U100 ( .A0(PCplus4_regI[16]), .A1(n137), .B0(PCplus4[16]), .B1(n1), 
        .Y(n51) );
  AO22X1 U101 ( .A0(PCplus4_regI[17]), .A1(n137), .B0(PCplus4[17]), .B1(n130), 
        .Y(n52) );
  AO22X1 U102 ( .A0(PCplus4_regI[18]), .A1(n137), .B0(PCplus4[18]), .B1(n1), 
        .Y(n53) );
  AO22X1 U103 ( .A0(PCplus4_regI[19]), .A1(n137), .B0(PCplus4[19]), .B1(n130), 
        .Y(n54) );
  AO22X1 U104 ( .A0(PCplus4_regI[20]), .A1(n137), .B0(PCplus4[20]), .B1(n130), 
        .Y(n55) );
  AO22X1 U105 ( .A0(PCplus4_regI[21]), .A1(n137), .B0(PCplus4[21]), .B1(n130), 
        .Y(n56) );
  AO22X1 U106 ( .A0(PCplus4_regI[22]), .A1(n137), .B0(PCplus4[22]), .B1(n1), 
        .Y(n57) );
  AO22X1 U107 ( .A0(PCplus4_regI[23]), .A1(n137), .B0(PCplus4[23]), .B1(n131), 
        .Y(n58) );
  AO22X1 U108 ( .A0(PCplus4_regI[24]), .A1(n137), .B0(PCplus4[24]), .B1(n130), 
        .Y(n59) );
  AO22X1 U109 ( .A0(PCplus4_regI[25]), .A1(n137), .B0(PCplus4[25]), .B1(n130), 
        .Y(n60) );
  AO22X1 U110 ( .A0(PCplus4_regI[26]), .A1(n137), .B0(PCplus4[26]), .B1(n131), 
        .Y(n61) );
  AO22X1 U111 ( .A0(PCplus4_regI[5]), .A1(n136), .B0(PCplus4[5]), .B1(n132), 
        .Y(n40) );
  AO22X1 U112 ( .A0(PCplus4_regI[0]), .A1(n134), .B0(PCplus4[0]), .B1(n132), 
        .Y(n35) );
  AO22X1 U113 ( .A0(PCplus4_regI[1]), .A1(n133), .B0(PCplus4[1]), .B1(n131), 
        .Y(n36) );
  AO22X1 U114 ( .A0(PCplus4_regI[2]), .A1(n133), .B0(PCplus4[2]), .B1(n131), 
        .Y(n37) );
  CLKBUFX3 U115 ( .A(funct[1]), .Y(immediate[1]) );
  CLKBUFX3 U116 ( .A(funct[0]), .Y(branchOffset[0]) );
  CLKBUFX3 U117 ( .A(funct[1]), .Y(branchOffset[1]) );
  CLKBUFX3 U118 ( .A(funct[0]), .Y(immediate[0]) );
  CLKBUFX3 U119 ( .A(Rd[4]), .Y(immediate[15]) );
  CLKBUFX3 U120 ( .A(Rd[4]), .Y(branchOffset[15]) );
  CLKBUFX3 U121 ( .A(Rd[3]), .Y(immediate[14]) );
  CLKBUFX3 U122 ( .A(Rd[3]), .Y(branchOffset[14]) );
  CLKBUFX3 U123 ( .A(Rd[2]), .Y(immediate[13]) );
  CLKBUFX3 U124 ( .A(Rd[2]), .Y(branchOffset[13]) );
  CLKBUFX3 U125 ( .A(Rd[1]), .Y(immediate[12]) );
  CLKBUFX3 U126 ( .A(Rd[1]), .Y(branchOffset[12]) );
  CLKBUFX3 U127 ( .A(Rd[0]), .Y(immediate[11]) );
  CLKBUFX3 U128 ( .A(Rd[0]), .Y(branchOffset[11]) );
  CLKBUFX3 U129 ( .A(shamt[4]), .Y(immediate[10]) );
  CLKBUFX3 U130 ( .A(shamt[4]), .Y(branchOffset[10]) );
  CLKBUFX3 U131 ( .A(shamt[3]), .Y(immediate[9]) );
  CLKBUFX3 U132 ( .A(shamt[3]), .Y(branchOffset[9]) );
  CLKBUFX3 U133 ( .A(shamt[2]), .Y(immediate[8]) );
  CLKBUFX3 U134 ( .A(shamt[2]), .Y(branchOffset[8]) );
  CLKBUFX3 U135 ( .A(shamt[1]), .Y(immediate[7]) );
  CLKBUFX3 U136 ( .A(shamt[1]), .Y(branchOffset[7]) );
  CLKBUFX3 U137 ( .A(shamt[0]), .Y(immediate[6]) );
  CLKBUFX3 U138 ( .A(shamt[0]), .Y(branchOffset[6]) );
  CLKBUFX3 U139 ( .A(funct[5]), .Y(immediate[5]) );
  CLKBUFX3 U140 ( .A(funct[5]), .Y(branchOffset[5]) );
  CLKBUFX3 U141 ( .A(funct[4]), .Y(immediate[4]) );
  CLKBUFX3 U142 ( .A(funct[4]), .Y(branchOffset[4]) );
  CLKBUFX3 U143 ( .A(funct[3]), .Y(immediate[3]) );
  CLKBUFX3 U144 ( .A(funct[3]), .Y(branchOffset[3]) );
  CLKBUFX3 U145 ( .A(funct[2]), .Y(immediate[2]) );
  CLKBUFX3 U146 ( .A(funct[2]), .Y(branchOffset[2]) );
  AO22X1 U147 ( .A0(PCplus4_regI[31]), .A1(n133), .B0(PCplus4[31]), .B1(n1), 
        .Y(n66) );
  AO22X1 U148 ( .A0(opcode[2]), .A1(n148), .B0(instruction_next[28]), .B1(n132), .Y(n31) );
  AO22X1 U149 ( .A0(opcode[5]), .A1(n136), .B0(instruction_next[31]), .B1(n132), .Y(n34) );
endmodule


module DEC_EX_regFile ( clk, rst_n, stallcache, MemtoReg, ALUOp, JumpReg, 
        MemRead, MemWrite, ALUsrc, RegWrite, Branch, PCplus4_regI, funct, 
        branchOffset_D, A, B, ExtOut, Rs, Rt, wsel, MemtoReg_regD, ALUOp_regD, 
        MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, funct_regD, 
        A_regD, B_regD, ExtOut_regD, Rs_regD, Rt_regD, wsel_regD, JumpReg_regD, 
        Branch_regD, PCplus4_regD, branchOffset_regD );
  input [1:0] MemtoReg;
  input [5:0] ALUOp;
  input [31:0] PCplus4_regI;
  input [5:0] funct;
  input [15:0] branchOffset_D;
  input [31:0] A;
  input [31:0] B;
  input [31:0] ExtOut;
  input [4:0] Rs;
  input [4:0] Rt;
  input [4:0] wsel;
  output [1:0] MemtoReg_regD;
  output [5:0] ALUOp_regD;
  output [5:0] funct_regD;
  output [31:0] A_regD;
  output [31:0] B_regD;
  output [31:0] ExtOut_regD;
  output [4:0] Rs_regD;
  output [4:0] Rt_regD;
  output [4:0] wsel_regD;
  output [31:0] PCplus4_regD;
  output [15:0] branchOffset_regD;
  input clk, rst_n, stallcache, JumpReg, MemRead, MemWrite, ALUsrc, RegWrite,
         Branch;
  output MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, JumpReg_regD,
         Branch_regD;
  wire   n4, n11, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n111, n112, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n1, n2, n3, n5, n6, n7, n8, n9, n10,
         n12, n13, n14, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88;

  DFFRX1 \MemtoReg_regD_reg[1]  ( .D(n300), .CK(clk), .RN(n77), .Q(
        MemtoReg_regD[1]), .QN(n121) );
  DFFRX1 \MemtoReg_regD_reg[0]  ( .D(n299), .CK(clk), .RN(n77), .Q(
        MemtoReg_regD[0]), .QN(n120) );
  DFFRX1 MemWrite_regD_reg ( .D(n291), .CK(clk), .RN(n76), .Q(MemWrite_regD), 
        .QN(n112) );
  DFFRX1 RegWrite_regD_reg ( .D(n290), .CK(clk), .RN(n76), .Q(RegWrite_regD), 
        .QN(n111) );
  DFFRX1 \wsel_regD_reg[2]  ( .D(n180), .CK(clk), .RN(n67), .Q(wsel_regD[2])
         );
  DFFRX1 \wsel_regD_reg[4]  ( .D(n182), .CK(clk), .RN(n67), .Q(wsel_regD[4])
         );
  DFFRX1 \wsel_regD_reg[3]  ( .D(n181), .CK(clk), .RN(n67), .Q(wsel_regD[3])
         );
  DFFRX1 \wsel_regD_reg[1]  ( .D(n179), .CK(clk), .RN(n67), .Q(wsel_regD[1])
         );
  DFFRX1 \wsel_regD_reg[0]  ( .D(n178), .CK(clk), .RN(n67), .Q(wsel_regD[0])
         );
  DFFRX1 \PCplus4_regD_reg[1]  ( .D(n324), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[1]), .QN(n145) );
  DFFRX1 \PCplus4_regD_reg[0]  ( .D(n323), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[0]), .QN(n144) );
  DFFRX1 \funct_regD_reg[4]  ( .D(n305), .CK(clk), .RN(n77), .Q(funct_regD[4]), 
        .QN(n126) );
  DFFRX1 \branchOffset_regD_reg[15]  ( .D(n322), .CK(clk), .RN(n79), .Q(
        branchOffset_regD[15]), .QN(n143) );
  DFFRX1 \branchOffset_regD_reg[12]  ( .D(n319), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[12]), .QN(n140) );
  DFFRX1 \branchOffset_regD_reg[14]  ( .D(n321), .CK(clk), .RN(n79), .Q(
        branchOffset_regD[14]), .QN(n142) );
  DFFRX1 \branchOffset_regD_reg[13]  ( .D(n320), .CK(clk), .RN(n79), .Q(
        branchOffset_regD[13]), .QN(n141) );
  DFFRX1 \branchOffset_regD_reg[10]  ( .D(n317), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[10]), .QN(n138) );
  DFFRX1 \branchOffset_regD_reg[8]  ( .D(n315), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[8]), .QN(n136) );
  DFFRX1 \branchOffset_regD_reg[7]  ( .D(n314), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[7]), .QN(n135) );
  DFFRX1 \branchOffset_regD_reg[6]  ( .D(n313), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[6]), .QN(n134) );
  DFFRX1 \branchOffset_regD_reg[5]  ( .D(n312), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[5]), .QN(n133) );
  DFFRX1 \branchOffset_regD_reg[4]  ( .D(n311), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[4]), .QN(n132) );
  DFFRX1 \branchOffset_regD_reg[2]  ( .D(n309), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[2]), .QN(n130) );
  DFFRX1 \branchOffset_regD_reg[0]  ( .D(n307), .CK(clk), .RN(n77), .Q(
        branchOffset_regD[0]), .QN(n128) );
  DFFRX1 \branchOffset_regD_reg[9]  ( .D(n316), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[9]), .QN(n137) );
  DFFRX1 \PCplus4_regD_reg[30]  ( .D(n353), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[30]), .QN(n174) );
  DFFRX1 \PCplus4_regD_reg[29]  ( .D(n352), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[29]), .QN(n173) );
  DFFRX1 \PCplus4_regD_reg[28]  ( .D(n351), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[28]), .QN(n172) );
  DFFRX1 \PCplus4_regD_reg[27]  ( .D(n350), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[27]), .QN(n171) );
  DFFRX1 \PCplus4_regD_reg[26]  ( .D(n349), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[26]), .QN(n170) );
  DFFRX1 \PCplus4_regD_reg[25]  ( .D(n348), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[25]), .QN(n169) );
  DFFRX1 \PCplus4_regD_reg[24]  ( .D(n347), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[24]), .QN(n168) );
  DFFRX1 \PCplus4_regD_reg[23]  ( .D(n346), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[23]), .QN(n167) );
  DFFRX1 \PCplus4_regD_reg[22]  ( .D(n345), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[22]), .QN(n166) );
  DFFRX1 \PCplus4_regD_reg[21]  ( .D(n344), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[21]), .QN(n165) );
  DFFRX1 \PCplus4_regD_reg[20]  ( .D(n343), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[20]), .QN(n164) );
  DFFRX1 \PCplus4_regD_reg[19]  ( .D(n342), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[19]), .QN(n163) );
  DFFRX1 \PCplus4_regD_reg[18]  ( .D(n341), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[18]), .QN(n162) );
  DFFRX1 \PCplus4_regD_reg[17]  ( .D(n340), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[17]), .QN(n161) );
  DFFRX1 \PCplus4_regD_reg[16]  ( .D(n339), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[16]), .QN(n160) );
  DFFRX1 \PCplus4_regD_reg[15]  ( .D(n338), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[15]), .QN(n159) );
  DFFRX1 \PCplus4_regD_reg[14]  ( .D(n337), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[14]), .QN(n158) );
  DFFRX1 \PCplus4_regD_reg[12]  ( .D(n335), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[12]), .QN(n156) );
  DFFRX1 \PCplus4_regD_reg[9]  ( .D(n332), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[9]), .QN(n153) );
  DFFRX1 \PCplus4_regD_reg[8]  ( .D(n331), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[8]), .QN(n152) );
  DFFRX1 \PCplus4_regD_reg[7]  ( .D(n330), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[7]), .QN(n151) );
  DFFRX1 \PCplus4_regD_reg[6]  ( .D(n329), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[6]), .QN(n150) );
  DFFRX1 \PCplus4_regD_reg[2]  ( .D(n325), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[2]), .QN(n146) );
  DFFRX1 \PCplus4_regD_reg[11]  ( .D(n334), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[11]), .QN(n155) );
  DFFRX2 \funct_regD_reg[1]  ( .D(n302), .CK(clk), .RN(n77), .Q(funct_regD[1]), 
        .QN(n123) );
  DFFRX2 \funct_regD_reg[5]  ( .D(n306), .CK(clk), .RN(n77), .Q(funct_regD[5]), 
        .QN(n127) );
  DFFRX1 \ExtOut_regD_reg[28]  ( .D(n221), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[28]), .QN(n42) );
  DFFRX1 \ExtOut_regD_reg[24]  ( .D(n217), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[24]), .QN(n38) );
  DFFRX1 \ExtOut_regD_reg[21]  ( .D(n214), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[21]), .QN(n35) );
  DFFRX1 \ExtOut_regD_reg[20]  ( .D(n213), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[20]), .QN(n34) );
  DFFRX1 \ExtOut_regD_reg[18]  ( .D(n211), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[18]), .QN(n32) );
  DFFRX1 \ExtOut_regD_reg[17]  ( .D(n210), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[17]), .QN(n31) );
  DFFRX1 \ExtOut_regD_reg[16]  ( .D(n209), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[16]), .QN(n30) );
  DFFRX1 \ExtOut_regD_reg[12]  ( .D(n205), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[12]), .QN(n26) );
  DFFRX1 \ExtOut_regD_reg[10]  ( .D(n203), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[10]), .QN(n24) );
  DFFRX1 \ExtOut_regD_reg[9]  ( .D(n202), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[9]), .QN(n23) );
  DFFRX1 \ExtOut_regD_reg[8]  ( .D(n201), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[8]), .QN(n22) );
  DFFRX1 \ExtOut_regD_reg[5]  ( .D(n198), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[5]), .QN(n19) );
  DFFRX1 \ExtOut_regD_reg[4]  ( .D(n197), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[4]), .QN(n18) );
  DFFRX1 \ExtOut_regD_reg[1]  ( .D(n194), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[1]), .QN(n15) );
  DFFRX1 MemRead_regD_reg ( .D(n292), .CK(clk), .RN(n76), .Q(MemRead_regD) );
  DFFRX1 JumpReg_regD_reg ( .D(n177), .CK(clk), .RN(n67), .Q(JumpReg_regD) );
  DFFRX1 \A_regD_reg[30]  ( .D(n287), .CK(clk), .RN(n76), .Q(A_regD[30]) );
  DFFRX1 \A_regD_reg[15]  ( .D(n272), .CK(clk), .RN(n75), .Q(A_regD[15]) );
  DFFRX1 \A_regD_reg[13]  ( .D(n270), .CK(clk), .RN(n74), .Q(A_regD[13]) );
  DFFRX1 \B_regD_reg[25]  ( .D(n250), .CK(clk), .RN(n73), .Q(B_regD[25]) );
  DFFRX1 \A_regD_reg[31]  ( .D(n288), .CK(clk), .RN(n76), .Q(A_regD[31]) );
  DFFRX1 \A_regD_reg[29]  ( .D(n286), .CK(clk), .RN(n76), .Q(A_regD[29]) );
  DFFRX1 \A_regD_reg[28]  ( .D(n285), .CK(clk), .RN(n76), .Q(A_regD[28]) );
  DFFRX1 \A_regD_reg[27]  ( .D(n284), .CK(clk), .RN(n76), .Q(A_regD[27]) );
  DFFRX1 \A_regD_reg[26]  ( .D(n283), .CK(clk), .RN(n75), .Q(A_regD[26]) );
  DFFRX1 \A_regD_reg[25]  ( .D(n282), .CK(clk), .RN(n75), .Q(A_regD[25]) );
  DFFRX1 \A_regD_reg[24]  ( .D(n281), .CK(clk), .RN(n75), .Q(A_regD[24]) );
  DFFRX1 \A_regD_reg[23]  ( .D(n280), .CK(clk), .RN(n75), .Q(A_regD[23]) );
  DFFRX1 \A_regD_reg[22]  ( .D(n279), .CK(clk), .RN(n75), .Q(A_regD[22]) );
  DFFRX1 \A_regD_reg[21]  ( .D(n278), .CK(clk), .RN(n75), .Q(A_regD[21]) );
  DFFRX1 \A_regD_reg[20]  ( .D(n277), .CK(clk), .RN(n75), .Q(A_regD[20]) );
  DFFRX1 \A_regD_reg[19]  ( .D(n276), .CK(clk), .RN(n75), .Q(A_regD[19]) );
  DFFRX1 \A_regD_reg[18]  ( .D(n275), .CK(clk), .RN(n75), .Q(A_regD[18]) );
  DFFRX1 \A_regD_reg[17]  ( .D(n274), .CK(clk), .RN(n75), .Q(A_regD[17]) );
  DFFRX1 \A_regD_reg[16]  ( .D(n273), .CK(clk), .RN(n75), .Q(A_regD[16]) );
  DFFRX1 \A_regD_reg[14]  ( .D(n271), .CK(clk), .RN(n74), .Q(A_regD[14]) );
  DFFRX1 \A_regD_reg[12]  ( .D(n269), .CK(clk), .RN(n74), .Q(A_regD[12]) );
  DFFRX1 \A_regD_reg[11]  ( .D(n268), .CK(clk), .RN(n74), .Q(A_regD[11]) );
  DFFRX1 \A_regD_reg[10]  ( .D(n267), .CK(clk), .RN(n74), .Q(A_regD[10]) );
  DFFRX1 \A_regD_reg[9]  ( .D(n266), .CK(clk), .RN(n74), .Q(A_regD[9]) );
  DFFRX1 \A_regD_reg[8]  ( .D(n265), .CK(clk), .RN(n74), .Q(A_regD[8]) );
  DFFRX1 \A_regD_reg[7]  ( .D(n264), .CK(clk), .RN(n74), .Q(A_regD[7]) );
  DFFRX1 \A_regD_reg[6]  ( .D(n263), .CK(clk), .RN(n74), .Q(A_regD[6]) );
  DFFRX1 \A_regD_reg[5]  ( .D(n262), .CK(clk), .RN(n74), .Q(A_regD[5]) );
  DFFRX1 \A_regD_reg[4]  ( .D(n261), .CK(clk), .RN(n74), .Q(A_regD[4]) );
  DFFRX1 \A_regD_reg[3]  ( .D(n260), .CK(clk), .RN(n74), .Q(A_regD[3]) );
  DFFRX1 \A_regD_reg[2]  ( .D(n259), .CK(clk), .RN(n73), .Q(A_regD[2]) );
  DFFRX1 \A_regD_reg[1]  ( .D(n258), .CK(clk), .RN(n73), .Q(A_regD[1]) );
  DFFRX1 \A_regD_reg[0]  ( .D(n257), .CK(clk), .RN(n73), .Q(A_regD[0]) );
  DFFRX1 \B_regD_reg[31]  ( .D(n256), .CK(clk), .RN(n73), .Q(B_regD[31]) );
  DFFRX1 \B_regD_reg[30]  ( .D(n255), .CK(clk), .RN(n73), .Q(B_regD[30]) );
  DFFRX1 \B_regD_reg[29]  ( .D(n254), .CK(clk), .RN(n73), .Q(B_regD[29]) );
  DFFRX1 \B_regD_reg[28]  ( .D(n253), .CK(clk), .RN(n73), .Q(B_regD[28]) );
  DFFRX1 \B_regD_reg[27]  ( .D(n252), .CK(clk), .RN(n73), .Q(B_regD[27]) );
  DFFRX1 \B_regD_reg[26]  ( .D(n251), .CK(clk), .RN(n73), .Q(B_regD[26]) );
  DFFRX1 \B_regD_reg[24]  ( .D(n249), .CK(clk), .RN(n73), .Q(B_regD[24]) );
  DFFRX1 \B_regD_reg[23]  ( .D(n248), .CK(clk), .RN(n73), .Q(B_regD[23]) );
  DFFRX1 \B_regD_reg[22]  ( .D(n247), .CK(clk), .RN(n72), .Q(B_regD[22]) );
  DFFRX1 \B_regD_reg[21]  ( .D(n246), .CK(clk), .RN(n72), .Q(B_regD[21]) );
  DFFRX1 \B_regD_reg[20]  ( .D(n245), .CK(clk), .RN(n72), .Q(B_regD[20]) );
  DFFRX1 \B_regD_reg[19]  ( .D(n244), .CK(clk), .RN(n72), .Q(B_regD[19]) );
  DFFRX1 \B_regD_reg[18]  ( .D(n243), .CK(clk), .RN(n72), .Q(B_regD[18]) );
  DFFRX1 \B_regD_reg[17]  ( .D(n242), .CK(clk), .RN(n72), .Q(B_regD[17]) );
  DFFRX1 \B_regD_reg[16]  ( .D(n241), .CK(clk), .RN(n72), .Q(B_regD[16]) );
  DFFRX1 \B_regD_reg[15]  ( .D(n240), .CK(clk), .RN(n72), .Q(B_regD[15]) );
  DFFRX1 \B_regD_reg[14]  ( .D(n239), .CK(clk), .RN(n72), .Q(B_regD[14]) );
  DFFRX1 \B_regD_reg[13]  ( .D(n238), .CK(clk), .RN(n72), .Q(B_regD[13]) );
  DFFRX1 \B_regD_reg[12]  ( .D(n237), .CK(clk), .RN(n72), .Q(B_regD[12]) );
  DFFRX1 \B_regD_reg[11]  ( .D(n236), .CK(clk), .RN(n72), .Q(B_regD[11]) );
  DFFRX1 \B_regD_reg[10]  ( .D(n235), .CK(clk), .RN(n71), .Q(B_regD[10]) );
  DFFRX1 \B_regD_reg[9]  ( .D(n234), .CK(clk), .RN(n71), .Q(B_regD[9]) );
  DFFRX1 \B_regD_reg[8]  ( .D(n233), .CK(clk), .RN(n71), .Q(B_regD[8]) );
  DFFRX1 \B_regD_reg[7]  ( .D(n232), .CK(clk), .RN(n71), .Q(B_regD[7]) );
  DFFRX1 \B_regD_reg[6]  ( .D(n231), .CK(clk), .RN(n71), .Q(B_regD[6]) );
  DFFRX1 \B_regD_reg[5]  ( .D(n230), .CK(clk), .RN(n71), .Q(B_regD[5]) );
  DFFRX1 \B_regD_reg[4]  ( .D(n229), .CK(clk), .RN(n71), .Q(B_regD[4]) );
  DFFRX1 \B_regD_reg[3]  ( .D(n228), .CK(clk), .RN(n71), .Q(B_regD[3]) );
  DFFRX1 \B_regD_reg[2]  ( .D(n227), .CK(clk), .RN(n71), .Q(B_regD[2]) );
  DFFRX1 \B_regD_reg[1]  ( .D(n226), .CK(clk), .RN(n71), .Q(B_regD[1]) );
  DFFRX1 \B_regD_reg[0]  ( .D(n225), .CK(clk), .RN(n71), .Q(B_regD[0]) );
  DFFRX1 \ExtOut_regD_reg[31]  ( .D(n224), .CK(clk), .RN(n71), .Q(
        ExtOut_regD[31]), .QN(n45) );
  DFFRX1 \ExtOut_regD_reg[30]  ( .D(n223), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[30]), .QN(n44) );
  DFFRX1 \ExtOut_regD_reg[29]  ( .D(n222), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[29]), .QN(n43) );
  DFFRX1 \ExtOut_regD_reg[27]  ( .D(n220), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[27]), .QN(n41) );
  DFFRX1 \ExtOut_regD_reg[26]  ( .D(n219), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[26]), .QN(n40) );
  DFFRX1 \ExtOut_regD_reg[25]  ( .D(n218), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[25]), .QN(n39) );
  DFFRX1 \ExtOut_regD_reg[23]  ( .D(n216), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[23]), .QN(n37) );
  DFFRX1 \ExtOut_regD_reg[22]  ( .D(n215), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[22]), .QN(n36) );
  DFFRX1 \ExtOut_regD_reg[19]  ( .D(n212), .CK(clk), .RN(n70), .Q(
        ExtOut_regD[19]), .QN(n33) );
  DFFRX1 \ExtOut_regD_reg[15]  ( .D(n208), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[15]), .QN(n29) );
  DFFRX1 \ExtOut_regD_reg[14]  ( .D(n207), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[14]), .QN(n28) );
  DFFRX1 \ExtOut_regD_reg[13]  ( .D(n206), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[13]), .QN(n27) );
  DFFRX1 \ExtOut_regD_reg[11]  ( .D(n204), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[11]), .QN(n25) );
  DFFRX1 \ExtOut_regD_reg[7]  ( .D(n200), .CK(clk), .RN(n69), .Q(
        ExtOut_regD[7]), .QN(n21) );
  DFFRX1 \ExtOut_regD_reg[6]  ( .D(n199), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[6]), .QN(n20) );
  DFFRX1 \ExtOut_regD_reg[3]  ( .D(n196), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[3]), .QN(n17) );
  DFFRX1 \ExtOut_regD_reg[2]  ( .D(n195), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[2]), .QN(n16) );
  DFFRX1 \ExtOut_regD_reg[0]  ( .D(n193), .CK(clk), .RN(n68), .Q(
        ExtOut_regD[0]) );
  DFFRX1 \Rs_regD_reg[4]  ( .D(n192), .CK(clk), .RN(n68), .Q(Rs_regD[4]) );
  DFFRX1 \Rs_regD_reg[3]  ( .D(n191), .CK(clk), .RN(n68), .Q(Rs_regD[3]) );
  DFFRX1 Branch_regD_reg ( .D(n176), .CK(clk), .RN(n67), .Q(Branch_regD) );
  DFFRX1 \PCplus4_regD_reg[31]  ( .D(n354), .CK(clk), .RN(n81), .Q(
        PCplus4_regD[31]), .QN(n175) );
  DFFRX1 \branchOffset_regD_reg[3]  ( .D(n310), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[3]), .QN(n131) );
  DFFRX1 \branchOffset_regD_reg[1]  ( .D(n308), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[1]), .QN(n129) );
  DFFRX1 \PCplus4_regD_reg[10]  ( .D(n333), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[10]), .QN(n154) );
  DFFRX1 \PCplus4_regD_reg[5]  ( .D(n328), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[5]), .QN(n149) );
  DFFRX1 \PCplus4_regD_reg[3]  ( .D(n326), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[3]), .QN(n147) );
  DFFRX1 \PCplus4_regD_reg[4]  ( .D(n327), .CK(clk), .RN(n79), .Q(
        PCplus4_regD[4]), .QN(n148) );
  DFFRX1 \ALUOp_regD_reg[4]  ( .D(n297), .CK(clk), .RN(n77), .Q(ALUOp_regD[4]), 
        .QN(n118) );
  DFFRX1 \ALUOp_regD_reg[5]  ( .D(n298), .CK(clk), .RN(n77), .Q(ALUOp_regD[5]), 
        .QN(n119) );
  DFFRX1 \ALUOp_regD_reg[3]  ( .D(n296), .CK(clk), .RN(n77), .Q(ALUOp_regD[3]), 
        .QN(n117) );
  DFFRX1 \ALUOp_regD_reg[0]  ( .D(n293), .CK(clk), .RN(n76), .Q(ALUOp_regD[0]), 
        .QN(n114) );
  DFFRX1 \ALUOp_regD_reg[1]  ( .D(n294), .CK(clk), .RN(n76), .Q(ALUOp_regD[1]), 
        .QN(n115) );
  DFFRX1 \ALUOp_regD_reg[2]  ( .D(n295), .CK(clk), .RN(n76), .Q(ALUOp_regD[2]), 
        .QN(n116) );
  DFFRX1 \funct_regD_reg[0]  ( .D(n301), .CK(clk), .RN(n77), .Q(funct_regD[0]), 
        .QN(n122) );
  DFFRX1 \branchOffset_regD_reg[11]  ( .D(n318), .CK(clk), .RN(n78), .Q(
        branchOffset_regD[11]), .QN(n139) );
  DFFRX1 \PCplus4_regD_reg[13]  ( .D(n336), .CK(clk), .RN(n80), .Q(
        PCplus4_regD[13]), .QN(n157) );
  DFFRX1 \funct_regD_reg[2]  ( .D(n303), .CK(clk), .RN(n77), .Q(funct_regD[2]), 
        .QN(n124) );
  DFFRX1 \funct_regD_reg[3]  ( .D(n304), .CK(clk), .RN(n77), .Q(funct_regD[3]), 
        .QN(n125) );
  DFFRX1 ALUsrc_regD_reg ( .D(n289), .CK(clk), .RN(n76), .Q(ALUsrc_regD) );
  DFFRX1 \Rs_regD_reg[2]  ( .D(n190), .CK(clk), .RN(n68), .Q(Rs_regD[2]), .QN(
        n11) );
  DFFRX1 \Rt_regD_reg[0]  ( .D(n183), .CK(clk), .RN(n67), .Q(Rt_regD[0]), .QN(
        n4) );
  DFFRX4 \Rt_regD_reg[1]  ( .D(n184), .CK(clk), .RN(n67), .Q(Rt_regD[1]) );
  DFFRX2 \Rs_regD_reg[0]  ( .D(n188), .CK(clk), .RN(n68), .Q(Rs_regD[0]) );
  DFFRX2 \Rt_regD_reg[4]  ( .D(n187), .CK(clk), .RN(n67), .Q(Rt_regD[4]) );
  DFFRX2 \Rt_regD_reg[2]  ( .D(n185), .CK(clk), .RN(n67), .Q(Rt_regD[2]) );
  DFFRX2 \Rs_regD_reg[1]  ( .D(n189), .CK(clk), .RN(n68), .Q(Rs_regD[1]) );
  DFFRX2 \Rt_regD_reg[3]  ( .D(n186), .CK(clk), .RN(n67), .Q(Rt_regD[3]) );
  CLKBUFX2 U2 ( .A(stallcache), .Y(n3) );
  INVX3 U3 ( .A(n50), .Y(n47) );
  CLKBUFX3 U4 ( .A(n63), .Y(n54) );
  CLKBUFX3 U5 ( .A(n60), .Y(n59) );
  CLKINVX3 U6 ( .A(n50), .Y(n48) );
  CLKBUFX2 U7 ( .A(n63), .Y(n53) );
  CLKBUFX2 U8 ( .A(n64), .Y(n52) );
  BUFX2 U9 ( .A(n65), .Y(n51) );
  MX2XL U10 ( .A(MemRead), .B(MemRead_regD), .S0(n59), .Y(n292) );
  INVXL U11 ( .A(n50), .Y(n49) );
  CLKBUFX2 U12 ( .A(n3), .Y(n2) );
  CLKBUFX2 U13 ( .A(n3), .Y(n1) );
  CLKBUFX2 U14 ( .A(rst_n), .Y(n66) );
  MX2XL U15 ( .A(ALUsrc), .B(ALUsrc_regD), .S0(n59), .Y(n289) );
  MX2XL U16 ( .A(Rs[2]), .B(n88), .S0(n54), .Y(n190) );
  MX2XL U17 ( .A(Rt[2]), .B(Rt_regD[2]), .S0(n53), .Y(n185) );
  MX2XL U18 ( .A(Rt[3]), .B(Rt_regD[3]), .S0(n53), .Y(n186) );
  MX2XL U19 ( .A(Rt[4]), .B(Rt_regD[4]), .S0(n53), .Y(n187) );
  MX2XL U20 ( .A(Rs[0]), .B(Rs_regD[0]), .S0(n53), .Y(n188) );
  MX2XL U21 ( .A(Rs[1]), .B(Rs_regD[1]), .S0(n53), .Y(n189) );
  MX2XL U22 ( .A(Rt[0]), .B(n87), .S0(n59), .Y(n183) );
  MX2XL U23 ( .A(Rt[1]), .B(Rt_regD[1]), .S0(n52), .Y(n184) );
  MX2XL U24 ( .A(JumpReg), .B(JumpReg_regD), .S0(n51), .Y(n177) );
  MX2XL U25 ( .A(Branch), .B(Branch_regD), .S0(n50), .Y(n176) );
  INVX3 U26 ( .A(n60), .Y(n12) );
  INVX3 U27 ( .A(n51), .Y(n46) );
  INVX3 U28 ( .A(n51), .Y(n14) );
  INVX3 U29 ( .A(n51), .Y(n13) );
  INVX3 U30 ( .A(n52), .Y(n9) );
  INVX3 U31 ( .A(n52), .Y(n8) );
  INVX3 U32 ( .A(n52), .Y(n7) );
  INVX3 U33 ( .A(n54), .Y(n10) );
  INVX3 U34 ( .A(n53), .Y(n6) );
  INVX3 U35 ( .A(n53), .Y(n5) );
  CLKBUFX3 U36 ( .A(n65), .Y(n50) );
  CLKBUFX3 U37 ( .A(n62), .Y(n55) );
  CLKBUFX3 U38 ( .A(n62), .Y(n56) );
  CLKBUFX3 U39 ( .A(n61), .Y(n57) );
  CLKBUFX3 U40 ( .A(n61), .Y(n58) );
  CLKBUFX3 U41 ( .A(n2), .Y(n63) );
  CLKBUFX3 U42 ( .A(n1), .Y(n65) );
  CLKBUFX3 U43 ( .A(n1), .Y(n64) );
  CLKBUFX3 U44 ( .A(n2), .Y(n62) );
  CLKBUFX3 U45 ( .A(n1), .Y(n61) );
  CLKBUFX3 U46 ( .A(n1), .Y(n60) );
  CLKBUFX3 U47 ( .A(n83), .Y(n68) );
  CLKBUFX3 U48 ( .A(n83), .Y(n69) );
  CLKBUFX3 U49 ( .A(n84), .Y(n70) );
  CLKBUFX3 U50 ( .A(n84), .Y(n71) );
  CLKBUFX3 U51 ( .A(n84), .Y(n72) );
  CLKBUFX3 U52 ( .A(n84), .Y(n73) );
  CLKBUFX3 U53 ( .A(n85), .Y(n74) );
  CLKBUFX3 U54 ( .A(n85), .Y(n75) );
  CLKBUFX3 U55 ( .A(n85), .Y(n76) );
  CLKBUFX3 U56 ( .A(n82), .Y(n77) );
  CLKBUFX3 U57 ( .A(n86), .Y(n78) );
  CLKBUFX3 U58 ( .A(n86), .Y(n79) );
  CLKBUFX3 U59 ( .A(n86), .Y(n80) );
  CLKBUFX3 U60 ( .A(n82), .Y(n81) );
  CLKBUFX3 U61 ( .A(n82), .Y(n67) );
  CLKBUFX3 U62 ( .A(n83), .Y(n82) );
  CLKBUFX3 U63 ( .A(n66), .Y(n83) );
  CLKBUFX3 U64 ( .A(n66), .Y(n84) );
  CLKBUFX3 U65 ( .A(n66), .Y(n85) );
  CLKBUFX3 U66 ( .A(n66), .Y(n86) );
  OAI2BB2XL U67 ( .B0(n15), .B1(n10), .A0N(ExtOut[1]), .A1N(n13), .Y(n194) );
  OAI2BB2XL U68 ( .B0(n16), .B1(n12), .A0N(ExtOut[2]), .A1N(n13), .Y(n195) );
  OAI2BB2XL U69 ( .B0(n17), .B1(n12), .A0N(ExtOut[3]), .A1N(n14), .Y(n196) );
  OAI2BB2XL U70 ( .B0(n18), .B1(n12), .A0N(ExtOut[4]), .A1N(n13), .Y(n197) );
  OAI2BB2XL U71 ( .B0(n19), .B1(n12), .A0N(ExtOut[5]), .A1N(n13), .Y(n198) );
  OAI2BB2XL U72 ( .B0(n20), .B1(n12), .A0N(ExtOut[6]), .A1N(n14), .Y(n199) );
  OAI2BB2XL U73 ( .B0(n21), .B1(n12), .A0N(ExtOut[7]), .A1N(n13), .Y(n200) );
  OAI2BB2XL U74 ( .B0(n22), .B1(n12), .A0N(ExtOut[8]), .A1N(n13), .Y(n201) );
  OAI2BB2XL U75 ( .B0(n23), .B1(n12), .A0N(ExtOut[9]), .A1N(n14), .Y(n202) );
  OAI2BB2XL U76 ( .B0(n24), .B1(n12), .A0N(ExtOut[10]), .A1N(n14), .Y(n203) );
  OAI2BB2XL U77 ( .B0(n25), .B1(n12), .A0N(ExtOut[11]), .A1N(n14), .Y(n204) );
  OAI2BB2XL U78 ( .B0(n26), .B1(n12), .A0N(ExtOut[12]), .A1N(n46), .Y(n205) );
  OAI2BB2XL U79 ( .B0(n27), .B1(n12), .A0N(ExtOut[13]), .A1N(n46), .Y(n206) );
  OAI2BB2XL U80 ( .B0(n28), .B1(n12), .A0N(ExtOut[14]), .A1N(n46), .Y(n207) );
  OAI2BB2XL U81 ( .B0(n29), .B1(n12), .A0N(ExtOut[15]), .A1N(n46), .Y(n208) );
  OAI2BB2XL U82 ( .B0(n30), .B1(n12), .A0N(ExtOut[16]), .A1N(n46), .Y(n209) );
  OAI2BB2XL U83 ( .B0(n31), .B1(n47), .A0N(ExtOut[17]), .A1N(n46), .Y(n210) );
  OAI2BB2XL U84 ( .B0(n32), .B1(n12), .A0N(ExtOut[18]), .A1N(n46), .Y(n211) );
  OAI2BB2XL U85 ( .B0(n33), .B1(n12), .A0N(ExtOut[19]), .A1N(n47), .Y(n212) );
  OAI2BB2XL U86 ( .B0(n34), .B1(n12), .A0N(ExtOut[20]), .A1N(n47), .Y(n213) );
  OAI2BB2XL U87 ( .B0(n35), .B1(n47), .A0N(ExtOut[21]), .A1N(n47), .Y(n214) );
  OAI2BB2XL U88 ( .B0(n36), .B1(n12), .A0N(ExtOut[22]), .A1N(n47), .Y(n215) );
  OAI2BB2XL U89 ( .B0(n37), .B1(n10), .A0N(ExtOut[23]), .A1N(n46), .Y(n216) );
  OAI2BB2XL U90 ( .B0(n38), .B1(n9), .A0N(ExtOut[24]), .A1N(n47), .Y(n217) );
  OAI2BB2XL U91 ( .B0(n39), .B1(n8), .A0N(ExtOut[25]), .A1N(n47), .Y(n218) );
  OAI2BB2XL U92 ( .B0(n40), .B1(n10), .A0N(ExtOut[26]), .A1N(n48), .Y(n219) );
  OAI2BB2XL U93 ( .B0(n41), .B1(n10), .A0N(ExtOut[27]), .A1N(n48), .Y(n220) );
  OAI2BB2XL U94 ( .B0(n42), .B1(n10), .A0N(ExtOut[28]), .A1N(n48), .Y(n221) );
  OAI2BB2XL U95 ( .B0(n43), .B1(n10), .A0N(ExtOut[29]), .A1N(n48), .Y(n222) );
  OAI2BB2XL U96 ( .B0(n44), .B1(n10), .A0N(ExtOut[30]), .A1N(n48), .Y(n223) );
  OAI2BB2XL U97 ( .B0(n45), .B1(n10), .A0N(ExtOut[31]), .A1N(n12), .Y(n224) );
  OAI2BB2XL U98 ( .B0(n111), .B1(n10), .A0N(RegWrite), .A1N(n48), .Y(n290) );
  OAI2BB2XL U99 ( .B0(n112), .B1(n10), .A0N(MemWrite), .A1N(n48), .Y(n291) );
  OAI2BB2XL U100 ( .B0(n114), .B1(n10), .A0N(ALUOp[0]), .A1N(n48), .Y(n293) );
  OAI2BB2XL U101 ( .B0(n115), .B1(n9), .A0N(ALUOp[1]), .A1N(n48), .Y(n294) );
  OAI2BB2XL U102 ( .B0(n116), .B1(n9), .A0N(ALUOp[2]), .A1N(n48), .Y(n295) );
  OAI2BB2XL U103 ( .B0(n117), .B1(n9), .A0N(ALUOp[3]), .A1N(n48), .Y(n296) );
  OAI2BB2XL U104 ( .B0(n118), .B1(n9), .A0N(ALUOp[4]), .A1N(n48), .Y(n297) );
  OAI2BB2XL U105 ( .B0(n119), .B1(n9), .A0N(ALUOp[5]), .A1N(n48), .Y(n298) );
  OAI2BB2XL U106 ( .B0(n120), .B1(n9), .A0N(MemtoReg[0]), .A1N(n48), .Y(n299)
         );
  OAI2BB2XL U107 ( .B0(n121), .B1(n9), .A0N(MemtoReg[1]), .A1N(n48), .Y(n300)
         );
  OAI2BB2XL U108 ( .B0(n122), .B1(n9), .A0N(funct[0]), .A1N(n48), .Y(n301) );
  OAI2BB2XL U109 ( .B0(n123), .B1(n9), .A0N(funct[1]), .A1N(n48), .Y(n302) );
  OAI2BB2XL U110 ( .B0(n124), .B1(n9), .A0N(funct[2]), .A1N(n47), .Y(n303) );
  OAI2BB2XL U111 ( .B0(n125), .B1(n9), .A0N(funct[3]), .A1N(n47), .Y(n304) );
  OAI2BB2XL U112 ( .B0(n126), .B1(n9), .A0N(funct[4]), .A1N(n47), .Y(n305) );
  OAI2BB2XL U113 ( .B0(n127), .B1(n8), .A0N(funct[5]), .A1N(n47), .Y(n306) );
  OAI2BB2XL U114 ( .B0(n128), .B1(n8), .A0N(branchOffset_D[0]), .A1N(n47), .Y(
        n307) );
  OAI2BB2XL U115 ( .B0(n129), .B1(n8), .A0N(branchOffset_D[1]), .A1N(n47), .Y(
        n308) );
  OAI2BB2XL U116 ( .B0(n130), .B1(n8), .A0N(branchOffset_D[2]), .A1N(n47), .Y(
        n309) );
  OAI2BB2XL U117 ( .B0(n131), .B1(n8), .A0N(branchOffset_D[3]), .A1N(n47), .Y(
        n310) );
  OAI2BB2XL U118 ( .B0(n132), .B1(n8), .A0N(branchOffset_D[4]), .A1N(n47), .Y(
        n311) );
  OAI2BB2XL U119 ( .B0(n133), .B1(n8), .A0N(branchOffset_D[5]), .A1N(n47), .Y(
        n312) );
  OAI2BB2XL U120 ( .B0(n134), .B1(n8), .A0N(branchOffset_D[6]), .A1N(n47), .Y(
        n313) );
  OAI2BB2XL U121 ( .B0(n135), .B1(n8), .A0N(branchOffset_D[7]), .A1N(n47), .Y(
        n314) );
  OAI2BB2XL U122 ( .B0(n136), .B1(n8), .A0N(branchOffset_D[8]), .A1N(n47), .Y(
        n315) );
  OAI2BB2XL U123 ( .B0(n137), .B1(n8), .A0N(branchOffset_D[9]), .A1N(n46), .Y(
        n316) );
  OAI2BB2XL U124 ( .B0(n138), .B1(n8), .A0N(branchOffset_D[10]), .A1N(n46), 
        .Y(n317) );
  OAI2BB2XL U125 ( .B0(n139), .B1(n7), .A0N(branchOffset_D[11]), .A1N(n46), 
        .Y(n318) );
  OAI2BB2XL U126 ( .B0(n140), .B1(n7), .A0N(branchOffset_D[12]), .A1N(n46), 
        .Y(n319) );
  OAI2BB2XL U127 ( .B0(n141), .B1(n7), .A0N(branchOffset_D[13]), .A1N(n46), 
        .Y(n320) );
  OAI2BB2XL U128 ( .B0(n142), .B1(n7), .A0N(branchOffset_D[14]), .A1N(n46), 
        .Y(n321) );
  OAI2BB2XL U129 ( .B0(n143), .B1(n7), .A0N(branchOffset_D[15]), .A1N(n46), 
        .Y(n322) );
  OAI2BB2XL U130 ( .B0(n144), .B1(n7), .A0N(PCplus4_regI[0]), .A1N(n46), .Y(
        n323) );
  OAI2BB2XL U131 ( .B0(n145), .B1(n7), .A0N(PCplus4_regI[1]), .A1N(n46), .Y(
        n324) );
  OAI2BB2XL U132 ( .B0(n146), .B1(n7), .A0N(PCplus4_regI[2]), .A1N(n46), .Y(
        n325) );
  OAI2BB2XL U133 ( .B0(n147), .B1(n7), .A0N(PCplus4_regI[3]), .A1N(n46), .Y(
        n326) );
  OAI2BB2XL U134 ( .B0(n148), .B1(n7), .A0N(PCplus4_regI[4]), .A1N(n14), .Y(
        n327) );
  OAI2BB2XL U135 ( .B0(n149), .B1(n7), .A0N(PCplus4_regI[5]), .A1N(n14), .Y(
        n328) );
  OAI2BB2XL U136 ( .B0(n150), .B1(n7), .A0N(PCplus4_regI[6]), .A1N(n14), .Y(
        n329) );
  OAI2BB2XL U137 ( .B0(n151), .B1(n6), .A0N(PCplus4_regI[7]), .A1N(n14), .Y(
        n330) );
  OAI2BB2XL U138 ( .B0(n152), .B1(n6), .A0N(PCplus4_regI[8]), .A1N(n14), .Y(
        n331) );
  OAI2BB2XL U139 ( .B0(n153), .B1(n6), .A0N(PCplus4_regI[9]), .A1N(n14), .Y(
        n332) );
  OAI2BB2XL U140 ( .B0(n154), .B1(n6), .A0N(PCplus4_regI[10]), .A1N(n14), .Y(
        n333) );
  OAI2BB2XL U141 ( .B0(n155), .B1(n6), .A0N(PCplus4_regI[11]), .A1N(n14), .Y(
        n334) );
  OAI2BB2XL U142 ( .B0(n156), .B1(n6), .A0N(PCplus4_regI[12]), .A1N(n14), .Y(
        n335) );
  OAI2BB2XL U143 ( .B0(n157), .B1(n6), .A0N(PCplus4_regI[13]), .A1N(n13), .Y(
        n336) );
  OAI2BB2XL U144 ( .B0(n158), .B1(n6), .A0N(PCplus4_regI[14]), .A1N(n13), .Y(
        n337) );
  OAI2BB2XL U145 ( .B0(n159), .B1(n6), .A0N(PCplus4_regI[15]), .A1N(n14), .Y(
        n338) );
  OAI2BB2XL U146 ( .B0(n160), .B1(n6), .A0N(PCplus4_regI[16]), .A1N(n13), .Y(
        n339) );
  OAI2BB2XL U147 ( .B0(n161), .B1(n6), .A0N(PCplus4_regI[17]), .A1N(n13), .Y(
        n340) );
  OAI2BB2XL U148 ( .B0(n162), .B1(n6), .A0N(PCplus4_regI[18]), .A1N(n14), .Y(
        n341) );
  OAI2BB2XL U149 ( .B0(n163), .B1(n5), .A0N(PCplus4_regI[19]), .A1N(n13), .Y(
        n342) );
  OAI2BB2XL U150 ( .B0(n164), .B1(n5), .A0N(PCplus4_regI[20]), .A1N(n13), .Y(
        n343) );
  OAI2BB2XL U151 ( .B0(n165), .B1(n5), .A0N(PCplus4_regI[21]), .A1N(n14), .Y(
        n344) );
  OAI2BB2XL U152 ( .B0(n166), .B1(n5), .A0N(PCplus4_regI[22]), .A1N(n13), .Y(
        n345) );
  OAI2BB2XL U153 ( .B0(n167), .B1(n5), .A0N(PCplus4_regI[23]), .A1N(n13), .Y(
        n346) );
  OAI2BB2XL U154 ( .B0(n168), .B1(n5), .A0N(PCplus4_regI[24]), .A1N(n14), .Y(
        n347) );
  OAI2BB2XL U155 ( .B0(n169), .B1(n5), .A0N(PCplus4_regI[25]), .A1N(n13), .Y(
        n348) );
  OAI2BB2XL U156 ( .B0(n170), .B1(n5), .A0N(PCplus4_regI[26]), .A1N(n13), .Y(
        n349) );
  OAI2BB2XL U157 ( .B0(n171), .B1(n5), .A0N(PCplus4_regI[27]), .A1N(n14), .Y(
        n350) );
  OAI2BB2XL U158 ( .B0(n172), .B1(n5), .A0N(PCplus4_regI[28]), .A1N(n13), .Y(
        n351) );
  OAI2BB2XL U159 ( .B0(n173), .B1(n5), .A0N(PCplus4_regI[29]), .A1N(n13), .Y(
        n352) );
  OAI2BB2XL U160 ( .B0(n174), .B1(n5), .A0N(PCplus4_regI[30]), .A1N(n13), .Y(
        n353) );
  OAI2BB2XL U161 ( .B0(n175), .B1(n10), .A0N(PCplus4_regI[31]), .A1N(n12), .Y(
        n354) );
  CLKINVX1 U162 ( .A(n11), .Y(n88) );
  CLKMX2X2 U163 ( .A(Rs[3]), .B(Rs_regD[3]), .S0(n54), .Y(n191) );
  CLKMX2X2 U164 ( .A(Rs[4]), .B(Rs_regD[4]), .S0(n54), .Y(n192) );
  CLKMX2X2 U165 ( .A(ExtOut[0]), .B(ExtOut_regD[0]), .S0(n54), .Y(n193) );
  CLKMX2X2 U166 ( .A(B[0]), .B(B_regD[0]), .S0(n54), .Y(n225) );
  CLKMX2X2 U167 ( .A(B[1]), .B(B_regD[1]), .S0(n54), .Y(n226) );
  CLKMX2X2 U168 ( .A(B[2]), .B(B_regD[2]), .S0(n54), .Y(n227) );
  CLKMX2X2 U169 ( .A(B[3]), .B(B_regD[3]), .S0(n54), .Y(n228) );
  CLKMX2X2 U170 ( .A(B[4]), .B(B_regD[4]), .S0(n54), .Y(n229) );
  CLKMX2X2 U171 ( .A(B[5]), .B(B_regD[5]), .S0(n54), .Y(n230) );
  CLKMX2X2 U172 ( .A(B[6]), .B(B_regD[6]), .S0(n54), .Y(n231) );
  CLKMX2X2 U173 ( .A(B[7]), .B(B_regD[7]), .S0(n54), .Y(n232) );
  CLKMX2X2 U174 ( .A(B[8]), .B(B_regD[8]), .S0(n55), .Y(n233) );
  CLKMX2X2 U175 ( .A(B[9]), .B(B_regD[9]), .S0(n55), .Y(n234) );
  CLKMX2X2 U176 ( .A(B[10]), .B(B_regD[10]), .S0(n55), .Y(n235) );
  CLKMX2X2 U177 ( .A(B[11]), .B(B_regD[11]), .S0(n55), .Y(n236) );
  CLKMX2X2 U178 ( .A(B[12]), .B(B_regD[12]), .S0(n55), .Y(n237) );
  CLKMX2X2 U179 ( .A(B[13]), .B(B_regD[13]), .S0(n55), .Y(n238) );
  CLKMX2X2 U180 ( .A(B[14]), .B(B_regD[14]), .S0(n55), .Y(n239) );
  CLKMX2X2 U181 ( .A(B[15]), .B(B_regD[15]), .S0(n55), .Y(n240) );
  CLKMX2X2 U182 ( .A(B[16]), .B(B_regD[16]), .S0(n55), .Y(n241) );
  CLKMX2X2 U183 ( .A(B[17]), .B(B_regD[17]), .S0(n55), .Y(n242) );
  CLKMX2X2 U184 ( .A(B[18]), .B(B_regD[18]), .S0(n55), .Y(n243) );
  CLKMX2X2 U185 ( .A(B[19]), .B(B_regD[19]), .S0(n55), .Y(n244) );
  CLKMX2X2 U186 ( .A(B[20]), .B(B_regD[20]), .S0(n56), .Y(n245) );
  CLKMX2X2 U187 ( .A(B[21]), .B(B_regD[21]), .S0(n56), .Y(n246) );
  CLKMX2X2 U188 ( .A(B[22]), .B(B_regD[22]), .S0(n56), .Y(n247) );
  CLKMX2X2 U189 ( .A(B[23]), .B(B_regD[23]), .S0(n56), .Y(n248) );
  CLKMX2X2 U190 ( .A(B[24]), .B(B_regD[24]), .S0(n56), .Y(n249) );
  CLKMX2X2 U191 ( .A(B[25]), .B(B_regD[25]), .S0(n56), .Y(n250) );
  CLKMX2X2 U192 ( .A(B[26]), .B(B_regD[26]), .S0(n56), .Y(n251) );
  CLKMX2X2 U193 ( .A(B[27]), .B(B_regD[27]), .S0(n56), .Y(n252) );
  CLKMX2X2 U194 ( .A(B[28]), .B(B_regD[28]), .S0(n56), .Y(n253) );
  CLKMX2X2 U195 ( .A(B[29]), .B(B_regD[29]), .S0(n56), .Y(n254) );
  CLKMX2X2 U196 ( .A(B[30]), .B(B_regD[30]), .S0(n56), .Y(n255) );
  CLKMX2X2 U197 ( .A(B[31]), .B(B_regD[31]), .S0(n56), .Y(n256) );
  CLKMX2X2 U198 ( .A(A[0]), .B(A_regD[0]), .S0(n57), .Y(n257) );
  CLKMX2X2 U199 ( .A(A[1]), .B(A_regD[1]), .S0(n57), .Y(n258) );
  CLKMX2X2 U200 ( .A(A[2]), .B(A_regD[2]), .S0(n57), .Y(n259) );
  CLKMX2X2 U201 ( .A(A[3]), .B(A_regD[3]), .S0(n57), .Y(n260) );
  CLKMX2X2 U202 ( .A(A[4]), .B(A_regD[4]), .S0(n57), .Y(n261) );
  CLKMX2X2 U203 ( .A(A[5]), .B(A_regD[5]), .S0(n57), .Y(n262) );
  CLKMX2X2 U204 ( .A(A[6]), .B(A_regD[6]), .S0(n57), .Y(n263) );
  CLKMX2X2 U205 ( .A(A[7]), .B(A_regD[7]), .S0(n57), .Y(n264) );
  CLKMX2X2 U206 ( .A(A[8]), .B(A_regD[8]), .S0(n57), .Y(n265) );
  CLKMX2X2 U207 ( .A(A[9]), .B(A_regD[9]), .S0(n57), .Y(n266) );
  CLKMX2X2 U208 ( .A(A[10]), .B(A_regD[10]), .S0(n57), .Y(n267) );
  CLKMX2X2 U209 ( .A(A[11]), .B(A_regD[11]), .S0(n57), .Y(n268) );
  CLKMX2X2 U210 ( .A(A[12]), .B(A_regD[12]), .S0(n58), .Y(n269) );
  CLKMX2X2 U211 ( .A(A[13]), .B(A_regD[13]), .S0(n58), .Y(n270) );
  CLKMX2X2 U212 ( .A(A[14]), .B(A_regD[14]), .S0(n58), .Y(n271) );
  CLKMX2X2 U213 ( .A(A[15]), .B(A_regD[15]), .S0(n58), .Y(n272) );
  CLKMX2X2 U214 ( .A(A[16]), .B(A_regD[16]), .S0(n58), .Y(n273) );
  CLKMX2X2 U215 ( .A(A[17]), .B(A_regD[17]), .S0(n58), .Y(n274) );
  CLKMX2X2 U216 ( .A(A[18]), .B(A_regD[18]), .S0(n58), .Y(n275) );
  CLKMX2X2 U217 ( .A(A[19]), .B(A_regD[19]), .S0(n58), .Y(n276) );
  CLKMX2X2 U218 ( .A(A[20]), .B(A_regD[20]), .S0(n58), .Y(n277) );
  CLKMX2X2 U219 ( .A(A[21]), .B(A_regD[21]), .S0(n58), .Y(n278) );
  CLKMX2X2 U220 ( .A(A[22]), .B(A_regD[22]), .S0(n58), .Y(n279) );
  CLKMX2X2 U221 ( .A(A[23]), .B(A_regD[23]), .S0(n58), .Y(n280) );
  CLKMX2X2 U222 ( .A(A[24]), .B(A_regD[24]), .S0(n59), .Y(n281) );
  CLKMX2X2 U223 ( .A(A[25]), .B(A_regD[25]), .S0(n59), .Y(n282) );
  CLKMX2X2 U224 ( .A(A[26]), .B(A_regD[26]), .S0(n59), .Y(n283) );
  CLKMX2X2 U225 ( .A(A[27]), .B(A_regD[27]), .S0(n59), .Y(n284) );
  CLKMX2X2 U226 ( .A(A[28]), .B(A_regD[28]), .S0(n59), .Y(n285) );
  CLKMX2X2 U227 ( .A(A[29]), .B(A_regD[29]), .S0(n59), .Y(n286) );
  CLKMX2X2 U228 ( .A(A[30]), .B(A_regD[30]), .S0(n59), .Y(n287) );
  CLKMX2X2 U229 ( .A(A[31]), .B(A_regD[31]), .S0(n59), .Y(n288) );
  CLKINVX1 U230 ( .A(n4), .Y(n87) );
  AO22X1 U231 ( .A0(wsel_regD[1]), .A1(n59), .B0(wsel[1]), .B1(n49), .Y(n179)
         );
  AO22X1 U232 ( .A0(wsel_regD[2]), .A1(n59), .B0(wsel[2]), .B1(n49), .Y(n180)
         );
  AO22X1 U233 ( .A0(wsel_regD[3]), .A1(n64), .B0(wsel[3]), .B1(n49), .Y(n181)
         );
  AO22X1 U234 ( .A0(wsel_regD[0]), .A1(n59), .B0(wsel[0]), .B1(n48), .Y(n178)
         );
  AO22X1 U235 ( .A0(wsel_regD[4]), .A1(n64), .B0(wsel[4]), .B1(n48), .Y(n182)
         );
endmodule


module EX_MEM_regFile ( clk, rst_n, stallcache, MemtoReg_regD, MemRead_regD, 
        MemWrite_regD, RegWrite_regD, B_regD, wsel_regD, ALUout, MemtoReg_regE, 
        MemRead_regE, MemWrite_regE, RegWrite_regE, B_regE, wsel_regE, 
        ALUout_regE );
  input [1:0] MemtoReg_regD;
  input [31:0] B_regD;
  input [4:0] wsel_regD;
  input [31:0] ALUout;
  output [1:0] MemtoReg_regE;
  output [31:0] B_regE;
  output [4:0] wsel_regE;
  output [31:0] ALUout_regE;
  input clk, rst_n, stallcache, MemRead_regD, MemWrite_regD, RegWrite_regD;
  output MemRead_regE, MemWrite_regE, RegWrite_regE;
  wire   n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n37, n38, n49, n54, n61, n64, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n1, n34, n35, n36, n40, n42,
         n44, n46, n48, n51, n53, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n206, n207;

  DFFRX4 \wsel_regE_reg[2]  ( .D(n110), .CK(clk), .RN(n194), .Q(wsel_regE[2])
         );
  DFFRX4 \wsel_regE_reg[1]  ( .D(n109), .CK(clk), .RN(n194), .Q(wsel_regE[1])
         );
  DFFRX4 \wsel_regE_reg[0]  ( .D(n108), .CK(clk), .RN(n194), .Q(wsel_regE[0])
         );
  DFFRX1 \MemtoReg_regE_reg[1]  ( .D(n107), .CK(clk), .RN(n194), .Q(
        MemtoReg_regE[1]), .QN(n38) );
  DFFRX1 \MemtoReg_regE_reg[0]  ( .D(n106), .CK(clk), .RN(n193), .Q(
        MemtoReg_regE[0]), .QN(n37) );
  DFFRX1 \ALUout_regE_reg[1]  ( .D(n114), .CK(clk), .RN(n194), .Q(
        ALUout_regE[1]) );
  DFFRX1 \ALUout_regE_reg[0]  ( .D(n113), .CK(clk), .RN(n194), .Q(
        ALUout_regE[0]) );
  DFFRX1 \ALUout_regE_reg[19]  ( .D(n132), .CK(clk), .RN(n196), .Q(
        ALUout_regE[19]) );
  DFFRX1 RegWrite_regE_reg ( .D(n103), .CK(clk), .RN(n193), .Q(RegWrite_regE)
         );
  DFFRX1 MemRead_regE_reg ( .D(n105), .CK(clk), .RN(n193), .Q(MemRead_regE) );
  DFFRX1 \ALUout_regE_reg[31]  ( .D(n144), .CK(clk), .RN(n197), .Q(
        ALUout_regE[31]) );
  DFFRX1 \ALUout_regE_reg[30]  ( .D(n143), .CK(clk), .RN(n197), .Q(
        ALUout_regE[30]) );
  DFFRX1 \ALUout_regE_reg[27]  ( .D(n140), .CK(clk), .RN(n196), .Q(
        ALUout_regE[27]) );
  DFFRX1 \ALUout_regE_reg[29]  ( .D(n142), .CK(clk), .RN(n196), .Q(
        ALUout_regE[29]) );
  DFFRX1 \ALUout_regE_reg[21]  ( .D(n134), .CK(clk), .RN(n196), .Q(
        ALUout_regE[21]) );
  DFFRX1 \ALUout_regE_reg[20]  ( .D(n133), .CK(clk), .RN(n196), .Q(
        ALUout_regE[20]) );
  DFFRX1 \ALUout_regE_reg[16]  ( .D(n129), .CK(clk), .RN(n195), .Q(
        ALUout_regE[16]) );
  DFFRX1 \ALUout_regE_reg[13]  ( .D(n126), .CK(clk), .RN(n195), .Q(
        ALUout_regE[13]) );
  DFFRX1 \ALUout_regE_reg[12]  ( .D(n125), .CK(clk), .RN(n195), .Q(
        ALUout_regE[12]) );
  DFFRX1 \ALUout_regE_reg[7]  ( .D(n120), .CK(clk), .RN(n195), .Q(
        ALUout_regE[7]) );
  DFFRX1 \ALUout_regE_reg[11]  ( .D(n124), .CK(clk), .RN(n195), .Q(
        ALUout_regE[11]) );
  DFFRX1 \ALUout_regE_reg[9]  ( .D(n122), .CK(clk), .RN(n195), .Q(
        ALUout_regE[9]) );
  DFFRX1 \ALUout_regE_reg[28]  ( .D(n141), .CK(clk), .RN(n196), .Q(
        ALUout_regE[28]) );
  DFFRX1 \ALUout_regE_reg[24]  ( .D(n137), .CK(clk), .RN(n196), .Q(
        ALUout_regE[24]) );
  DFFRX1 \ALUout_regE_reg[2]  ( .D(n115), .CK(clk), .RN(n194), .Q(
        ALUout_regE[2]) );
  DFFRX1 \B_regE_reg[0]  ( .D(n71), .CK(clk), .RN(n191), .Q(n239), .QN(n2) );
  DFFRX1 \B_regE_reg[1]  ( .D(n72), .CK(clk), .RN(n191), .Q(n238), .QN(n3) );
  DFFRX1 \B_regE_reg[2]  ( .D(n73), .CK(clk), .RN(n191), .Q(n237), .QN(n4) );
  DFFRX1 \B_regE_reg[3]  ( .D(n74), .CK(clk), .RN(n191), .Q(n236), .QN(n5) );
  DFFRX1 \B_regE_reg[4]  ( .D(n75), .CK(clk), .RN(n191), .Q(n235), .QN(n6) );
  DFFRX1 \B_regE_reg[5]  ( .D(n76), .CK(clk), .RN(n191), .Q(n234), .QN(n7) );
  DFFRX1 \B_regE_reg[6]  ( .D(n77), .CK(clk), .RN(n191), .Q(n233), .QN(n8) );
  DFFRX1 \B_regE_reg[7]  ( .D(n78), .CK(clk), .RN(n191), .Q(n232), .QN(n9) );
  DFFRX1 \B_regE_reg[8]  ( .D(n79), .CK(clk), .RN(n191), .Q(n231), .QN(n10) );
  DFFRX1 \B_regE_reg[9]  ( .D(n80), .CK(clk), .RN(n191), .Q(n230), .QN(n11) );
  DFFRX1 \B_regE_reg[10]  ( .D(n81), .CK(clk), .RN(n191), .Q(n229), .QN(n12)
         );
  DFFRX1 \B_regE_reg[11]  ( .D(n82), .CK(clk), .RN(n191), .Q(n228), .QN(n13)
         );
  DFFRX1 \B_regE_reg[12]  ( .D(n83), .CK(clk), .RN(n192), .Q(n227), .QN(n14)
         );
  DFFRX1 \B_regE_reg[13]  ( .D(n84), .CK(clk), .RN(n192), .Q(n226), .QN(n15)
         );
  DFFRX1 \B_regE_reg[14]  ( .D(n85), .CK(clk), .RN(n192), .Q(n225), .QN(n16)
         );
  DFFRX1 \B_regE_reg[15]  ( .D(n86), .CK(clk), .RN(n192), .Q(n224), .QN(n17)
         );
  DFFRX1 \B_regE_reg[16]  ( .D(n87), .CK(clk), .RN(n192), .Q(n223), .QN(n18)
         );
  DFFRX1 \B_regE_reg[17]  ( .D(n88), .CK(clk), .RN(n192), .Q(n222), .QN(n19)
         );
  DFFRX1 \B_regE_reg[18]  ( .D(n89), .CK(clk), .RN(n192), .Q(n221), .QN(n20)
         );
  DFFRX1 \B_regE_reg[19]  ( .D(n90), .CK(clk), .RN(n192), .Q(n220), .QN(n21)
         );
  DFFRX1 \B_regE_reg[20]  ( .D(n91), .CK(clk), .RN(n192), .Q(n219), .QN(n22)
         );
  DFFRX1 \B_regE_reg[21]  ( .D(n92), .CK(clk), .RN(n192), .Q(n218), .QN(n23)
         );
  DFFRX1 \B_regE_reg[22]  ( .D(n93), .CK(clk), .RN(n192), .Q(n217), .QN(n24)
         );
  DFFRX1 \B_regE_reg[23]  ( .D(n94), .CK(clk), .RN(n192), .Q(n216), .QN(n25)
         );
  DFFRX1 \B_regE_reg[24]  ( .D(n95), .CK(clk), .RN(n193), .Q(n215), .QN(n26)
         );
  DFFRX1 \B_regE_reg[25]  ( .D(n96), .CK(clk), .RN(n193), .Q(n214), .QN(n27)
         );
  DFFRX1 \B_regE_reg[26]  ( .D(n97), .CK(clk), .RN(n193), .Q(n213), .QN(n28)
         );
  DFFRX1 \B_regE_reg[27]  ( .D(n98), .CK(clk), .RN(n193), .Q(n212), .QN(n29)
         );
  DFFRX1 \B_regE_reg[28]  ( .D(n99), .CK(clk), .RN(n193), .Q(n211), .QN(n30)
         );
  DFFRX1 \B_regE_reg[29]  ( .D(n100), .CK(clk), .RN(n193), .Q(n210), .QN(n31)
         );
  DFFRX1 \B_regE_reg[30]  ( .D(n101), .CK(clk), .RN(n193), .Q(n209), .QN(n32)
         );
  DFFRX1 \B_regE_reg[31]  ( .D(n102), .CK(clk), .RN(n193), .Q(n208), .QN(n33)
         );
  DFFRX2 \ALUout_regE_reg[6]  ( .D(n119), .CK(clk), .RN(n195), .Q(
        ALUout_regE[6]) );
  DFFRX1 \ALUout_regE_reg[10]  ( .D(n123), .CK(clk), .RN(n195), .Q(n35), .QN(
        n49) );
  DFFRX1 \ALUout_regE_reg[15]  ( .D(n128), .CK(clk), .RN(n195), .Q(n34), .QN(
        n54) );
  DFFRX1 \ALUout_regE_reg[22]  ( .D(n135), .CK(clk), .RN(n196), .Q(n1), .QN(
        n61) );
  DFFRX2 \ALUout_regE_reg[25]  ( .D(n138), .CK(clk), .RN(n196), .QN(n64) );
  DFFRHQX2 \ALUout_regE_reg[4]  ( .D(n117), .CK(clk), .RN(n194), .Q(
        ALUout_regE[4]) );
  DFFRX2 \wsel_regE_reg[4]  ( .D(n112), .CK(clk), .RN(n194), .Q(wsel_regE[4])
         );
  DFFRX2 \wsel_regE_reg[3]  ( .D(n111), .CK(clk), .RN(n194), .Q(wsel_regE[3])
         );
  DFFSRHQX1 MemWrite_regE_reg ( .D(n104), .CK(clk), .SN(1'b1), .RN(rst_n), .Q(
        n207) );
  DFFSRHQX1 \ALUout_regE_reg[8]  ( .D(n121), .CK(clk), .SN(1'b1), .RN(rst_n), 
        .Q(n200) );
  DFFSRHQX1 \ALUout_regE_reg[14]  ( .D(n127), .CK(clk), .SN(1'b1), .RN(n195), 
        .Q(n201) );
  DFFSRHQX1 \ALUout_regE_reg[17]  ( .D(n130), .CK(clk), .SN(1'b1), .RN(n195), 
        .Q(n202) );
  DFFSRHQX1 \ALUout_regE_reg[3]  ( .D(n116), .CK(clk), .SN(1'b1), .RN(n194), 
        .Q(n199) );
  DFFSRHQX1 \ALUout_regE_reg[26]  ( .D(n139), .CK(clk), .SN(1'b1), .RN(n196), 
        .Q(n206) );
  DFFSRHQX2 \ALUout_regE_reg[18]  ( .D(n131), .CK(clk), .SN(1'b1), .RN(n196), 
        .Q(n203) );
  DFFSRHQX2 \ALUout_regE_reg[23]  ( .D(n136), .CK(clk), .SN(1'b1), .RN(n196), 
        .Q(n204) );
  DFFRX4 \ALUout_regE_reg[5]  ( .D(n118), .CK(clk), .RN(n194), .Q(
        ALUout_regE[5]) );
  CLKMX2X4 U2 ( .A(ALUout[28]), .B(ALUout_regE[28]), .S0(n183), .Y(n141) );
  MX2X2 U3 ( .A(ALUout[1]), .B(ALUout_regE[1]), .S0(n180), .Y(n114) );
  CLKMX2X2 U4 ( .A(ALUout[18]), .B(ALUout_regE[18]), .S0(n181), .Y(n131) );
  MX2X1 U5 ( .A(ALUout[29]), .B(ALUout_regE[29]), .S0(n183), .Y(n142) );
  MX2XL U6 ( .A(ALUout[5]), .B(ALUout_regE[5]), .S0(n184), .Y(n118) );
  INVX16 U7 ( .A(n48), .Y(ALUout_regE[8]) );
  CLKINVX1 U8 ( .A(n200), .Y(n48) );
  INVX16 U9 ( .A(n42), .Y(ALUout_regE[17]) );
  CLKINVX1 U10 ( .A(n202), .Y(n42) );
  INVX16 U11 ( .A(n53), .Y(ALUout_regE[18]) );
  CLKINVX1 U12 ( .A(n203), .Y(n53) );
  INVX16 U13 ( .A(n51), .Y(ALUout_regE[23]) );
  CLKINVX1 U14 ( .A(n204), .Y(n51) );
  INVX16 U15 ( .A(n36), .Y(MemWrite_regE) );
  CLKINVX1 U16 ( .A(n207), .Y(n36) );
  INVX16 U17 ( .A(n49), .Y(ALUout_regE[10]) );
  INVX16 U18 ( .A(n54), .Y(ALUout_regE[15]) );
  INVX16 U19 ( .A(n61), .Y(ALUout_regE[22]) );
  INVX16 U20 ( .A(n64), .Y(ALUout_regE[25]) );
  CLKMX2X2 U21 ( .A(ALUout[22]), .B(n1), .S0(n182), .Y(n135) );
  CLKMX2X2 U22 ( .A(ALUout[23]), .B(ALUout_regE[23]), .S0(n182), .Y(n136) );
  CLKMX2X2 U23 ( .A(ALUout[3]), .B(ALUout_regE[3]), .S0(n182), .Y(n116) );
  CLKMX2X2 U24 ( .A(ALUout[17]), .B(ALUout_regE[17]), .S0(n186), .Y(n130) );
  CLKMX2X2 U25 ( .A(ALUout[8]), .B(ALUout_regE[8]), .S0(n181), .Y(n121) );
  CLKMX2X2 U26 ( .A(ALUout[4]), .B(ALUout_regE[4]), .S0(n180), .Y(n117) );
  MX2X1 U27 ( .A(ALUout[12]), .B(ALUout_regE[12]), .S0(n181), .Y(n125) );
  CLKMX2X2 U28 ( .A(ALUout[21]), .B(ALUout_regE[21]), .S0(n182), .Y(n134) );
  CLKMX2X2 U29 ( .A(ALUout[27]), .B(ALUout_regE[27]), .S0(n183), .Y(n140) );
  CLKMX2X2 U30 ( .A(ALUout[31]), .B(ALUout_regE[31]), .S0(n184), .Y(n144) );
  INVX3 U31 ( .A(n180), .Y(n177) );
  INVX3 U32 ( .A(n188), .Y(n178) );
  INVX6 U33 ( .A(n188), .Y(n179) );
  INVX12 U34 ( .A(n199), .Y(n40) );
  CLKINVX20 U35 ( .A(n40), .Y(ALUout_regE[3]) );
  INVX12 U36 ( .A(n201), .Y(n44) );
  CLKINVX20 U37 ( .A(n44), .Y(ALUout_regE[14]) );
  INVX12 U38 ( .A(n206), .Y(n46) );
  CLKINVX20 U39 ( .A(n46), .Y(ALUout_regE[26]) );
  CLKMX2X2 U48 ( .A(ALUout[7]), .B(ALUout_regE[7]), .S0(n188), .Y(n120) );
  CLKMX2X6 U49 ( .A(ALUout[2]), .B(ALUout_regE[2]), .S0(n188), .Y(n115) );
  CLKMX2X6 U50 ( .A(ALUout[19]), .B(ALUout_regE[19]), .S0(n185), .Y(n132) );
  BUFX12 U51 ( .A(n208), .Y(B_regE[31]) );
  BUFX12 U52 ( .A(n209), .Y(B_regE[30]) );
  BUFX12 U53 ( .A(n210), .Y(B_regE[29]) );
  BUFX12 U54 ( .A(n211), .Y(B_regE[28]) );
  BUFX12 U55 ( .A(n212), .Y(B_regE[27]) );
  BUFX12 U56 ( .A(n213), .Y(B_regE[26]) );
  BUFX12 U57 ( .A(n214), .Y(B_regE[25]) );
  BUFX12 U58 ( .A(n215), .Y(B_regE[24]) );
  BUFX12 U59 ( .A(n216), .Y(B_regE[23]) );
  BUFX12 U60 ( .A(n217), .Y(B_regE[22]) );
  BUFX12 U61 ( .A(n218), .Y(B_regE[21]) );
  BUFX12 U62 ( .A(n219), .Y(B_regE[20]) );
  BUFX12 U63 ( .A(n220), .Y(B_regE[19]) );
  BUFX12 U64 ( .A(n221), .Y(B_regE[18]) );
  BUFX12 U65 ( .A(n222), .Y(B_regE[17]) );
  BUFX12 U66 ( .A(n223), .Y(B_regE[16]) );
  BUFX12 U67 ( .A(n224), .Y(B_regE[15]) );
  BUFX12 U68 ( .A(n225), .Y(B_regE[14]) );
  BUFX12 U69 ( .A(n226), .Y(B_regE[13]) );
  BUFX12 U70 ( .A(n227), .Y(B_regE[12]) );
  BUFX12 U71 ( .A(n228), .Y(B_regE[11]) );
  BUFX12 U72 ( .A(n229), .Y(B_regE[10]) );
  BUFX12 U73 ( .A(n230), .Y(B_regE[9]) );
  BUFX12 U74 ( .A(n231), .Y(B_regE[8]) );
  BUFX12 U75 ( .A(n232), .Y(B_regE[7]) );
  BUFX12 U76 ( .A(n233), .Y(B_regE[6]) );
  BUFX12 U77 ( .A(n234), .Y(B_regE[5]) );
  BUFX12 U78 ( .A(n235), .Y(B_regE[4]) );
  BUFX12 U79 ( .A(n236), .Y(B_regE[3]) );
  BUFX12 U80 ( .A(n237), .Y(B_regE[2]) );
  BUFX12 U81 ( .A(n238), .Y(B_regE[1]) );
  BUFX12 U82 ( .A(n239), .Y(B_regE[0]) );
  BUFX2 U83 ( .A(n176), .Y(n188) );
  CLKMX2X2 U84 ( .A(ALUout[30]), .B(ALUout_regE[30]), .S0(n184), .Y(n143) );
  CLKMX2X2 U85 ( .A(ALUout[14]), .B(ALUout_regE[14]), .S0(n181), .Y(n127) );
  CLKMX2X2 U86 ( .A(ALUout[26]), .B(ALUout_regE[26]), .S0(n183), .Y(n139) );
  CLKBUFX2 U87 ( .A(n176), .Y(n187) );
  CLKBUFX2 U88 ( .A(n176), .Y(n186) );
  CLKBUFX2 U89 ( .A(n176), .Y(n185) );
  CLKBUFX2 U90 ( .A(rst_n), .Y(n190) );
  CLKBUFX2 U91 ( .A(rst_n), .Y(n189) );
  MX2X1 U92 ( .A(ALUout[25]), .B(ALUout_regE[25]), .S0(n183), .Y(n138) );
  MX2X1 U93 ( .A(ALUout[10]), .B(n35), .S0(n181), .Y(n123) );
  MX2XL U94 ( .A(ALUout[24]), .B(ALUout_regE[24]), .S0(n182), .Y(n137) );
  MX2XL U95 ( .A(ALUout[20]), .B(ALUout_regE[20]), .S0(n182), .Y(n133) );
  MX2XL U96 ( .A(ALUout[11]), .B(ALUout_regE[11]), .S0(n181), .Y(n124) );
  MX2XL U97 ( .A(ALUout[9]), .B(ALUout_regE[9]), .S0(n185), .Y(n122) );
  MX2XL U98 ( .A(ALUout[13]), .B(ALUout_regE[13]), .S0(n181), .Y(n126) );
  MX2XL U99 ( .A(ALUout[16]), .B(ALUout_regE[16]), .S0(n182), .Y(n129) );
  MX2XL U100 ( .A(wsel_regD[0]), .B(wsel_regE[0]), .S0(n184), .Y(n108) );
  MX2XL U101 ( .A(wsel_regD[1]), .B(wsel_regE[1]), .S0(n184), .Y(n109) );
  MX2XL U102 ( .A(wsel_regD[2]), .B(wsel_regE[2]), .S0(n184), .Y(n110) );
  MX2XL U103 ( .A(wsel_regD[3]), .B(wsel_regE[3]), .S0(n184), .Y(n111) );
  MX2XL U104 ( .A(wsel_regD[4]), .B(wsel_regE[4]), .S0(n183), .Y(n112) );
  MX2XL U105 ( .A(ALUout[6]), .B(ALUout_regE[6]), .S0(n183), .Y(n119) );
  MX2XL U106 ( .A(MemRead_regD), .B(MemRead_regE), .S0(n184), .Y(n105) );
  CLKBUFX3 U107 ( .A(n187), .Y(n180) );
  CLKBUFX3 U108 ( .A(n186), .Y(n181) );
  CLKBUFX3 U109 ( .A(n186), .Y(n182) );
  CLKBUFX3 U110 ( .A(n185), .Y(n183) );
  CLKBUFX3 U111 ( .A(n185), .Y(n184) );
  CLKBUFX3 U112 ( .A(stallcache), .Y(n176) );
  CLKBUFX3 U113 ( .A(n190), .Y(n192) );
  CLKBUFX3 U114 ( .A(n190), .Y(n193) );
  CLKBUFX3 U115 ( .A(n189), .Y(n194) );
  CLKBUFX3 U116 ( .A(n189), .Y(n196) );
  CLKBUFX3 U117 ( .A(n189), .Y(n195) );
  CLKBUFX3 U118 ( .A(n198), .Y(n197) );
  CLKBUFX3 U119 ( .A(n198), .Y(n191) );
  CLKBUFX3 U120 ( .A(n190), .Y(n198) );
  CLKMX2X2 U121 ( .A(ALUout[0]), .B(ALUout_regE[0]), .S0(n188), .Y(n113) );
  CLKMX2X2 U122 ( .A(ALUout[15]), .B(n34), .S0(n186), .Y(n128) );
  OAI2BB2XL U123 ( .B0(n2), .B1(n178), .A0N(B_regD[0]), .A1N(n179), .Y(n71) );
  OAI2BB2XL U124 ( .B0(n3), .B1(n178), .A0N(B_regD[1]), .A1N(n179), .Y(n72) );
  OAI2BB2XL U125 ( .B0(n4), .B1(n178), .A0N(B_regD[2]), .A1N(n179), .Y(n73) );
  OAI2BB2XL U126 ( .B0(n5), .B1(n178), .A0N(B_regD[3]), .A1N(n179), .Y(n74) );
  OAI2BB2XL U127 ( .B0(n6), .B1(n177), .A0N(B_regD[4]), .A1N(n179), .Y(n75) );
  OAI2BB2XL U128 ( .B0(n7), .B1(n178), .A0N(B_regD[5]), .A1N(n179), .Y(n76) );
  OAI2BB2XL U129 ( .B0(n8), .B1(n178), .A0N(B_regD[6]), .A1N(n179), .Y(n77) );
  OAI2BB2XL U130 ( .B0(n9), .B1(n178), .A0N(B_regD[7]), .A1N(n179), .Y(n78) );
  OAI2BB2XL U131 ( .B0(n10), .B1(n178), .A0N(B_regD[8]), .A1N(n179), .Y(n79)
         );
  OAI2BB2XL U132 ( .B0(n11), .B1(n178), .A0N(B_regD[9]), .A1N(n179), .Y(n80)
         );
  OAI2BB2XL U133 ( .B0(n12), .B1(n178), .A0N(B_regD[10]), .A1N(n179), .Y(n81)
         );
  OAI2BB2XL U134 ( .B0(n13), .B1(n177), .A0N(B_regD[11]), .A1N(n178), .Y(n82)
         );
  OAI2BB2XL U135 ( .B0(n14), .B1(n177), .A0N(B_regD[12]), .A1N(n178), .Y(n83)
         );
  OAI2BB2XL U136 ( .B0(n15), .B1(n177), .A0N(B_regD[13]), .A1N(n178), .Y(n84)
         );
  OAI2BB2XL U137 ( .B0(n16), .B1(n177), .A0N(B_regD[14]), .A1N(n178), .Y(n85)
         );
  OAI2BB2XL U138 ( .B0(n17), .B1(n177), .A0N(B_regD[15]), .A1N(n179), .Y(n86)
         );
  OAI2BB2XL U139 ( .B0(n18), .B1(n177), .A0N(B_regD[16]), .A1N(n179), .Y(n87)
         );
  OAI2BB2XL U140 ( .B0(n19), .B1(n177), .A0N(B_regD[17]), .A1N(n179), .Y(n88)
         );
  OAI2BB2XL U141 ( .B0(n20), .B1(n177), .A0N(B_regD[18]), .A1N(n179), .Y(n89)
         );
  OAI2BB2XL U142 ( .B0(n21), .B1(n177), .A0N(B_regD[19]), .A1N(n179), .Y(n90)
         );
  OAI2BB2XL U143 ( .B0(n22), .B1(n177), .A0N(B_regD[20]), .A1N(n179), .Y(n91)
         );
  OAI2BB2XL U144 ( .B0(n23), .B1(n177), .A0N(B_regD[21]), .A1N(n179), .Y(n92)
         );
  OAI2BB2XL U145 ( .B0(n24), .B1(n178), .A0N(B_regD[22]), .A1N(n179), .Y(n93)
         );
  OAI2BB2XL U146 ( .B0(n25), .B1(n177), .A0N(B_regD[23]), .A1N(n179), .Y(n94)
         );
  OAI2BB2XL U147 ( .B0(n26), .B1(n178), .A0N(B_regD[24]), .A1N(n179), .Y(n95)
         );
  OAI2BB2XL U148 ( .B0(n28), .B1(n177), .A0N(B_regD[26]), .A1N(n179), .Y(n97)
         );
  OAI2BB2XL U149 ( .B0(n29), .B1(n178), .A0N(B_regD[27]), .A1N(n179), .Y(n98)
         );
  OAI2BB2XL U150 ( .B0(n30), .B1(n177), .A0N(B_regD[28]), .A1N(n179), .Y(n99)
         );
  OAI2BB2XL U151 ( .B0(n31), .B1(n178), .A0N(B_regD[29]), .A1N(n179), .Y(n100)
         );
  OAI2BB2XL U152 ( .B0(n32), .B1(n177), .A0N(B_regD[30]), .A1N(n179), .Y(n101)
         );
  OAI2BB2XL U153 ( .B0(n33), .B1(n178), .A0N(B_regD[31]), .A1N(n179), .Y(n102)
         );
  OAI2BB2XL U154 ( .B0(n37), .B1(n178), .A0N(MemtoReg_regD[0]), .A1N(n179), 
        .Y(n106) );
  OAI2BB2XL U155 ( .B0(n38), .B1(n177), .A0N(MemtoReg_regD[1]), .A1N(n179), 
        .Y(n107) );
  CLKMX2X2 U156 ( .A(RegWrite_regD), .B(RegWrite_regE), .S0(n181), .Y(n103) );
  CLKMX2X2 U157 ( .A(MemWrite_regD), .B(MemWrite_regE), .S0(n185), .Y(n104) );
  OAI2BB2XL U158 ( .B0(n27), .B1(n177), .A0N(B_regD[25]), .A1N(n179), .Y(n96)
         );
endmodule


module MEM_WB_regFile ( clk, rst_n, stallcache, MemtoReg_regE, RegWrite_regE, 
        ALUout_regE, wsel_regE, dataOut, MemtoReg_regM, RegWrite_regM, 
        ALUout_regM, wsel_regM, dataOut_regM );
  input [1:0] MemtoReg_regE;
  input [31:0] ALUout_regE;
  input [4:0] wsel_regE;
  input [31:0] dataOut;
  output [1:0] MemtoReg_regM;
  output [31:0] ALUout_regM;
  output [4:0] wsel_regM;
  output [31:0] dataOut_regM;
  input clk, rst_n, stallcache, RegWrite_regE;
  output RegWrite_regM;
  wire   n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  DFFRX4 \wsel_regM_reg[2]  ( .D(n106), .CK(clk), .RN(n13), .Q(wsel_regM[2])
         );
  DFFRX4 \wsel_regM_reg[1]  ( .D(n105), .CK(clk), .RN(n13), .Q(wsel_regM[1])
         );
  DFFRX4 \wsel_regM_reg[0]  ( .D(n104), .CK(clk), .RN(n12), .Q(wsel_regM[0])
         );
  DFFRX1 \ALUout_regM_reg[25]  ( .D(n94), .CK(clk), .RN(n12), .Q(
        ALUout_regM[25]) );
  DFFRX1 \dataOut_regM_reg[30]  ( .D(n139), .CK(clk), .RN(n15), .Q(
        dataOut_regM[30]) );
  DFFRX1 \dataOut_regM_reg[19]  ( .D(n128), .CK(clk), .RN(n14), .Q(
        dataOut_regM[19]) );
  DFFRX1 \dataOut_regM_reg[15]  ( .D(n124), .CK(clk), .RN(n14), .Q(
        dataOut_regM[15]) );
  DFFRX1 \dataOut_regM_reg[13]  ( .D(n122), .CK(clk), .RN(n14), .Q(
        dataOut_regM[13]) );
  DFFRX1 \dataOut_regM_reg[2]  ( .D(n111), .CK(clk), .RN(n13), .Q(
        dataOut_regM[2]) );
  DFFRX1 \dataOut_regM_reg[31]  ( .D(n140), .CK(clk), .RN(n15), .Q(
        dataOut_regM[31]) );
  DFFRX1 \dataOut_regM_reg[29]  ( .D(n138), .CK(clk), .RN(n15), .Q(
        dataOut_regM[29]) );
  DFFRX1 \dataOut_regM_reg[28]  ( .D(n137), .CK(clk), .RN(n15), .Q(
        dataOut_regM[28]) );
  DFFRX1 \dataOut_regM_reg[27]  ( .D(n136), .CK(clk), .RN(n15), .Q(
        dataOut_regM[27]) );
  DFFRX1 \dataOut_regM_reg[26]  ( .D(n135), .CK(clk), .RN(n15), .Q(
        dataOut_regM[26]) );
  DFFRX1 \dataOut_regM_reg[25]  ( .D(n134), .CK(clk), .RN(n15), .Q(
        dataOut_regM[25]) );
  DFFRX1 \dataOut_regM_reg[24]  ( .D(n133), .CK(clk), .RN(n15), .Q(
        dataOut_regM[24]) );
  DFFRX1 \dataOut_regM_reg[23]  ( .D(n132), .CK(clk), .RN(n15), .Q(
        dataOut_regM[23]) );
  DFFRX1 \dataOut_regM_reg[21]  ( .D(n130), .CK(clk), .RN(n15), .Q(
        dataOut_regM[21]) );
  DFFRX1 \dataOut_regM_reg[20]  ( .D(n129), .CK(clk), .RN(n15), .Q(
        dataOut_regM[20]) );
  DFFRX1 \dataOut_regM_reg[18]  ( .D(n127), .CK(clk), .RN(n14), .Q(
        dataOut_regM[18]) );
  DFFRX1 \dataOut_regM_reg[17]  ( .D(n126), .CK(clk), .RN(n14), .Q(
        dataOut_regM[17]) );
  DFFRX1 \dataOut_regM_reg[16]  ( .D(n125), .CK(clk), .RN(n14), .Q(
        dataOut_regM[16]) );
  DFFRX1 \dataOut_regM_reg[14]  ( .D(n123), .CK(clk), .RN(n14), .Q(
        dataOut_regM[14]) );
  DFFRX1 \dataOut_regM_reg[12]  ( .D(n121), .CK(clk), .RN(n14), .Q(
        dataOut_regM[12]) );
  DFFRX1 \dataOut_regM_reg[11]  ( .D(n120), .CK(clk), .RN(n14), .Q(
        dataOut_regM[11]) );
  DFFRX1 \dataOut_regM_reg[10]  ( .D(n119), .CK(clk), .RN(n14), .Q(
        dataOut_regM[10]) );
  DFFRX1 \dataOut_regM_reg[9]  ( .D(n118), .CK(clk), .RN(n14), .Q(
        dataOut_regM[9]) );
  DFFRX1 \dataOut_regM_reg[8]  ( .D(n117), .CK(clk), .RN(n14), .Q(
        dataOut_regM[8]) );
  DFFRX1 \dataOut_regM_reg[7]  ( .D(n116), .CK(clk), .RN(n13), .Q(
        dataOut_regM[7]) );
  DFFRX1 \dataOut_regM_reg[6]  ( .D(n115), .CK(clk), .RN(n13), .Q(
        dataOut_regM[6]) );
  DFFRX1 \dataOut_regM_reg[5]  ( .D(n114), .CK(clk), .RN(n13), .Q(
        dataOut_regM[5]) );
  DFFRX1 \dataOut_regM_reg[4]  ( .D(n113), .CK(clk), .RN(n13), .Q(
        dataOut_regM[4]) );
  DFFRX1 \dataOut_regM_reg[3]  ( .D(n112), .CK(clk), .RN(n13), .Q(
        dataOut_regM[3]) );
  DFFRX1 \dataOut_regM_reg[1]  ( .D(n110), .CK(clk), .RN(n13), .Q(
        dataOut_regM[1]) );
  DFFRX1 \dataOut_regM_reg[0]  ( .D(n109), .CK(clk), .RN(n13), .Q(
        dataOut_regM[0]) );
  DFFRX1 \ALUout_regM_reg[31]  ( .D(n100), .CK(clk), .RN(n12), .Q(
        ALUout_regM[31]) );
  DFFRX1 \ALUout_regM_reg[30]  ( .D(n99), .CK(clk), .RN(n12), .Q(
        ALUout_regM[30]) );
  DFFRX1 \ALUout_regM_reg[29]  ( .D(n98), .CK(clk), .RN(n12), .Q(
        ALUout_regM[29]) );
  DFFRX1 \ALUout_regM_reg[28]  ( .D(n97), .CK(clk), .RN(n12), .Q(
        ALUout_regM[28]) );
  DFFRX1 \ALUout_regM_reg[27]  ( .D(n96), .CK(clk), .RN(n12), .Q(
        ALUout_regM[27]) );
  DFFRX1 \ALUout_regM_reg[26]  ( .D(n95), .CK(clk), .RN(n12), .Q(
        ALUout_regM[26]) );
  DFFRX1 \ALUout_regM_reg[24]  ( .D(n93), .CK(clk), .RN(n12), .Q(
        ALUout_regM[24]) );
  DFFRX1 \ALUout_regM_reg[23]  ( .D(n92), .CK(clk), .RN(n11), .Q(
        ALUout_regM[23]) );
  DFFRX1 \ALUout_regM_reg[22]  ( .D(n91), .CK(clk), .RN(n11), .Q(
        ALUout_regM[22]) );
  DFFRX1 \ALUout_regM_reg[21]  ( .D(n90), .CK(clk), .RN(n11), .Q(
        ALUout_regM[21]) );
  DFFRX1 \ALUout_regM_reg[20]  ( .D(n89), .CK(clk), .RN(n11), .Q(
        ALUout_regM[20]) );
  DFFRX1 \ALUout_regM_reg[19]  ( .D(n88), .CK(clk), .RN(n11), .Q(
        ALUout_regM[19]) );
  DFFRX1 \ALUout_regM_reg[18]  ( .D(n87), .CK(clk), .RN(n11), .Q(
        ALUout_regM[18]) );
  DFFRX1 \ALUout_regM_reg[17]  ( .D(n86), .CK(clk), .RN(n11), .Q(
        ALUout_regM[17]) );
  DFFRX1 \ALUout_regM_reg[16]  ( .D(n85), .CK(clk), .RN(n11), .Q(
        ALUout_regM[16]) );
  DFFRX1 \ALUout_regM_reg[15]  ( .D(n84), .CK(clk), .RN(n11), .Q(
        ALUout_regM[15]) );
  DFFRX1 \ALUout_regM_reg[14]  ( .D(n83), .CK(clk), .RN(n11), .Q(
        ALUout_regM[14]) );
  DFFRX1 \ALUout_regM_reg[13]  ( .D(n82), .CK(clk), .RN(n11), .Q(
        ALUout_regM[13]) );
  DFFRX1 \ALUout_regM_reg[12]  ( .D(n81), .CK(clk), .RN(n11), .Q(
        ALUout_regM[12]) );
  DFFRX1 \ALUout_regM_reg[11]  ( .D(n80), .CK(clk), .RN(n10), .Q(
        ALUout_regM[11]) );
  DFFRX1 \ALUout_regM_reg[10]  ( .D(n79), .CK(clk), .RN(n10), .Q(
        ALUout_regM[10]) );
  DFFRX1 \ALUout_regM_reg[9]  ( .D(n78), .CK(clk), .RN(n10), .Q(ALUout_regM[9]) );
  DFFRX1 \ALUout_regM_reg[8]  ( .D(n77), .CK(clk), .RN(n10), .Q(ALUout_regM[8]) );
  DFFRX1 \ALUout_regM_reg[7]  ( .D(n76), .CK(clk), .RN(n10), .Q(ALUout_regM[7]) );
  DFFRX1 \ALUout_regM_reg[6]  ( .D(n75), .CK(clk), .RN(n10), .Q(ALUout_regM[6]) );
  DFFRX1 \ALUout_regM_reg[5]  ( .D(n74), .CK(clk), .RN(n10), .Q(ALUout_regM[5]) );
  DFFRX1 \ALUout_regM_reg[4]  ( .D(n73), .CK(clk), .RN(n10), .Q(ALUout_regM[4]) );
  DFFRX1 \ALUout_regM_reg[3]  ( .D(n72), .CK(clk), .RN(n10), .Q(ALUout_regM[3]) );
  DFFRX1 \ALUout_regM_reg[2]  ( .D(n71), .CK(clk), .RN(n10), .Q(ALUout_regM[2]) );
  DFFRX1 \ALUout_regM_reg[1]  ( .D(n70), .CK(clk), .RN(n10), .Q(ALUout_regM[1]) );
  DFFRX1 \ALUout_regM_reg[0]  ( .D(n69), .CK(clk), .RN(n10), .Q(ALUout_regM[0]) );
  DFFRX2 \wsel_regM_reg[4]  ( .D(n108), .CK(clk), .RN(n13), .Q(wsel_regM[4])
         );
  DFFRX1 RegWrite_regM_reg ( .D(n101), .CK(clk), .RN(n12), .Q(RegWrite_regM)
         );
  DFFRX4 \MemtoReg_regM_reg[0]  ( .D(n102), .CK(clk), .RN(n12), .Q(
        MemtoReg_regM[0]) );
  DFFRX1 \dataOut_regM_reg[22]  ( .D(n131), .CK(clk), .RN(n15), .Q(
        dataOut_regM[22]) );
  DFFRX2 \wsel_regM_reg[3]  ( .D(n107), .CK(clk), .RN(n13), .Q(wsel_regM[3])
         );
  DFFSRHQX2 \MemtoReg_regM_reg[1]  ( .D(n103), .CK(clk), .SN(1'b1), .RN(rst_n), 
        .Q(MemtoReg_regM[1]) );
  CLKBUFX3 U2 ( .A(n2), .Y(n7) );
  CLKBUFX2 U4 ( .A(n2), .Y(n8) );
  CLKBUFX2 U5 ( .A(rst_n), .Y(n9) );
  MX2X1 U6 ( .A(dataOut[0]), .B(dataOut_regM[0]), .S0(n3), .Y(n109) );
  MX2X1 U7 ( .A(dataOut[1]), .B(dataOut_regM[1]), .S0(n3), .Y(n110) );
  MX2X1 U8 ( .A(dataOut[2]), .B(dataOut_regM[2]), .S0(n3), .Y(n111) );
  MX2X1 U9 ( .A(dataOut[3]), .B(dataOut_regM[3]), .S0(n3), .Y(n112) );
  MX2X1 U10 ( .A(dataOut[4]), .B(dataOut_regM[4]), .S0(n3), .Y(n113) );
  MX2X1 U11 ( .A(dataOut[5]), .B(dataOut_regM[5]), .S0(n3), .Y(n114) );
  MX2X1 U12 ( .A(dataOut[6]), .B(dataOut_regM[6]), .S0(n3), .Y(n115) );
  MX2X1 U13 ( .A(dataOut[7]), .B(dataOut_regM[7]), .S0(n3), .Y(n116) );
  MX2X1 U14 ( .A(dataOut[8]), .B(dataOut_regM[8]), .S0(n3), .Y(n117) );
  MX2X1 U15 ( .A(dataOut[9]), .B(dataOut_regM[9]), .S0(n3), .Y(n118) );
  MX2X1 U16 ( .A(dataOut[10]), .B(dataOut_regM[10]), .S0(n3), .Y(n119) );
  MX2X1 U17 ( .A(dataOut[11]), .B(dataOut_regM[11]), .S0(n3), .Y(n120) );
  MX2X1 U18 ( .A(dataOut[12]), .B(dataOut_regM[12]), .S0(n3), .Y(n121) );
  MX2X1 U19 ( .A(dataOut[13]), .B(dataOut_regM[13]), .S0(n4), .Y(n122) );
  MX2X1 U20 ( .A(dataOut[14]), .B(dataOut_regM[14]), .S0(n4), .Y(n123) );
  MX2X1 U21 ( .A(dataOut[15]), .B(dataOut_regM[15]), .S0(n4), .Y(n124) );
  MX2X1 U22 ( .A(dataOut[16]), .B(dataOut_regM[16]), .S0(n4), .Y(n125) );
  MX2X1 U23 ( .A(dataOut[17]), .B(dataOut_regM[17]), .S0(n4), .Y(n126) );
  MX2X1 U24 ( .A(dataOut[18]), .B(dataOut_regM[18]), .S0(n4), .Y(n127) );
  MX2X1 U25 ( .A(dataOut[19]), .B(dataOut_regM[19]), .S0(n4), .Y(n128) );
  MX2X1 U26 ( .A(dataOut[20]), .B(dataOut_regM[20]), .S0(n4), .Y(n129) );
  MX2X1 U27 ( .A(dataOut[21]), .B(dataOut_regM[21]), .S0(n4), .Y(n130) );
  MX2X1 U28 ( .A(dataOut[22]), .B(dataOut_regM[22]), .S0(n4), .Y(n131) );
  MX2X1 U29 ( .A(dataOut[23]), .B(dataOut_regM[23]), .S0(n4), .Y(n132) );
  MX2X1 U30 ( .A(dataOut[24]), .B(dataOut_regM[24]), .S0(n4), .Y(n133) );
  MX2X1 U31 ( .A(dataOut[25]), .B(dataOut_regM[25]), .S0(n4), .Y(n134) );
  MX2X1 U32 ( .A(dataOut[26]), .B(dataOut_regM[26]), .S0(n5), .Y(n135) );
  MX2X1 U33 ( .A(dataOut[27]), .B(dataOut_regM[27]), .S0(n5), .Y(n136) );
  MX2X1 U34 ( .A(dataOut[28]), .B(dataOut_regM[28]), .S0(n5), .Y(n137) );
  MX2X1 U35 ( .A(dataOut[29]), .B(dataOut_regM[29]), .S0(n5), .Y(n138) );
  MX2X1 U36 ( .A(dataOut[30]), .B(dataOut_regM[30]), .S0(n5), .Y(n139) );
  MX2X1 U37 ( .A(dataOut[31]), .B(dataOut_regM[31]), .S0(n5), .Y(n140) );
  MX2XL U38 ( .A(wsel_regE[0]), .B(wsel_regM[0]), .S0(n5), .Y(n104) );
  MX2XL U39 ( .A(wsel_regE[1]), .B(wsel_regM[1]), .S0(n5), .Y(n105) );
  MX2XL U40 ( .A(wsel_regE[2]), .B(wsel_regM[2]), .S0(n5), .Y(n106) );
  MX2XL U41 ( .A(wsel_regE[3]), .B(wsel_regM[3]), .S0(n5), .Y(n107) );
  MX2XL U42 ( .A(wsel_regE[4]), .B(wsel_regM[4]), .S0(n5), .Y(n108) );
  MX2XL U43 ( .A(ALUout_regE[4]), .B(ALUout_regM[4]), .S0(n6), .Y(n73) );
  MX2XL U44 ( .A(ALUout_regE[5]), .B(ALUout_regM[5]), .S0(n6), .Y(n74) );
  MX2XL U45 ( .A(ALUout_regE[6]), .B(ALUout_regM[6]), .S0(n6), .Y(n75) );
  MX2XL U46 ( .A(RegWrite_regE), .B(RegWrite_regM), .S0(n6), .Y(n101) );
  MX2XL U47 ( .A(MemtoReg_regE[0]), .B(MemtoReg_regM[0]), .S0(n6), .Y(n102) );
  MX2XL U48 ( .A(MemtoReg_regE[1]), .B(MemtoReg_regM[1]), .S0(n5), .Y(n103) );
  CLKBUFX3 U49 ( .A(n8), .Y(n3) );
  CLKBUFX3 U50 ( .A(n8), .Y(n4) );
  CLKBUFX3 U51 ( .A(stallcache), .Y(n5) );
  CLKBUFX3 U52 ( .A(stallcache), .Y(n6) );
  CLKBUFX3 U53 ( .A(stallcache), .Y(n2) );
  CLKBUFX3 U54 ( .A(n17), .Y(n10) );
  CLKBUFX3 U55 ( .A(n17), .Y(n11) );
  CLKBUFX3 U56 ( .A(n9), .Y(n13) );
  CLKBUFX3 U57 ( .A(n16), .Y(n14) );
  CLKBUFX3 U58 ( .A(n16), .Y(n15) );
  CLKBUFX3 U59 ( .A(n17), .Y(n12) );
  CLKBUFX3 U60 ( .A(n9), .Y(n17) );
  CLKBUFX3 U61 ( .A(n9), .Y(n16) );
  MX2XL U62 ( .A(ALUout_regE[15]), .B(ALUout_regM[15]), .S0(n7), .Y(n84) );
  CLKMX2X2 U63 ( .A(ALUout_regE[17]), .B(ALUout_regM[17]), .S0(n7), .Y(n86) );
  CLKMX2X2 U64 ( .A(ALUout_regE[31]), .B(ALUout_regM[31]), .S0(n5), .Y(n100)
         );
  CLKMX2X2 U65 ( .A(ALUout_regE[7]), .B(ALUout_regM[7]), .S0(n6), .Y(n76) );
  CLKMX2X2 U66 ( .A(ALUout_regE[11]), .B(ALUout_regM[11]), .S0(n6), .Y(n80) );
  CLKMX2X2 U67 ( .A(ALUout_regE[21]), .B(ALUout_regM[21]), .S0(n7), .Y(n90) );
  CLKMX2X2 U68 ( .A(ALUout_regE[30]), .B(ALUout_regM[30]), .S0(n5), .Y(n99) );
  CLKMX2X2 U69 ( .A(ALUout_regE[16]), .B(ALUout_regM[16]), .S0(n7), .Y(n85) );
  CLKMX2X2 U70 ( .A(ALUout_regE[20]), .B(ALUout_regM[20]), .S0(n7), .Y(n89) );
  CLKMX2X2 U71 ( .A(ALUout_regE[18]), .B(ALUout_regM[18]), .S0(n7), .Y(n87) );
  CLKMX2X2 U72 ( .A(ALUout_regE[26]), .B(ALUout_regM[26]), .S0(n7), .Y(n95) );
  CLKMX2X2 U73 ( .A(ALUout_regE[27]), .B(ALUout_regM[27]), .S0(n6), .Y(n96) );
  CLKMX2X2 U74 ( .A(ALUout_regE[12]), .B(ALUout_regM[12]), .S0(n6), .Y(n81) );
  CLKMX2X2 U75 ( .A(ALUout_regE[29]), .B(ALUout_regM[29]), .S0(n6), .Y(n98) );
  CLKMX2X2 U76 ( .A(ALUout_regE[23]), .B(ALUout_regM[23]), .S0(n7), .Y(n92) );
  CLKMX2X2 U77 ( .A(ALUout_regE[19]), .B(ALUout_regM[19]), .S0(n6), .Y(n88) );
  CLKMX2X2 U78 ( .A(ALUout_regE[24]), .B(ALUout_regM[24]), .S0(n7), .Y(n93) );
  CLKMX2X2 U79 ( .A(ALUout_regE[0]), .B(ALUout_regM[0]), .S0(n5), .Y(n69) );
  CLKMX2X2 U80 ( .A(ALUout_regE[1]), .B(ALUout_regM[1]), .S0(n5), .Y(n70) );
  MX2XL U81 ( .A(ALUout_regE[25]), .B(ALUout_regM[25]), .S0(n7), .Y(n94) );
  MX2XL U82 ( .A(ALUout_regE[8]), .B(ALUout_regM[8]), .S0(n6), .Y(n77) );
  MX2XL U83 ( .A(ALUout_regE[14]), .B(ALUout_regM[14]), .S0(n6), .Y(n83) );
  MX2XL U84 ( .A(ALUout_regE[9]), .B(ALUout_regM[9]), .S0(n6), .Y(n78) );
  MX2XL U85 ( .A(ALUout_regE[13]), .B(ALUout_regM[13]), .S0(n6), .Y(n82) );
  MX2XL U86 ( .A(ALUout_regE[10]), .B(ALUout_regM[10]), .S0(n6), .Y(n79) );
  MX2XL U87 ( .A(ALUout_regE[28]), .B(ALUout_regM[28]), .S0(n5), .Y(n97) );
  MX2XL U88 ( .A(ALUout_regE[2]), .B(ALUout_regM[2]), .S0(n6), .Y(n71) );
  MX2XL U89 ( .A(ALUout_regE[3]), .B(ALUout_regM[3]), .S0(n6), .Y(n72) );
  MX2XL U90 ( .A(ALUout_regE[22]), .B(ALUout_regM[22]), .S0(n7), .Y(n91) );
endmodule


module maincontrol ( opcode, funct, RegDst, MemtoReg, ALUOp, Branch, MemRead, 
        MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp );
  input [5:0] opcode;
  input [5:0] funct;
  output [1:0] RegDst;
  output [1:0] MemtoReg;
  output [5:0] ALUOp;
  output Branch, MemRead, MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n8, n9, n29, n30, n31, n32, n33, n34, n35;

  NOR2X1 U3 ( .A(n13), .B(ALUOp[4]), .Y(RegDst[1]) );
  OAI221XL U4 ( .A0(n27), .A1(n32), .B0(n23), .B1(n30), .C0(n28), .Y(n19) );
  CLKINVX1 U5 ( .A(opcode[5]), .Y(n30) );
  OAI22XL U6 ( .A0(opcode[0]), .A1(n31), .B0(opcode[1]), .B1(n20), .Y(n14) );
  CLKBUFX3 U7 ( .A(RegDst[0]), .Y(ExtOp) );
  NAND2X1 U8 ( .A(n8), .B(n29), .Y(RegDst[0]) );
  CLKINVX1 U9 ( .A(n19), .Y(n8) );
  NAND3X1 U10 ( .A(n32), .B(n30), .C(n33), .Y(n11) );
  CLKINVX1 U11 ( .A(n25), .Y(n29) );
  OAI31XL U12 ( .A0(n29), .A1(ALUOp[4]), .A2(n16), .B0(n9), .Y(MemtoReg[1]) );
  CLKINVX1 U13 ( .A(RegDst[1]), .Y(n9) );
  CLKINVX1 U14 ( .A(n21), .Y(n34) );
  NOR2BX1 U15 ( .AN(n10), .B(ALUOp[4]), .Y(RegWrite) );
  OAI211X1 U16 ( .A0(n11), .A1(opcode[2]), .B0(n12), .C0(n13), .Y(n10) );
  NOR3X1 U17 ( .A(n31), .B(ALUOp[4]), .C(n15), .Y(MemWrite) );
  CLKBUFX3 U18 ( .A(opcode[0]), .Y(ALUOp[0]) );
  CLKBUFX3 U19 ( .A(opcode[1]), .Y(ALUOp[1]) );
  CLKBUFX3 U20 ( .A(opcode[2]), .Y(ALUOp[2]) );
  CLKBUFX3 U21 ( .A(opcode[3]), .Y(ALUOp[3]) );
  CLKBUFX3 U22 ( .A(opcode[5]), .Y(ALUOp[5]) );
  NAND3X1 U23 ( .A(n26), .B(n13), .C(n8), .Y(ALUsrc) );
  OAI31XL U24 ( .A0(n34), .A1(funct[3]), .A2(n22), .B0(n25), .Y(n26) );
  NOR3X1 U25 ( .A(n15), .B(ALUOp[4]), .C(opcode[3]), .Y(MemRead) );
  NOR4BX1 U26 ( .AN(opcode[2]), .B(ALUOp[4]), .C(opcode[3]), .D(n11), .Y(
        Branch) );
  AND3X2 U27 ( .A(funct[3]), .B(n24), .C(n25), .Y(JumpReg) );
  AOI31X1 U28 ( .A0(n20), .A1(n32), .A2(opcode[0]), .B0(ALUOp[4]), .Y(n28) );
  AOI32X1 U29 ( .A0(opcode[0]), .A1(n30), .A2(opcode[3]), .B0(opcode[2]), .B1(
        n31), .Y(n27) );
  NOR3X1 U30 ( .A(opcode[2]), .B(opcode[3]), .C(n11), .Y(n25) );
  CLKINVX1 U31 ( .A(opcode[3]), .Y(n31) );
  NOR2X1 U32 ( .A(n33), .B(opcode[2]), .Y(n23) );
  CLKINVX1 U33 ( .A(opcode[1]), .Y(n32) );
  CLKINVX1 U34 ( .A(opcode[0]), .Y(n33) );
  NAND2X1 U35 ( .A(opcode[3]), .B(opcode[2]), .Y(n20) );
  OAI211X1 U36 ( .A0(n35), .A1(n29), .B0(n17), .C0(n18), .Y(MemtoReg[0]) );
  OAI21XL U37 ( .A0(opcode[2]), .A1(opcode[1]), .B0(n33), .Y(n17) );
  CLKINVX1 U38 ( .A(n16), .Y(n35) );
  NOR2X1 U39 ( .A(n19), .B(n14), .Y(n18) );
  NOR3X1 U40 ( .A(funct[5]), .B(funct[4]), .C(funct[2]), .Y(n21) );
  NAND4X1 U41 ( .A(opcode[1]), .B(n23), .C(n31), .D(n30), .Y(n13) );
  NOR2BX1 U42 ( .AN(funct[0]), .B(funct[1]), .Y(n22) );
  NAND3X1 U43 ( .A(opcode[1]), .B(n23), .C(opcode[5]), .Y(n15) );
  NOR3X1 U44 ( .A(ALUOp[4]), .B(funct[1]), .C(n34), .Y(n24) );
  NAND3X1 U45 ( .A(n21), .B(n22), .C(funct[3]), .Y(n16) );
  AOI2BB2X1 U46 ( .B0(n30), .B1(n14), .A0N(opcode[3]), .A1N(n15), .Y(n12) );
  CLKBUFX3 U47 ( .A(opcode[4]), .Y(ALUOp[4]) );
endmodule


module registerFile ( clk, rst_n, rsel1, rsel2, wsel, wen, wdata, rdata1, 
        rdata2 );
  input [4:0] rsel1;
  input [4:0] rsel2;
  input [4:0] wsel;
  input [31:0] wdata;
  output [31:0] rdata1;
  output [31:0] rdata2;
  input clk, rst_n, wen;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, \register[31][31] ,
         \register[31][30] , \register[31][29] , \register[31][28] ,
         \register[31][27] , \register[31][26] , \register[31][25] ,
         \register[31][24] , \register[31][23] , \register[31][22] ,
         \register[31][21] , \register[31][20] , \register[31][19] ,
         \register[31][18] , \register[31][17] , \register[31][16] ,
         \register[31][15] , \register[31][14] , \register[31][13] ,
         \register[31][12] , \register[31][11] , \register[31][10] ,
         \register[31][9] , \register[31][8] , \register[31][7] ,
         \register[31][6] , \register[31][5] , \register[31][4] ,
         \register[31][3] , \register[31][2] , \register[31][1] ,
         \register[31][0] , \register[30][31] , \register[30][30] ,
         \register[30][29] , \register[30][28] , \register[30][27] ,
         \register[30][26] , \register[30][25] , \register[30][24] ,
         \register[30][23] , \register[30][22] , \register[30][21] ,
         \register[30][20] , \register[30][19] , \register[30][18] ,
         \register[30][17] , \register[30][16] , \register[30][15] ,
         \register[30][14] , \register[30][13] , \register[30][12] ,
         \register[30][11] , \register[30][10] , \register[30][9] ,
         \register[30][8] , \register[30][7] , \register[30][6] ,
         \register[30][5] , \register[30][4] , \register[30][3] ,
         \register[30][2] , \register[30][1] , \register[30][0] ,
         \register[29][31] , \register[29][30] , \register[29][29] ,
         \register[29][28] , \register[29][27] , \register[29][26] ,
         \register[29][25] , \register[29][24] , \register[29][23] ,
         \register[29][22] , \register[29][21] , \register[29][20] ,
         \register[29][19] , \register[29][18] , \register[29][17] ,
         \register[29][16] , \register[29][15] , \register[29][14] ,
         \register[29][13] , \register[29][12] , \register[29][11] ,
         \register[29][10] , \register[29][9] , \register[29][8] ,
         \register[29][7] , \register[29][6] , \register[29][5] ,
         \register[29][4] , \register[29][3] , \register[29][2] ,
         \register[29][1] , \register[29][0] , \register[28][31] ,
         \register[28][30] , \register[28][29] , \register[28][28] ,
         \register[28][27] , \register[28][26] , \register[28][25] ,
         \register[28][24] , \register[28][23] , \register[28][22] ,
         \register[28][21] , \register[28][20] , \register[28][19] ,
         \register[28][18] , \register[28][17] , \register[28][16] ,
         \register[28][15] , \register[28][14] , \register[28][13] ,
         \register[28][12] , \register[28][11] , \register[28][10] ,
         \register[28][9] , \register[28][8] , \register[28][7] ,
         \register[28][6] , \register[28][5] , \register[28][4] ,
         \register[28][3] , \register[28][2] , \register[28][1] ,
         \register[28][0] , \register[27][31] , \register[27][30] ,
         \register[27][29] , \register[27][28] , \register[27][27] ,
         \register[27][26] , \register[27][25] , \register[27][24] ,
         \register[27][23] , \register[27][22] , \register[27][21] ,
         \register[27][20] , \register[27][19] , \register[27][18] ,
         \register[27][17] , \register[27][16] , \register[27][15] ,
         \register[27][14] , \register[27][13] , \register[27][12] ,
         \register[27][11] , \register[27][10] , \register[27][9] ,
         \register[27][8] , \register[27][7] , \register[27][6] ,
         \register[27][5] , \register[27][4] , \register[27][3] ,
         \register[27][2] , \register[27][1] , \register[27][0] ,
         \register[26][31] , \register[26][30] , \register[26][29] ,
         \register[26][28] , \register[26][27] , \register[26][26] ,
         \register[26][25] , \register[26][24] , \register[26][23] ,
         \register[26][22] , \register[26][21] , \register[26][20] ,
         \register[26][19] , \register[26][18] , \register[26][17] ,
         \register[26][16] , \register[26][15] , \register[26][14] ,
         \register[26][13] , \register[26][12] , \register[26][11] ,
         \register[26][10] , \register[26][9] , \register[26][8] ,
         \register[26][7] , \register[26][6] , \register[26][5] ,
         \register[26][4] , \register[26][3] , \register[26][2] ,
         \register[26][1] , \register[26][0] , \register[25][31] ,
         \register[25][30] , \register[25][29] , \register[25][28] ,
         \register[25][27] , \register[25][26] , \register[25][25] ,
         \register[25][24] , \register[25][23] , \register[25][22] ,
         \register[25][21] , \register[25][20] , \register[25][19] ,
         \register[25][18] , \register[25][17] , \register[25][16] ,
         \register[25][15] , \register[25][14] , \register[25][13] ,
         \register[25][12] , \register[25][11] , \register[25][10] ,
         \register[25][9] , \register[25][8] , \register[25][7] ,
         \register[25][6] , \register[25][5] , \register[25][4] ,
         \register[25][3] , \register[25][2] , \register[25][1] ,
         \register[25][0] , \register[24][31] , \register[24][30] ,
         \register[24][29] , \register[24][28] , \register[24][27] ,
         \register[24][26] , \register[24][25] , \register[24][24] ,
         \register[24][23] , \register[24][22] , \register[24][21] ,
         \register[24][20] , \register[24][19] , \register[24][18] ,
         \register[24][17] , \register[24][16] , \register[24][15] ,
         \register[24][14] , \register[24][13] , \register[24][12] ,
         \register[24][11] , \register[24][10] , \register[24][9] ,
         \register[24][8] , \register[24][7] , \register[24][6] ,
         \register[24][5] , \register[24][4] , \register[24][3] ,
         \register[24][2] , \register[24][1] , \register[24][0] ,
         \register[23][31] , \register[23][30] , \register[23][29] ,
         \register[23][28] , \register[23][27] , \register[23][26] ,
         \register[23][25] , \register[23][24] , \register[23][23] ,
         \register[23][22] , \register[23][21] , \register[23][20] ,
         \register[23][19] , \register[23][18] , \register[23][17] ,
         \register[23][16] , \register[23][15] , \register[23][14] ,
         \register[23][13] , \register[23][12] , \register[23][11] ,
         \register[23][10] , \register[23][9] , \register[23][8] ,
         \register[23][7] , \register[23][6] , \register[23][5] ,
         \register[23][4] , \register[23][3] , \register[23][2] ,
         \register[23][1] , \register[23][0] , \register[22][31] ,
         \register[22][30] , \register[22][29] , \register[22][28] ,
         \register[22][27] , \register[22][26] , \register[22][25] ,
         \register[22][24] , \register[22][23] , \register[22][22] ,
         \register[22][21] , \register[22][20] , \register[22][19] ,
         \register[22][18] , \register[22][17] , \register[22][16] ,
         \register[22][15] , \register[22][14] , \register[22][13] ,
         \register[22][12] , \register[22][11] , \register[22][10] ,
         \register[22][9] , \register[22][8] , \register[22][7] ,
         \register[22][6] , \register[22][5] , \register[22][4] ,
         \register[22][3] , \register[22][2] , \register[22][1] ,
         \register[22][0] , \register[21][31] , \register[21][30] ,
         \register[21][29] , \register[21][28] , \register[21][27] ,
         \register[21][26] , \register[21][25] , \register[21][24] ,
         \register[21][23] , \register[21][22] , \register[21][21] ,
         \register[21][20] , \register[21][19] , \register[21][18] ,
         \register[21][17] , \register[21][16] , \register[21][15] ,
         \register[21][14] , \register[21][13] , \register[21][12] ,
         \register[21][11] , \register[21][10] , \register[21][9] ,
         \register[21][8] , \register[21][7] , \register[21][6] ,
         \register[21][5] , \register[21][4] , \register[21][3] ,
         \register[21][2] , \register[21][1] , \register[21][0] ,
         \register[20][31] , \register[20][30] , \register[20][29] ,
         \register[20][28] , \register[20][27] , \register[20][26] ,
         \register[20][25] , \register[20][24] , \register[20][23] ,
         \register[20][22] , \register[20][21] , \register[20][20] ,
         \register[20][19] , \register[20][18] , \register[20][17] ,
         \register[20][16] , \register[20][15] , \register[20][14] ,
         \register[20][13] , \register[20][12] , \register[20][11] ,
         \register[20][10] , \register[20][9] , \register[20][8] ,
         \register[20][7] , \register[20][6] , \register[20][5] ,
         \register[20][4] , \register[20][3] , \register[20][2] ,
         \register[20][1] , \register[20][0] , \register[19][31] ,
         \register[19][30] , \register[19][29] , \register[19][28] ,
         \register[19][27] , \register[19][26] , \register[19][25] ,
         \register[19][24] , \register[19][23] , \register[19][22] ,
         \register[19][21] , \register[19][20] , \register[19][19] ,
         \register[19][18] , \register[19][17] , \register[19][16] ,
         \register[19][15] , \register[19][14] , \register[19][13] ,
         \register[19][12] , \register[19][11] , \register[19][10] ,
         \register[19][9] , \register[19][8] , \register[19][7] ,
         \register[19][6] , \register[19][5] , \register[19][4] ,
         \register[19][3] , \register[19][2] , \register[19][1] ,
         \register[19][0] , \register[18][31] , \register[18][30] ,
         \register[18][29] , \register[18][28] , \register[18][27] ,
         \register[18][26] , \register[18][25] , \register[18][24] ,
         \register[18][23] , \register[18][22] , \register[18][21] ,
         \register[18][20] , \register[18][19] , \register[18][18] ,
         \register[18][17] , \register[18][16] , \register[18][15] ,
         \register[18][14] , \register[18][13] , \register[18][12] ,
         \register[18][11] , \register[18][10] , \register[18][9] ,
         \register[18][8] , \register[18][7] , \register[18][6] ,
         \register[18][5] , \register[18][4] , \register[18][3] ,
         \register[18][2] , \register[18][1] , \register[18][0] ,
         \register[17][31] , \register[17][30] , \register[17][29] ,
         \register[17][28] , \register[17][27] , \register[17][26] ,
         \register[17][25] , \register[17][24] , \register[17][23] ,
         \register[17][22] , \register[17][21] , \register[17][20] ,
         \register[17][19] , \register[17][18] , \register[17][17] ,
         \register[17][16] , \register[17][15] , \register[17][14] ,
         \register[17][13] , \register[17][12] , \register[17][11] ,
         \register[17][10] , \register[17][9] , \register[17][8] ,
         \register[17][7] , \register[17][6] , \register[17][5] ,
         \register[17][4] , \register[17][3] , \register[17][2] ,
         \register[17][1] , \register[17][0] , \register[16][31] ,
         \register[16][30] , \register[16][29] , \register[16][28] ,
         \register[16][27] , \register[16][26] , \register[16][25] ,
         \register[16][24] , \register[16][23] , \register[16][22] ,
         \register[16][21] , \register[16][20] , \register[16][19] ,
         \register[16][18] , \register[16][17] , \register[16][16] ,
         \register[16][15] , \register[16][14] , \register[16][13] ,
         \register[16][12] , \register[16][11] , \register[16][10] ,
         \register[16][9] , \register[16][8] , \register[16][7] ,
         \register[16][6] , \register[16][5] , \register[16][4] ,
         \register[16][3] , \register[16][2] , \register[16][1] ,
         \register[16][0] , \register[15][31] , \register[15][30] ,
         \register[15][29] , \register[15][28] , \register[15][27] ,
         \register[15][26] , \register[15][25] , \register[15][24] ,
         \register[15][23] , \register[15][22] , \register[15][21] ,
         \register[15][20] , \register[15][19] , \register[15][18] ,
         \register[15][17] , \register[15][16] , \register[15][15] ,
         \register[15][14] , \register[15][13] , \register[15][12] ,
         \register[15][11] , \register[15][10] , \register[15][9] ,
         \register[15][8] , \register[15][7] , \register[15][6] ,
         \register[15][5] , \register[15][4] , \register[15][3] ,
         \register[15][2] , \register[15][1] , \register[15][0] ,
         \register[14][31] , \register[14][30] , \register[14][29] ,
         \register[14][28] , \register[14][27] , \register[14][26] ,
         \register[14][25] , \register[14][24] , \register[14][23] ,
         \register[14][22] , \register[14][21] , \register[14][20] ,
         \register[14][19] , \register[14][18] , \register[14][17] ,
         \register[14][16] , \register[14][15] , \register[14][14] ,
         \register[14][13] , \register[14][12] , \register[14][11] ,
         \register[14][10] , \register[14][9] , \register[14][8] ,
         \register[14][7] , \register[14][6] , \register[14][5] ,
         \register[14][4] , \register[14][3] , \register[14][2] ,
         \register[14][1] , \register[14][0] , \register[13][31] ,
         \register[13][30] , \register[13][29] , \register[13][28] ,
         \register[13][27] , \register[13][26] , \register[13][25] ,
         \register[13][24] , \register[13][23] , \register[13][22] ,
         \register[13][21] , \register[13][20] , \register[13][19] ,
         \register[13][18] , \register[13][17] , \register[13][16] ,
         \register[13][15] , \register[13][14] , \register[13][13] ,
         \register[13][12] , \register[13][11] , \register[13][10] ,
         \register[13][9] , \register[13][8] , \register[13][7] ,
         \register[13][6] , \register[13][5] , \register[13][4] ,
         \register[13][3] , \register[13][2] , \register[13][1] ,
         \register[13][0] , \register[12][31] , \register[12][30] ,
         \register[12][29] , \register[12][28] , \register[12][27] ,
         \register[12][26] , \register[12][25] , \register[12][24] ,
         \register[12][23] , \register[12][22] , \register[12][21] ,
         \register[12][20] , \register[12][19] , \register[12][18] ,
         \register[12][17] , \register[12][16] , \register[12][15] ,
         \register[12][14] , \register[12][13] , \register[12][12] ,
         \register[12][11] , \register[12][10] , \register[12][9] ,
         \register[12][8] , \register[12][7] , \register[12][6] ,
         \register[12][5] , \register[12][4] , \register[12][3] ,
         \register[12][2] , \register[12][1] , \register[12][0] ,
         \register[11][31] , \register[11][30] , \register[11][29] ,
         \register[11][28] , \register[11][27] , \register[11][26] ,
         \register[11][25] , \register[11][24] , \register[11][23] ,
         \register[11][22] , \register[11][21] , \register[11][20] ,
         \register[11][19] , \register[11][18] , \register[11][17] ,
         \register[11][16] , \register[11][15] , \register[11][14] ,
         \register[11][13] , \register[11][12] , \register[11][11] ,
         \register[11][10] , \register[11][9] , \register[11][8] ,
         \register[11][7] , \register[11][6] , \register[11][5] ,
         \register[11][4] , \register[11][3] , \register[11][2] ,
         \register[11][1] , \register[11][0] , \register[10][31] ,
         \register[10][30] , \register[10][29] , \register[10][28] ,
         \register[10][27] , \register[10][26] , \register[10][25] ,
         \register[10][24] , \register[10][23] , \register[10][22] ,
         \register[10][21] , \register[10][20] , \register[10][19] ,
         \register[10][18] , \register[10][17] , \register[10][16] ,
         \register[10][15] , \register[10][14] , \register[10][13] ,
         \register[10][12] , \register[10][11] , \register[10][10] ,
         \register[10][9] , \register[10][8] , \register[10][7] ,
         \register[10][6] , \register[10][5] , \register[10][4] ,
         \register[10][3] , \register[10][2] , \register[10][1] ,
         \register[10][0] , \register[9][31] , \register[9][30] ,
         \register[9][29] , \register[9][28] , \register[9][27] ,
         \register[9][26] , \register[9][25] , \register[9][24] ,
         \register[9][23] , \register[9][22] , \register[9][21] ,
         \register[9][20] , \register[9][19] , \register[9][18] ,
         \register[9][17] , \register[9][16] , \register[9][15] ,
         \register[9][14] , \register[9][13] , \register[9][12] ,
         \register[9][11] , \register[9][10] , \register[9][9] ,
         \register[9][8] , \register[9][7] , \register[9][6] ,
         \register[9][5] , \register[9][4] , \register[9][3] ,
         \register[9][2] , \register[9][1] , \register[9][0] ,
         \register[8][31] , \register[8][30] , \register[8][29] ,
         \register[8][28] , \register[8][27] , \register[8][26] ,
         \register[8][25] , \register[8][24] , \register[8][23] ,
         \register[8][22] , \register[8][21] , \register[8][20] ,
         \register[8][19] , \register[8][18] , \register[8][17] ,
         \register[8][16] , \register[8][15] , \register[8][14] ,
         \register[8][13] , \register[8][12] , \register[8][11] ,
         \register[8][10] , \register[8][9] , \register[8][8] ,
         \register[8][7] , \register[8][6] , \register[8][5] ,
         \register[8][4] , \register[8][3] , \register[8][2] ,
         \register[8][1] , \register[8][0] , \register[7][31] ,
         \register[7][30] , \register[7][29] , \register[7][28] ,
         \register[7][27] , \register[7][26] , \register[7][25] ,
         \register[7][24] , \register[7][23] , \register[7][22] ,
         \register[7][21] , \register[7][20] , \register[7][19] ,
         \register[7][18] , \register[7][17] , \register[7][16] ,
         \register[7][15] , \register[7][14] , \register[7][13] ,
         \register[7][12] , \register[7][11] , \register[7][10] ,
         \register[7][9] , \register[7][8] , \register[7][7] ,
         \register[7][6] , \register[7][5] , \register[7][4] ,
         \register[7][3] , \register[7][2] , \register[7][1] ,
         \register[7][0] , \register[6][31] , \register[6][30] ,
         \register[6][29] , \register[6][28] , \register[6][27] ,
         \register[6][26] , \register[6][25] , \register[6][24] ,
         \register[6][23] , \register[6][22] , \register[6][21] ,
         \register[6][20] , \register[6][19] , \register[6][18] ,
         \register[6][17] , \register[6][16] , \register[6][15] ,
         \register[6][14] , \register[6][13] , \register[6][12] ,
         \register[6][11] , \register[6][10] , \register[6][9] ,
         \register[6][8] , \register[6][7] , \register[6][6] ,
         \register[6][5] , \register[6][4] , \register[6][3] ,
         \register[6][2] , \register[6][1] , \register[6][0] ,
         \register[5][31] , \register[5][30] , \register[5][29] ,
         \register[5][28] , \register[5][27] , \register[5][26] ,
         \register[5][25] , \register[5][24] , \register[5][23] ,
         \register[5][22] , \register[5][21] , \register[5][20] ,
         \register[5][19] , \register[5][18] , \register[5][17] ,
         \register[5][16] , \register[5][15] , \register[5][14] ,
         \register[5][13] , \register[5][12] , \register[5][11] ,
         \register[5][10] , \register[5][9] , \register[5][8] ,
         \register[5][7] , \register[5][6] , \register[5][5] ,
         \register[5][4] , \register[5][3] , \register[5][2] ,
         \register[5][1] , \register[5][0] , \register[4][31] ,
         \register[4][30] , \register[4][29] , \register[4][28] ,
         \register[4][27] , \register[4][26] , \register[4][25] ,
         \register[4][24] , \register[4][23] , \register[4][22] ,
         \register[4][21] , \register[4][20] , \register[4][19] ,
         \register[4][18] , \register[4][17] , \register[4][16] ,
         \register[4][15] , \register[4][14] , \register[4][13] ,
         \register[4][12] , \register[4][11] , \register[4][10] ,
         \register[4][9] , \register[4][8] , \register[4][7] ,
         \register[4][6] , \register[4][5] , \register[4][4] ,
         \register[4][3] , \register[4][2] , \register[4][1] ,
         \register[4][0] , \register[3][31] , \register[3][30] ,
         \register[3][29] , \register[3][28] , \register[3][27] ,
         \register[3][26] , \register[3][25] , \register[3][24] ,
         \register[3][23] , \register[3][22] , \register[3][21] ,
         \register[3][20] , \register[3][19] , \register[3][18] ,
         \register[3][17] , \register[3][16] , \register[3][15] ,
         \register[3][14] , \register[3][13] , \register[3][12] ,
         \register[3][11] , \register[3][10] , \register[3][9] ,
         \register[3][8] , \register[3][7] , \register[3][6] ,
         \register[3][5] , \register[3][4] , \register[3][3] ,
         \register[3][2] , \register[3][1] , \register[3][0] ,
         \register[2][31] , \register[2][30] , \register[2][29] ,
         \register[2][28] , \register[2][27] , \register[2][26] ,
         \register[2][25] , \register[2][24] , \register[2][23] ,
         \register[2][22] , \register[2][21] , \register[2][20] ,
         \register[2][19] , \register[2][18] , \register[2][17] ,
         \register[2][16] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[1][31] ,
         \register[1][30] , \register[1][29] , \register[1][28] ,
         \register[1][27] , \register[1][26] , \register[1][25] ,
         \register[1][24] , \register[1][23] , \register[1][22] ,
         \register[1][21] , \register[1][20] , \register[1][19] ,
         \register[1][18] , \register[1][17] , \register[1][16] ,
         \register[1][15] , \register[1][14] , \register[1][13] ,
         \register[1][12] , \register[1][11] , \register[1][10] ,
         \register[1][9] , \register[1][8] , \register[1][7] ,
         \register[1][6] , \register[1][5] , \register[1][4] ,
         \register[1][3] , \register[1][2] , \register[1][1] ,
         \register[1][0] , N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n66, n67, n69, n71, n73, n75, n77, n79, n81, n82, n91, n100,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n65, n68, n70, n72, n74, n76, n78, n80, n83, n84,
         n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99,
         n101, n102, n103, n104, n105, n106, n107, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455;
  assign N12 = rsel1[0];
  assign N13 = rsel1[1];
  assign N14 = rsel1[2];
  assign N15 = rsel1[3];
  assign N16 = rsel1[4];
  assign N17 = rsel2[0];
  assign N18 = rsel2[1];
  assign N19 = rsel2[2];
  assign N20 = rsel2[3];
  assign N21 = rsel2[4];

  DFFRX1 \register_reg[2][31]  ( .D(n171), .CK(clk), .RN(n2279), .Q(
        \register[2][31] ), .QN(n2417) );
  DFFRX1 \register_reg[2][30]  ( .D(n170), .CK(clk), .RN(n2279), .Q(
        \register[2][30] ), .QN(n2416) );
  DFFRX1 \register_reg[2][29]  ( .D(n169), .CK(clk), .RN(n2279), .Q(
        \register[2][29] ), .QN(n2415) );
  DFFRX1 \register_reg[2][28]  ( .D(n168), .CK(clk), .RN(n2279), .Q(
        \register[2][28] ), .QN(n2414) );
  DFFRX1 \register_reg[2][27]  ( .D(n167), .CK(clk), .RN(n2278), .Q(
        \register[2][27] ), .QN(n2413) );
  DFFRX1 \register_reg[2][26]  ( .D(n166), .CK(clk), .RN(n2278), .Q(
        \register[2][26] ), .QN(n2412) );
  DFFRX1 \register_reg[2][25]  ( .D(n165), .CK(clk), .RN(n2278), .Q(
        \register[2][25] ), .QN(n2411) );
  DFFRX1 \register_reg[2][24]  ( .D(n164), .CK(clk), .RN(n2278), .Q(
        \register[2][24] ), .QN(n2410) );
  DFFRX1 \register_reg[2][23]  ( .D(n163), .CK(clk), .RN(n2278), .Q(
        \register[2][23] ), .QN(n2409) );
  DFFRX1 \register_reg[2][22]  ( .D(n162), .CK(clk), .RN(n2278), .Q(
        \register[2][22] ), .QN(n2408) );
  DFFRX1 \register_reg[2][21]  ( .D(n161), .CK(clk), .RN(n2278), .Q(
        \register[2][21] ), .QN(n2407) );
  DFFRX1 \register_reg[2][20]  ( .D(n160), .CK(clk), .RN(n2278), .Q(
        \register[2][20] ), .QN(n2406) );
  DFFRX1 \register_reg[2][19]  ( .D(n159), .CK(clk), .RN(n2278), .Q(
        \register[2][19] ), .QN(n2405) );
  DFFRX1 \register_reg[2][18]  ( .D(n158), .CK(clk), .RN(n2278), .Q(
        \register[2][18] ), .QN(n2404) );
  DFFRX1 \register_reg[2][17]  ( .D(n157), .CK(clk), .RN(n2278), .Q(
        \register[2][17] ), .QN(n2403) );
  DFFRX1 \register_reg[2][16]  ( .D(n156), .CK(clk), .RN(n2278), .Q(
        \register[2][16] ), .QN(n2402) );
  DFFRX1 \register_reg[2][15]  ( .D(n155), .CK(clk), .RN(n2277), .Q(
        \register[2][15] ), .QN(n2401) );
  DFFRX1 \register_reg[2][14]  ( .D(n154), .CK(clk), .RN(n2277), .Q(
        \register[2][14] ), .QN(n2400) );
  DFFRX1 \register_reg[2][13]  ( .D(n153), .CK(clk), .RN(n2277), .Q(
        \register[2][13] ), .QN(n2399) );
  DFFRX1 \register_reg[2][12]  ( .D(n152), .CK(clk), .RN(n2277), .Q(
        \register[2][12] ), .QN(n2398) );
  DFFRX1 \register_reg[2][11]  ( .D(n151), .CK(clk), .RN(n2277), .Q(
        \register[2][11] ), .QN(n2397) );
  DFFRX1 \register_reg[2][10]  ( .D(n150), .CK(clk), .RN(n2277), .Q(
        \register[2][10] ), .QN(n2396) );
  DFFRX1 \register_reg[2][9]  ( .D(n149), .CK(clk), .RN(n2277), .Q(
        \register[2][9] ), .QN(n2395) );
  DFFRX1 \register_reg[2][8]  ( .D(n148), .CK(clk), .RN(n2277), .Q(
        \register[2][8] ), .QN(n2394) );
  DFFRX1 \register_reg[2][7]  ( .D(n147), .CK(clk), .RN(n2277), .Q(
        \register[2][7] ), .QN(n2393) );
  DFFRX1 \register_reg[2][6]  ( .D(n146), .CK(clk), .RN(n2277), .Q(
        \register[2][6] ), .QN(n2392) );
  DFFRX1 \register_reg[2][5]  ( .D(n145), .CK(clk), .RN(n2277), .Q(
        \register[2][5] ), .QN(n2391) );
  DFFRX1 \register_reg[2][4]  ( .D(n144), .CK(clk), .RN(n2277), .Q(
        \register[2][4] ), .QN(n2390) );
  DFFRX1 \register_reg[2][3]  ( .D(n143), .CK(clk), .RN(n2276), .Q(
        \register[2][3] ), .QN(n2389) );
  DFFRX1 \register_reg[2][2]  ( .D(n142), .CK(clk), .RN(n2276), .Q(
        \register[2][2] ), .QN(n2388) );
  DFFRX1 \register_reg[2][1]  ( .D(n141), .CK(clk), .RN(n2276), .Q(
        \register[2][1] ), .QN(n2387) );
  DFFRX1 \register_reg[2][0]  ( .D(n140), .CK(clk), .RN(n2276), .Q(
        \register[2][0] ), .QN(n2386) );
  DFFRX1 \register_reg[31][31]  ( .D(n1099), .CK(clk), .RN(n2356), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n1098), .CK(clk), .RN(n2356), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n1097), .CK(clk), .RN(n2356), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n1096), .CK(clk), .RN(n2356), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n1095), .CK(clk), .RN(n2356), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n1094), .CK(clk), .RN(n2356), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n1093), .CK(clk), .RN(n2356), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n1092), .CK(clk), .RN(n2356), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n1091), .CK(clk), .RN(n2355), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n1090), .CK(clk), .RN(n2355), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n1089), .CK(clk), .RN(n2355), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n1088), .CK(clk), .RN(n2355), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n1087), .CK(clk), .RN(n2355), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n1086), .CK(clk), .RN(n2355), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n1085), .CK(clk), .RN(n2355), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n1084), .CK(clk), .RN(n2355), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n1083), .CK(clk), .RN(n2355), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n1082), .CK(clk), .RN(n2355), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n1081), .CK(clk), .RN(n2355), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n1080), .CK(clk), .RN(n2355), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n1079), .CK(clk), .RN(n2354), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n1078), .CK(clk), .RN(n2354), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n1077), .CK(clk), .RN(n2354), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n1076), .CK(clk), .RN(n2354), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n1075), .CK(clk), .RN(n2354), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n1074), .CK(clk), .RN(n2354), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n1073), .CK(clk), .RN(n2354), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n1072), .CK(clk), .RN(n2354), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n1071), .CK(clk), .RN(n2354), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n1070), .CK(clk), .RN(n2354), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n1069), .CK(clk), .RN(n2354), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n1068), .CK(clk), .RN(n2354), .Q(
        \register[31][0] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n971), .CK(clk), .RN(n2345), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n970), .CK(clk), .RN(n2345), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n969), .CK(clk), .RN(n2345), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n968), .CK(clk), .RN(n2345), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n967), .CK(clk), .RN(n2345), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n966), .CK(clk), .RN(n2345), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n965), .CK(clk), .RN(n2345), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n964), .CK(clk), .RN(n2345), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n963), .CK(clk), .RN(n2345), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n962), .CK(clk), .RN(n2345), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n961), .CK(clk), .RN(n2345), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n960), .CK(clk), .RN(n2345), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n959), .CK(clk), .RN(n2344), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n958), .CK(clk), .RN(n2344), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n957), .CK(clk), .RN(n2344), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n956), .CK(clk), .RN(n2344), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n955), .CK(clk), .RN(n2344), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n954), .CK(clk), .RN(n2344), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n953), .CK(clk), .RN(n2344), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n952), .CK(clk), .RN(n2344), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n951), .CK(clk), .RN(n2344), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n950), .CK(clk), .RN(n2344), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n949), .CK(clk), .RN(n2344), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n948), .CK(clk), .RN(n2344), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n947), .CK(clk), .RN(n2343), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n946), .CK(clk), .RN(n2343), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n945), .CK(clk), .RN(n2343), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n944), .CK(clk), .RN(n2343), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n943), .CK(clk), .RN(n2343), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n942), .CK(clk), .RN(n2343), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n941), .CK(clk), .RN(n2343), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n940), .CK(clk), .RN(n2343), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n843), .CK(clk), .RN(n2335), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n842), .CK(clk), .RN(n2335), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n841), .CK(clk), .RN(n2335), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n840), .CK(clk), .RN(n2335), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n839), .CK(clk), .RN(n2334), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n838), .CK(clk), .RN(n2334), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n837), .CK(clk), .RN(n2334), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n836), .CK(clk), .RN(n2334), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n835), .CK(clk), .RN(n2334), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n834), .CK(clk), .RN(n2334), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n833), .CK(clk), .RN(n2334), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n832), .CK(clk), .RN(n2334), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n831), .CK(clk), .RN(n2334), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n830), .CK(clk), .RN(n2334), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n829), .CK(clk), .RN(n2334), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n828), .CK(clk), .RN(n2334), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n827), .CK(clk), .RN(n2333), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n826), .CK(clk), .RN(n2333), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n825), .CK(clk), .RN(n2333), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n824), .CK(clk), .RN(n2333), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n823), .CK(clk), .RN(n2333), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n822), .CK(clk), .RN(n2333), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n821), .CK(clk), .RN(n2333), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n820), .CK(clk), .RN(n2333), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n819), .CK(clk), .RN(n2333), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n818), .CK(clk), .RN(n2333), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n817), .CK(clk), .RN(n2333), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n816), .CK(clk), .RN(n2333), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n815), .CK(clk), .RN(n2332), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n814), .CK(clk), .RN(n2332), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n813), .CK(clk), .RN(n2332), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n812), .CK(clk), .RN(n2332), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n715), .CK(clk), .RN(n2324), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n714), .CK(clk), .RN(n2324), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n713), .CK(clk), .RN(n2324), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n712), .CK(clk), .RN(n2324), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n711), .CK(clk), .RN(n2324), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n710), .CK(clk), .RN(n2324), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n709), .CK(clk), .RN(n2324), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n708), .CK(clk), .RN(n2324), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n707), .CK(clk), .RN(n2323), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n706), .CK(clk), .RN(n2323), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n705), .CK(clk), .RN(n2323), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n704), .CK(clk), .RN(n2323), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n703), .CK(clk), .RN(n2323), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n702), .CK(clk), .RN(n2323), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n701), .CK(clk), .RN(n2323), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n700), .CK(clk), .RN(n2323), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n699), .CK(clk), .RN(n2323), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n698), .CK(clk), .RN(n2323), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n697), .CK(clk), .RN(n2323), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n696), .CK(clk), .RN(n2323), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n695), .CK(clk), .RN(n2322), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n694), .CK(clk), .RN(n2322), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n693), .CK(clk), .RN(n2322), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n692), .CK(clk), .RN(n2322), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n691), .CK(clk), .RN(n2322), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n690), .CK(clk), .RN(n2322), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n689), .CK(clk), .RN(n2322), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n688), .CK(clk), .RN(n2322), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n687), .CK(clk), .RN(n2322), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n686), .CK(clk), .RN(n2322), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n685), .CK(clk), .RN(n2322), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n684), .CK(clk), .RN(n2322), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n587), .CK(clk), .RN(n2313), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n586), .CK(clk), .RN(n2313), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n585), .CK(clk), .RN(n2313), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n584), .CK(clk), .RN(n2313), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n583), .CK(clk), .RN(n2313), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n582), .CK(clk), .RN(n2313), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n581), .CK(clk), .RN(n2313), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n580), .CK(clk), .RN(n2313), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n579), .CK(clk), .RN(n2313), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n578), .CK(clk), .RN(n2313), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n577), .CK(clk), .RN(n2313), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n576), .CK(clk), .RN(n2313), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n575), .CK(clk), .RN(n2312), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n574), .CK(clk), .RN(n2312), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n573), .CK(clk), .RN(n2312), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n572), .CK(clk), .RN(n2312), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n571), .CK(clk), .RN(n2312), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n570), .CK(clk), .RN(n2312), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n569), .CK(clk), .RN(n2312), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n568), .CK(clk), .RN(n2312), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n567), .CK(clk), .RN(n2312), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n566), .CK(clk), .RN(n2312), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n565), .CK(clk), .RN(n2312), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n564), .CK(clk), .RN(n2312), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n563), .CK(clk), .RN(n2311), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n562), .CK(clk), .RN(n2311), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n561), .CK(clk), .RN(n2311), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n560), .CK(clk), .RN(n2311), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n559), .CK(clk), .RN(n2311), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n558), .CK(clk), .RN(n2311), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n557), .CK(clk), .RN(n2311), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n556), .CK(clk), .RN(n2311), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n459), .CK(clk), .RN(n2303), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n458), .CK(clk), .RN(n2303), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n457), .CK(clk), .RN(n2303), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n456), .CK(clk), .RN(n2303), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n455), .CK(clk), .RN(n2302), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n454), .CK(clk), .RN(n2302), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n453), .CK(clk), .RN(n2302), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n452), .CK(clk), .RN(n2302), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n451), .CK(clk), .RN(n2302), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n450), .CK(clk), .RN(n2302), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n449), .CK(clk), .RN(n2302), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n448), .CK(clk), .RN(n2302), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n447), .CK(clk), .RN(n2302), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n446), .CK(clk), .RN(n2302), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n445), .CK(clk), .RN(n2302), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n444), .CK(clk), .RN(n2302), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n443), .CK(clk), .RN(n2301), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n442), .CK(clk), .RN(n2301), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n441), .CK(clk), .RN(n2301), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n440), .CK(clk), .RN(n2301), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n439), .CK(clk), .RN(n2301), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n438), .CK(clk), .RN(n2301), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n437), .CK(clk), .RN(n2301), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n436), .CK(clk), .RN(n2301), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n435), .CK(clk), .RN(n2301), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n434), .CK(clk), .RN(n2301), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n433), .CK(clk), .RN(n2301), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n432), .CK(clk), .RN(n2301), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n431), .CK(clk), .RN(n2300), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n430), .CK(clk), .RN(n2300), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n429), .CK(clk), .RN(n2300), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n428), .CK(clk), .RN(n2300), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n331), .CK(clk), .RN(n2292), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n330), .CK(clk), .RN(n2292), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n329), .CK(clk), .RN(n2292), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n328), .CK(clk), .RN(n2292), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n327), .CK(clk), .RN(n2292), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n326), .CK(clk), .RN(n2292), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n325), .CK(clk), .RN(n2292), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n324), .CK(clk), .RN(n2292), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n323), .CK(clk), .RN(n2291), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n322), .CK(clk), .RN(n2291), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n321), .CK(clk), .RN(n2291), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n320), .CK(clk), .RN(n2291), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n319), .CK(clk), .RN(n2291), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n318), .CK(clk), .RN(n2291), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n317), .CK(clk), .RN(n2291), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n316), .CK(clk), .RN(n2291), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n315), .CK(clk), .RN(n2291), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n314), .CK(clk), .RN(n2291), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n313), .CK(clk), .RN(n2291), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n312), .CK(clk), .RN(n2291), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n311), .CK(clk), .RN(n2290), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n310), .CK(clk), .RN(n2290), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n309), .CK(clk), .RN(n2290), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n308), .CK(clk), .RN(n2290), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n307), .CK(clk), .RN(n2290), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n306), .CK(clk), .RN(n2290), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n305), .CK(clk), .RN(n2290), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n304), .CK(clk), .RN(n2290), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n303), .CK(clk), .RN(n2290), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n302), .CK(clk), .RN(n2290), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n301), .CK(clk), .RN(n2290), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n300), .CK(clk), .RN(n2290), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n1035), .CK(clk), .RN(n2351), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n1034), .CK(clk), .RN(n2351), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n1033), .CK(clk), .RN(n2351), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n1032), .CK(clk), .RN(n2351), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n1031), .CK(clk), .RN(n2350), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n1030), .CK(clk), .RN(n2350), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n1029), .CK(clk), .RN(n2350), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n1028), .CK(clk), .RN(n2350), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n1027), .CK(clk), .RN(n2350), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n1026), .CK(clk), .RN(n2350), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n1025), .CK(clk), .RN(n2350), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n1024), .CK(clk), .RN(n2350), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n1023), .CK(clk), .RN(n2350), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n1022), .CK(clk), .RN(n2350), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n1021), .CK(clk), .RN(n2350), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n1020), .CK(clk), .RN(n2350), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n1019), .CK(clk), .RN(n2349), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n1018), .CK(clk), .RN(n2349), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n1017), .CK(clk), .RN(n2349), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n1016), .CK(clk), .RN(n2349), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n1015), .CK(clk), .RN(n2349), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n1014), .CK(clk), .RN(n2349), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n1013), .CK(clk), .RN(n2349), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n1012), .CK(clk), .RN(n2349), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n1011), .CK(clk), .RN(n2349), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n1010), .CK(clk), .RN(n2349), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n1009), .CK(clk), .RN(n2349), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n1008), .CK(clk), .RN(n2349), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n1007), .CK(clk), .RN(n2348), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n1006), .CK(clk), .RN(n2348), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n1005), .CK(clk), .RN(n2348), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n1004), .CK(clk), .RN(n2348), .Q(
        \register[29][0] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n907), .CK(clk), .RN(n2340), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n906), .CK(clk), .RN(n2340), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n905), .CK(clk), .RN(n2340), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n904), .CK(clk), .RN(n2340), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n903), .CK(clk), .RN(n2340), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n902), .CK(clk), .RN(n2340), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n901), .CK(clk), .RN(n2340), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n900), .CK(clk), .RN(n2340), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n899), .CK(clk), .RN(n2339), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n898), .CK(clk), .RN(n2339), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n897), .CK(clk), .RN(n2339), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n896), .CK(clk), .RN(n2339), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n895), .CK(clk), .RN(n2339), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n894), .CK(clk), .RN(n2339), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n893), .CK(clk), .RN(n2339), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n892), .CK(clk), .RN(n2339), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n891), .CK(clk), .RN(n2339), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n890), .CK(clk), .RN(n2339), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n889), .CK(clk), .RN(n2339), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n888), .CK(clk), .RN(n2339), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n887), .CK(clk), .RN(n2338), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n886), .CK(clk), .RN(n2338), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n885), .CK(clk), .RN(n2338), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n884), .CK(clk), .RN(n2338), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n883), .CK(clk), .RN(n2338), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n882), .CK(clk), .RN(n2338), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n881), .CK(clk), .RN(n2338), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n880), .CK(clk), .RN(n2338), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n879), .CK(clk), .RN(n2338), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n878), .CK(clk), .RN(n2338), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n877), .CK(clk), .RN(n2338), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n876), .CK(clk), .RN(n2338), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n779), .CK(clk), .RN(n2329), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n778), .CK(clk), .RN(n2329), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n777), .CK(clk), .RN(n2329), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n776), .CK(clk), .RN(n2329), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n775), .CK(clk), .RN(n2329), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n774), .CK(clk), .RN(n2329), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n773), .CK(clk), .RN(n2329), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n772), .CK(clk), .RN(n2329), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n771), .CK(clk), .RN(n2329), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n770), .CK(clk), .RN(n2329), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n769), .CK(clk), .RN(n2329), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n768), .CK(clk), .RN(n2329), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n767), .CK(clk), .RN(n2328), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n766), .CK(clk), .RN(n2328), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n765), .CK(clk), .RN(n2328), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n764), .CK(clk), .RN(n2328), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n763), .CK(clk), .RN(n2328), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n762), .CK(clk), .RN(n2328), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n761), .CK(clk), .RN(n2328), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n760), .CK(clk), .RN(n2328), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n759), .CK(clk), .RN(n2328), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n758), .CK(clk), .RN(n2328), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n757), .CK(clk), .RN(n2328), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n756), .CK(clk), .RN(n2328), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n755), .CK(clk), .RN(n2327), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n754), .CK(clk), .RN(n2327), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n753), .CK(clk), .RN(n2327), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n752), .CK(clk), .RN(n2327), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n751), .CK(clk), .RN(n2327), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n750), .CK(clk), .RN(n2327), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n749), .CK(clk), .RN(n2327), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n748), .CK(clk), .RN(n2327), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n651), .CK(clk), .RN(n2319), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n650), .CK(clk), .RN(n2319), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n649), .CK(clk), .RN(n2319), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n648), .CK(clk), .RN(n2319), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n647), .CK(clk), .RN(n2318), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n646), .CK(clk), .RN(n2318), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n645), .CK(clk), .RN(n2318), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n644), .CK(clk), .RN(n2318), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n643), .CK(clk), .RN(n2318), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n642), .CK(clk), .RN(n2318), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n641), .CK(clk), .RN(n2318), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n640), .CK(clk), .RN(n2318), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n639), .CK(clk), .RN(n2318), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n638), .CK(clk), .RN(n2318), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n637), .CK(clk), .RN(n2318), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n636), .CK(clk), .RN(n2318), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n635), .CK(clk), .RN(n2317), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n634), .CK(clk), .RN(n2317), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n633), .CK(clk), .RN(n2317), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n632), .CK(clk), .RN(n2317), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n631), .CK(clk), .RN(n2317), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n630), .CK(clk), .RN(n2317), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n629), .CK(clk), .RN(n2317), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n628), .CK(clk), .RN(n2317), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n627), .CK(clk), .RN(n2317), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n626), .CK(clk), .RN(n2317), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n625), .CK(clk), .RN(n2317), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n624), .CK(clk), .RN(n2317), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n623), .CK(clk), .RN(n2316), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n622), .CK(clk), .RN(n2316), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n621), .CK(clk), .RN(n2316), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n620), .CK(clk), .RN(n2316), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n523), .CK(clk), .RN(n2308), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n522), .CK(clk), .RN(n2308), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n521), .CK(clk), .RN(n2308), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n520), .CK(clk), .RN(n2308), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n519), .CK(clk), .RN(n2308), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n518), .CK(clk), .RN(n2308), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n517), .CK(clk), .RN(n2308), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n516), .CK(clk), .RN(n2308), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n515), .CK(clk), .RN(n2307), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n514), .CK(clk), .RN(n2307), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n513), .CK(clk), .RN(n2307), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n512), .CK(clk), .RN(n2307), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n511), .CK(clk), .RN(n2307), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n510), .CK(clk), .RN(n2307), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n509), .CK(clk), .RN(n2307), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n508), .CK(clk), .RN(n2307), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n507), .CK(clk), .RN(n2307), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n506), .CK(clk), .RN(n2307), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n505), .CK(clk), .RN(n2307), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n504), .CK(clk), .RN(n2307), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n503), .CK(clk), .RN(n2306), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n502), .CK(clk), .RN(n2306), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n501), .CK(clk), .RN(n2306), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n500), .CK(clk), .RN(n2306), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n499), .CK(clk), .RN(n2306), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n498), .CK(clk), .RN(n2306), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n497), .CK(clk), .RN(n2306), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n496), .CK(clk), .RN(n2306), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n495), .CK(clk), .RN(n2306), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n494), .CK(clk), .RN(n2306), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n493), .CK(clk), .RN(n2306), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n492), .CK(clk), .RN(n2306), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n395), .CK(clk), .RN(n2297), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n394), .CK(clk), .RN(n2297), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n393), .CK(clk), .RN(n2297), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n392), .CK(clk), .RN(n2297), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n391), .CK(clk), .RN(n2297), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n390), .CK(clk), .RN(n2297), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n389), .CK(clk), .RN(n2297), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n388), .CK(clk), .RN(n2297), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n387), .CK(clk), .RN(n2297), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n386), .CK(clk), .RN(n2297), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n385), .CK(clk), .RN(n2297), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n384), .CK(clk), .RN(n2297), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n383), .CK(clk), .RN(n2296), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n382), .CK(clk), .RN(n2296), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n381), .CK(clk), .RN(n2296), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n380), .CK(clk), .RN(n2296), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n379), .CK(clk), .RN(n2296), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n378), .CK(clk), .RN(n2296), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n377), .CK(clk), .RN(n2296), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n376), .CK(clk), .RN(n2296), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n375), .CK(clk), .RN(n2296), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n374), .CK(clk), .RN(n2296), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n373), .CK(clk), .RN(n2296), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n372), .CK(clk), .RN(n2296), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n371), .CK(clk), .RN(n2295), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n370), .CK(clk), .RN(n2295), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n369), .CK(clk), .RN(n2295), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n368), .CK(clk), .RN(n2295), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n367), .CK(clk), .RN(n2295), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n366), .CK(clk), .RN(n2295), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n365), .CK(clk), .RN(n2295), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n364), .CK(clk), .RN(n2295), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n267), .CK(clk), .RN(n2287), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n266), .CK(clk), .RN(n2287), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n265), .CK(clk), .RN(n2287), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n264), .CK(clk), .RN(n2287), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n263), .CK(clk), .RN(n2286), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n262), .CK(clk), .RN(n2286), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n261), .CK(clk), .RN(n2286), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n260), .CK(clk), .RN(n2286), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n259), .CK(clk), .RN(n2286), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n258), .CK(clk), .RN(n2286), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n257), .CK(clk), .RN(n2286), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n256), .CK(clk), .RN(n2286), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n255), .CK(clk), .RN(n2286), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n254), .CK(clk), .RN(n2286), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n253), .CK(clk), .RN(n2286), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n252), .CK(clk), .RN(n2286), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n251), .CK(clk), .RN(n2285), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n250), .CK(clk), .RN(n2285), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n249), .CK(clk), .RN(n2285), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n248), .CK(clk), .RN(n2285), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n247), .CK(clk), .RN(n2285), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n246), .CK(clk), .RN(n2285), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n245), .CK(clk), .RN(n2285), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n244), .CK(clk), .RN(n2285), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n243), .CK(clk), .RN(n2285), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n242), .CK(clk), .RN(n2285), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n241), .CK(clk), .RN(n2285), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n240), .CK(clk), .RN(n2285), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n239), .CK(clk), .RN(n2284), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n238), .CK(clk), .RN(n2284), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n237), .CK(clk), .RN(n2284), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n236), .CK(clk), .RN(n2284), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n1003), .CK(clk), .RN(n2348), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n1002), .CK(clk), .RN(n2348), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n1001), .CK(clk), .RN(n2348), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n1000), .CK(clk), .RN(n2348), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n999), .CK(clk), .RN(n2348), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n998), .CK(clk), .RN(n2348), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n997), .CK(clk), .RN(n2348), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n996), .CK(clk), .RN(n2348), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n995), .CK(clk), .RN(n2347), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n994), .CK(clk), .RN(n2347), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n993), .CK(clk), .RN(n2347), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n992), .CK(clk), .RN(n2347), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n991), .CK(clk), .RN(n2347), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n990), .CK(clk), .RN(n2347), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n989), .CK(clk), .RN(n2347), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n988), .CK(clk), .RN(n2347), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n987), .CK(clk), .RN(n2347), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n986), .CK(clk), .RN(n2347), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n985), .CK(clk), .RN(n2347), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n984), .CK(clk), .RN(n2347), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n983), .CK(clk), .RN(n2346), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n982), .CK(clk), .RN(n2346), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n981), .CK(clk), .RN(n2346), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n980), .CK(clk), .RN(n2346), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n979), .CK(clk), .RN(n2346), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n978), .CK(clk), .RN(n2346), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n977), .CK(clk), .RN(n2346), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n976), .CK(clk), .RN(n2346), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n975), .CK(clk), .RN(n2346), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n974), .CK(clk), .RN(n2346), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n973), .CK(clk), .RN(n2346), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][0]  ( .D(n972), .CK(clk), .RN(n2346), .Q(
        \register[28][0] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n875), .CK(clk), .RN(n2337), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n874), .CK(clk), .RN(n2337), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n873), .CK(clk), .RN(n2337), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n872), .CK(clk), .RN(n2337), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n871), .CK(clk), .RN(n2337), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n870), .CK(clk), .RN(n2337), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n869), .CK(clk), .RN(n2337), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n868), .CK(clk), .RN(n2337), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n867), .CK(clk), .RN(n2337), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n866), .CK(clk), .RN(n2337), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n865), .CK(clk), .RN(n2337), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n864), .CK(clk), .RN(n2337), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n863), .CK(clk), .RN(n2336), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n862), .CK(clk), .RN(n2336), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n861), .CK(clk), .RN(n2336), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n860), .CK(clk), .RN(n2336), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n859), .CK(clk), .RN(n2336), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n858), .CK(clk), .RN(n2336), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n857), .CK(clk), .RN(n2336), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n856), .CK(clk), .RN(n2336), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n855), .CK(clk), .RN(n2336), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n854), .CK(clk), .RN(n2336), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n853), .CK(clk), .RN(n2336), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n852), .CK(clk), .RN(n2336), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n851), .CK(clk), .RN(n2335), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n850), .CK(clk), .RN(n2335), .Q(
        \register[24][6] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n849), .CK(clk), .RN(n2335), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n848), .CK(clk), .RN(n2335), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n847), .CK(clk), .RN(n2335), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n846), .CK(clk), .RN(n2335), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n845), .CK(clk), .RN(n2335), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n844), .CK(clk), .RN(n2335), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n747), .CK(clk), .RN(n2327), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n746), .CK(clk), .RN(n2327), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n745), .CK(clk), .RN(n2327), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n744), .CK(clk), .RN(n2327), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n743), .CK(clk), .RN(n2326), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n742), .CK(clk), .RN(n2326), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n741), .CK(clk), .RN(n2326), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n740), .CK(clk), .RN(n2326), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n739), .CK(clk), .RN(n2326), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n738), .CK(clk), .RN(n2326), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n737), .CK(clk), .RN(n2326), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n736), .CK(clk), .RN(n2326), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n735), .CK(clk), .RN(n2326), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n734), .CK(clk), .RN(n2326), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n733), .CK(clk), .RN(n2326), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n732), .CK(clk), .RN(n2326), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n731), .CK(clk), .RN(n2325), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n730), .CK(clk), .RN(n2325), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n729), .CK(clk), .RN(n2325), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n728), .CK(clk), .RN(n2325), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n727), .CK(clk), .RN(n2325), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n726), .CK(clk), .RN(n2325), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n725), .CK(clk), .RN(n2325), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n724), .CK(clk), .RN(n2325), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n723), .CK(clk), .RN(n2325), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n722), .CK(clk), .RN(n2325), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n721), .CK(clk), .RN(n2325), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n720), .CK(clk), .RN(n2325), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n719), .CK(clk), .RN(n2324), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n718), .CK(clk), .RN(n2324), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n717), .CK(clk), .RN(n2324), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[20][0]  ( .D(n716), .CK(clk), .RN(n2324), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n619), .CK(clk), .RN(n2316), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n618), .CK(clk), .RN(n2316), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n617), .CK(clk), .RN(n2316), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n616), .CK(clk), .RN(n2316), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n615), .CK(clk), .RN(n2316), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n614), .CK(clk), .RN(n2316), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n613), .CK(clk), .RN(n2316), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n612), .CK(clk), .RN(n2316), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n611), .CK(clk), .RN(n2315), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n610), .CK(clk), .RN(n2315), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n609), .CK(clk), .RN(n2315), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n608), .CK(clk), .RN(n2315), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n607), .CK(clk), .RN(n2315), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n606), .CK(clk), .RN(n2315), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n605), .CK(clk), .RN(n2315), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n604), .CK(clk), .RN(n2315), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n603), .CK(clk), .RN(n2315), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n602), .CK(clk), .RN(n2315), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n601), .CK(clk), .RN(n2315), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n600), .CK(clk), .RN(n2315), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n599), .CK(clk), .RN(n2314), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n598), .CK(clk), .RN(n2314), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n597), .CK(clk), .RN(n2314), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n596), .CK(clk), .RN(n2314), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n595), .CK(clk), .RN(n2314), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n594), .CK(clk), .RN(n2314), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n593), .CK(clk), .RN(n2314), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n592), .CK(clk), .RN(n2314), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n591), .CK(clk), .RN(n2314), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n590), .CK(clk), .RN(n2314), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n589), .CK(clk), .RN(n2314), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n588), .CK(clk), .RN(n2314), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n491), .CK(clk), .RN(n2305), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n490), .CK(clk), .RN(n2305), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n489), .CK(clk), .RN(n2305), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n488), .CK(clk), .RN(n2305), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n487), .CK(clk), .RN(n2305), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n486), .CK(clk), .RN(n2305), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n485), .CK(clk), .RN(n2305), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n484), .CK(clk), .RN(n2305), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n483), .CK(clk), .RN(n2305), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n482), .CK(clk), .RN(n2305), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n481), .CK(clk), .RN(n2305), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n480), .CK(clk), .RN(n2305), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n479), .CK(clk), .RN(n2304), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n478), .CK(clk), .RN(n2304), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n477), .CK(clk), .RN(n2304), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n476), .CK(clk), .RN(n2304), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n475), .CK(clk), .RN(n2304), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n474), .CK(clk), .RN(n2304), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n473), .CK(clk), .RN(n2304), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n472), .CK(clk), .RN(n2304), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n471), .CK(clk), .RN(n2304), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n470), .CK(clk), .RN(n2304), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n469), .CK(clk), .RN(n2304), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n468), .CK(clk), .RN(n2304), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n467), .CK(clk), .RN(n2303), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n466), .CK(clk), .RN(n2303), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n465), .CK(clk), .RN(n2303), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n464), .CK(clk), .RN(n2303), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n463), .CK(clk), .RN(n2303), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n462), .CK(clk), .RN(n2303), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n461), .CK(clk), .RN(n2303), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n460), .CK(clk), .RN(n2303), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n363), .CK(clk), .RN(n2295), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n362), .CK(clk), .RN(n2295), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n361), .CK(clk), .RN(n2295), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n360), .CK(clk), .RN(n2295), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n359), .CK(clk), .RN(n2294), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n358), .CK(clk), .RN(n2294), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n357), .CK(clk), .RN(n2294), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n356), .CK(clk), .RN(n2294), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n355), .CK(clk), .RN(n2294), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n354), .CK(clk), .RN(n2294), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n353), .CK(clk), .RN(n2294), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n352), .CK(clk), .RN(n2294), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n351), .CK(clk), .RN(n2294), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n350), .CK(clk), .RN(n2294), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n349), .CK(clk), .RN(n2294), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n348), .CK(clk), .RN(n2294), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n347), .CK(clk), .RN(n2293), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n346), .CK(clk), .RN(n2293), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n345), .CK(clk), .RN(n2293), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n344), .CK(clk), .RN(n2293), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n343), .CK(clk), .RN(n2293), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n342), .CK(clk), .RN(n2293), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n341), .CK(clk), .RN(n2293), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n340), .CK(clk), .RN(n2293), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n339), .CK(clk), .RN(n2293), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n338), .CK(clk), .RN(n2293), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n337), .CK(clk), .RN(n2293), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n336), .CK(clk), .RN(n2293), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n335), .CK(clk), .RN(n2292), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n334), .CK(clk), .RN(n2292), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n333), .CK(clk), .RN(n2292), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n332), .CK(clk), .RN(n2292), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n235), .CK(clk), .RN(n2284), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n234), .CK(clk), .RN(n2284), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n233), .CK(clk), .RN(n2284), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n232), .CK(clk), .RN(n2284), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n231), .CK(clk), .RN(n2284), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n230), .CK(clk), .RN(n2284), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n229), .CK(clk), .RN(n2284), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n228), .CK(clk), .RN(n2284), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n227), .CK(clk), .RN(n2283), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n226), .CK(clk), .RN(n2283), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n225), .CK(clk), .RN(n2283), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n224), .CK(clk), .RN(n2283), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n223), .CK(clk), .RN(n2283), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n222), .CK(clk), .RN(n2283), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n221), .CK(clk), .RN(n2283), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n220), .CK(clk), .RN(n2283), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n219), .CK(clk), .RN(n2283), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n218), .CK(clk), .RN(n2283), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n217), .CK(clk), .RN(n2283), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n216), .CK(clk), .RN(n2283), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n215), .CK(clk), .RN(n2282), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n214), .CK(clk), .RN(n2282), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n213), .CK(clk), .RN(n2282), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n212), .CK(clk), .RN(n2282), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n211), .CK(clk), .RN(n2282), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n210), .CK(clk), .RN(n2282), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n209), .CK(clk), .RN(n2282), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n208), .CK(clk), .RN(n2282), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n207), .CK(clk), .RN(n2282), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n206), .CK(clk), .RN(n2282), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n205), .CK(clk), .RN(n2282), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n204), .CK(clk), .RN(n2282), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n1067), .CK(clk), .RN(n2353), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n1066), .CK(clk), .RN(n2353), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n1065), .CK(clk), .RN(n2353), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n1064), .CK(clk), .RN(n2353), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n1063), .CK(clk), .RN(n2353), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n1062), .CK(clk), .RN(n2353), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n1061), .CK(clk), .RN(n2353), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n1060), .CK(clk), .RN(n2353), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n1059), .CK(clk), .RN(n2353), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n1058), .CK(clk), .RN(n2353), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n1057), .CK(clk), .RN(n2353), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n1056), .CK(clk), .RN(n2353), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n1055), .CK(clk), .RN(n2352), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n1054), .CK(clk), .RN(n2352), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n1053), .CK(clk), .RN(n2352), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n1052), .CK(clk), .RN(n2352), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n1051), .CK(clk), .RN(n2352), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n1050), .CK(clk), .RN(n2352), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n1049), .CK(clk), .RN(n2352), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n1048), .CK(clk), .RN(n2352), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n1047), .CK(clk), .RN(n2352), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n1046), .CK(clk), .RN(n2352), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n1045), .CK(clk), .RN(n2352), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n1044), .CK(clk), .RN(n2352), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n1043), .CK(clk), .RN(n2351), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n1042), .CK(clk), .RN(n2351), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n1041), .CK(clk), .RN(n2351), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n1040), .CK(clk), .RN(n2351), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n1039), .CK(clk), .RN(n2351), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n1038), .CK(clk), .RN(n2351), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n1037), .CK(clk), .RN(n2351), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][0]  ( .D(n1036), .CK(clk), .RN(n2351), .Q(
        \register[30][0] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n939), .CK(clk), .RN(n2343), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n938), .CK(clk), .RN(n2343), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n937), .CK(clk), .RN(n2343), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n936), .CK(clk), .RN(n2343), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n935), .CK(clk), .RN(n2342), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n934), .CK(clk), .RN(n2342), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n933), .CK(clk), .RN(n2342), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n932), .CK(clk), .RN(n2342), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n931), .CK(clk), .RN(n2342), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n930), .CK(clk), .RN(n2342), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n929), .CK(clk), .RN(n2342), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n928), .CK(clk), .RN(n2342), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n927), .CK(clk), .RN(n2342), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n926), .CK(clk), .RN(n2342), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n925), .CK(clk), .RN(n2342), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n924), .CK(clk), .RN(n2342), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n923), .CK(clk), .RN(n2341), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n922), .CK(clk), .RN(n2341), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n921), .CK(clk), .RN(n2341), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n920), .CK(clk), .RN(n2341), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n919), .CK(clk), .RN(n2341), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n918), .CK(clk), .RN(n2341), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n917), .CK(clk), .RN(n2341), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n916), .CK(clk), .RN(n2341), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n915), .CK(clk), .RN(n2341), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n914), .CK(clk), .RN(n2341), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n913), .CK(clk), .RN(n2341), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n912), .CK(clk), .RN(n2341), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n911), .CK(clk), .RN(n2340), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n910), .CK(clk), .RN(n2340), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n909), .CK(clk), .RN(n2340), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n908), .CK(clk), .RN(n2340), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n811), .CK(clk), .RN(n2332), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n810), .CK(clk), .RN(n2332), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n809), .CK(clk), .RN(n2332), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n808), .CK(clk), .RN(n2332), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n807), .CK(clk), .RN(n2332), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n806), .CK(clk), .RN(n2332), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n805), .CK(clk), .RN(n2332), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n804), .CK(clk), .RN(n2332), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n803), .CK(clk), .RN(n2331), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n802), .CK(clk), .RN(n2331), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n801), .CK(clk), .RN(n2331), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n800), .CK(clk), .RN(n2331), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n799), .CK(clk), .RN(n2331), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n798), .CK(clk), .RN(n2331), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n797), .CK(clk), .RN(n2331), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n796), .CK(clk), .RN(n2331), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n795), .CK(clk), .RN(n2331), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n794), .CK(clk), .RN(n2331), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n793), .CK(clk), .RN(n2331), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n792), .CK(clk), .RN(n2331), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n791), .CK(clk), .RN(n2330), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n790), .CK(clk), .RN(n2330), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n789), .CK(clk), .RN(n2330), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n788), .CK(clk), .RN(n2330), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n787), .CK(clk), .RN(n2330), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n786), .CK(clk), .RN(n2330), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n785), .CK(clk), .RN(n2330), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n784), .CK(clk), .RN(n2330), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n783), .CK(clk), .RN(n2330), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n782), .CK(clk), .RN(n2330), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n781), .CK(clk), .RN(n2330), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n780), .CK(clk), .RN(n2330), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n683), .CK(clk), .RN(n2321), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n682), .CK(clk), .RN(n2321), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n681), .CK(clk), .RN(n2321), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n680), .CK(clk), .RN(n2321), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n679), .CK(clk), .RN(n2321), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n678), .CK(clk), .RN(n2321), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n677), .CK(clk), .RN(n2321), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n676), .CK(clk), .RN(n2321), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n675), .CK(clk), .RN(n2321), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n674), .CK(clk), .RN(n2321), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n673), .CK(clk), .RN(n2321), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n672), .CK(clk), .RN(n2321), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n671), .CK(clk), .RN(n2320), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n670), .CK(clk), .RN(n2320), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n669), .CK(clk), .RN(n2320), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n668), .CK(clk), .RN(n2320), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n667), .CK(clk), .RN(n2320), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n666), .CK(clk), .RN(n2320), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n665), .CK(clk), .RN(n2320), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n664), .CK(clk), .RN(n2320), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n663), .CK(clk), .RN(n2320), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n662), .CK(clk), .RN(n2320), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n661), .CK(clk), .RN(n2320), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n660), .CK(clk), .RN(n2320), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n659), .CK(clk), .RN(n2319), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n658), .CK(clk), .RN(n2319), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n657), .CK(clk), .RN(n2319), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n656), .CK(clk), .RN(n2319), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n655), .CK(clk), .RN(n2319), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n654), .CK(clk), .RN(n2319), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n653), .CK(clk), .RN(n2319), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n652), .CK(clk), .RN(n2319), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n555), .CK(clk), .RN(n2311), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n554), .CK(clk), .RN(n2311), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n553), .CK(clk), .RN(n2311), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n552), .CK(clk), .RN(n2311), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n551), .CK(clk), .RN(n2310), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n550), .CK(clk), .RN(n2310), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n549), .CK(clk), .RN(n2310), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n548), .CK(clk), .RN(n2310), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n547), .CK(clk), .RN(n2310), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n546), .CK(clk), .RN(n2310), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n545), .CK(clk), .RN(n2310), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n544), .CK(clk), .RN(n2310), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n543), .CK(clk), .RN(n2310), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n542), .CK(clk), .RN(n2310), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n541), .CK(clk), .RN(n2310), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n540), .CK(clk), .RN(n2310), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n539), .CK(clk), .RN(n2309), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n538), .CK(clk), .RN(n2309), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n537), .CK(clk), .RN(n2309), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n536), .CK(clk), .RN(n2309), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n535), .CK(clk), .RN(n2309), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n534), .CK(clk), .RN(n2309), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n533), .CK(clk), .RN(n2309), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n532), .CK(clk), .RN(n2309), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n531), .CK(clk), .RN(n2309), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n530), .CK(clk), .RN(n2309), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n529), .CK(clk), .RN(n2309), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n528), .CK(clk), .RN(n2309), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n527), .CK(clk), .RN(n2308), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n526), .CK(clk), .RN(n2308), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n525), .CK(clk), .RN(n2308), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n524), .CK(clk), .RN(n2308), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n427), .CK(clk), .RN(n2300), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n426), .CK(clk), .RN(n2300), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n425), .CK(clk), .RN(n2300), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n424), .CK(clk), .RN(n2300), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n423), .CK(clk), .RN(n2300), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n422), .CK(clk), .RN(n2300), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n421), .CK(clk), .RN(n2300), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n420), .CK(clk), .RN(n2300), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n419), .CK(clk), .RN(n2299), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n418), .CK(clk), .RN(n2299), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n417), .CK(clk), .RN(n2299), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n416), .CK(clk), .RN(n2299), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n415), .CK(clk), .RN(n2299), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n414), .CK(clk), .RN(n2299), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n413), .CK(clk), .RN(n2299), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n412), .CK(clk), .RN(n2299), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n411), .CK(clk), .RN(n2299), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n410), .CK(clk), .RN(n2299), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n409), .CK(clk), .RN(n2299), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n408), .CK(clk), .RN(n2299), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n407), .CK(clk), .RN(n2298), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n406), .CK(clk), .RN(n2298), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n405), .CK(clk), .RN(n2298), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n404), .CK(clk), .RN(n2298), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n403), .CK(clk), .RN(n2298), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n402), .CK(clk), .RN(n2298), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n401), .CK(clk), .RN(n2298), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n400), .CK(clk), .RN(n2298), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n399), .CK(clk), .RN(n2298), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n398), .CK(clk), .RN(n2298), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n397), .CK(clk), .RN(n2298), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n396), .CK(clk), .RN(n2298), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n299), .CK(clk), .RN(n2289), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n298), .CK(clk), .RN(n2289), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n297), .CK(clk), .RN(n2289), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n296), .CK(clk), .RN(n2289), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n295), .CK(clk), .RN(n2289), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n294), .CK(clk), .RN(n2289), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n293), .CK(clk), .RN(n2289), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n292), .CK(clk), .RN(n2289), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n291), .CK(clk), .RN(n2289), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n290), .CK(clk), .RN(n2289), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n289), .CK(clk), .RN(n2289), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n288), .CK(clk), .RN(n2289), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n287), .CK(clk), .RN(n2288), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n286), .CK(clk), .RN(n2288), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n285), .CK(clk), .RN(n2288), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n284), .CK(clk), .RN(n2288), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n283), .CK(clk), .RN(n2288), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n282), .CK(clk), .RN(n2288), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n281), .CK(clk), .RN(n2288), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n280), .CK(clk), .RN(n2288), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n279), .CK(clk), .RN(n2288), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n278), .CK(clk), .RN(n2288), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n277), .CK(clk), .RN(n2288), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n276), .CK(clk), .RN(n2288), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n275), .CK(clk), .RN(n2287), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n274), .CK(clk), .RN(n2287), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n273), .CK(clk), .RN(n2287), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n272), .CK(clk), .RN(n2287), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n271), .CK(clk), .RN(n2287), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n270), .CK(clk), .RN(n2287), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n269), .CK(clk), .RN(n2287), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n268), .CK(clk), .RN(n2287), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[3][31]  ( .D(n203), .CK(clk), .RN(n2281), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n202), .CK(clk), .RN(n2281), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n201), .CK(clk), .RN(n2281), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n200), .CK(clk), .RN(n2281), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n199), .CK(clk), .RN(n2281), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n198), .CK(clk), .RN(n2281), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n197), .CK(clk), .RN(n2281), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n196), .CK(clk), .RN(n2281), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n195), .CK(clk), .RN(n2281), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n194), .CK(clk), .RN(n2281), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n193), .CK(clk), .RN(n2281), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n192), .CK(clk), .RN(n2281), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n191), .CK(clk), .RN(n2280), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n190), .CK(clk), .RN(n2280), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n189), .CK(clk), .RN(n2280), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n188), .CK(clk), .RN(n2280), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n187), .CK(clk), .RN(n2280), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n186), .CK(clk), .RN(n2280), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n185), .CK(clk), .RN(n2280), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n184), .CK(clk), .RN(n2280), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n183), .CK(clk), .RN(n2280), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n182), .CK(clk), .RN(n2280), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n181), .CK(clk), .RN(n2280), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n180), .CK(clk), .RN(n2280), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n179), .CK(clk), .RN(n2279), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n178), .CK(clk), .RN(n2279), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n177), .CK(clk), .RN(n2279), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n176), .CK(clk), .RN(n2279), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n175), .CK(clk), .RN(n2279), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n174), .CK(clk), .RN(n2279), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n173), .CK(clk), .RN(n2279), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n172), .CK(clk), .RN(n2279), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n139), .CK(clk), .RN(n2276), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n138), .CK(clk), .RN(n2276), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n137), .CK(clk), .RN(n2276), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n136), .CK(clk), .RN(n2276), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n135), .CK(clk), .RN(n2276), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n134), .CK(clk), .RN(n2276), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n133), .CK(clk), .RN(n2276), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n132), .CK(clk), .RN(n2276), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n131), .CK(clk), .RN(n2275), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n130), .CK(clk), .RN(n2275), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n129), .CK(clk), .RN(n2275), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n128), .CK(clk), .RN(n2275), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n127), .CK(clk), .RN(n2275), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n126), .CK(clk), .RN(n2275), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n125), .CK(clk), .RN(n2275), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n124), .CK(clk), .RN(n2275), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n123), .CK(clk), .RN(n2275), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n122), .CK(clk), .RN(n2275), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n121), .CK(clk), .RN(n2275), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n120), .CK(clk), .RN(n2275), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n119), .CK(clk), .RN(n2274), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n118), .CK(clk), .RN(n2274), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n117), .CK(clk), .RN(n2274), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n116), .CK(clk), .RN(n2274), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n115), .CK(clk), .RN(n2274), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n114), .CK(clk), .RN(n2274), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n113), .CK(clk), .RN(n2274), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n112), .CK(clk), .RN(n2274), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n111), .CK(clk), .RN(n2274), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n110), .CK(clk), .RN(n2274), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][1]  ( .D(n109), .CK(clk), .RN(n2274), .Q(
        \register[1][1] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n108), .CK(clk), .RN(n2274), .Q(
        \register[1][0] ) );
  NOR3X1 U3 ( .A(wsel[0]), .B(wsel[1]), .C(n2452), .Y(n73) );
  NOR3X1 U4 ( .A(n2454), .B(wsel[1]), .C(n2452), .Y(n75) );
  NOR3X2 U5 ( .A(n2451), .B(wsel[4]), .C(n2455), .Y(n81) );
  NOR3X2 U6 ( .A(n2450), .B(wsel[3]), .C(n2455), .Y(n91) );
  NOR3X1 U7 ( .A(n2454), .B(wsel[2]), .C(n2453), .Y(n71) );
  NOR3X1 U8 ( .A(wsel[0]), .B(wsel[2]), .C(n2453), .Y(n69) );
  NOR3X2 U9 ( .A(wsel[3]), .B(wsel[4]), .C(n2455), .Y(n67) );
  NAND2X1 U10 ( .A(n100), .B(n66), .Y(n1) );
  NAND2X1 U11 ( .A(n100), .B(n82), .Y(n2) );
  NAND2X1 U12 ( .A(n100), .B(n69), .Y(n3) );
  NAND2X1 U13 ( .A(n100), .B(n71), .Y(n4) );
  NAND2X1 U14 ( .A(n100), .B(n73), .Y(n5) );
  NAND2X1 U15 ( .A(n100), .B(n75), .Y(n6) );
  NAND2X1 U16 ( .A(n100), .B(n77), .Y(n7) );
  NAND2X1 U17 ( .A(n100), .B(n79), .Y(n8) );
  NAND2X1 U18 ( .A(n81), .B(n66), .Y(n9) );
  NAND2X1 U19 ( .A(n91), .B(n66), .Y(n10) );
  NAND2X1 U20 ( .A(n66), .B(n67), .Y(n11) );
  NAND2X1 U21 ( .A(n81), .B(n82), .Y(n12) );
  NAND2X1 U22 ( .A(n81), .B(n69), .Y(n13) );
  NAND2X1 U23 ( .A(n81), .B(n71), .Y(n14) );
  NAND2X1 U24 ( .A(n81), .B(n73), .Y(n15) );
  NAND2X1 U25 ( .A(n81), .B(n75), .Y(n16) );
  NAND2X1 U26 ( .A(n81), .B(n77), .Y(n17) );
  NAND2X1 U27 ( .A(n81), .B(n79), .Y(n18) );
  NAND2X1 U28 ( .A(n91), .B(n82), .Y(n19) );
  NAND2X1 U29 ( .A(n91), .B(n69), .Y(n20) );
  NAND2X1 U30 ( .A(n91), .B(n71), .Y(n21) );
  NAND2X1 U31 ( .A(n91), .B(n73), .Y(n22) );
  NAND2X1 U32 ( .A(n91), .B(n75), .Y(n23) );
  NAND2X1 U33 ( .A(n91), .B(n77), .Y(n24) );
  NAND2X1 U34 ( .A(n91), .B(n79), .Y(n25) );
  NAND2X1 U35 ( .A(n69), .B(n67), .Y(n26) );
  NAND2X1 U36 ( .A(n71), .B(n67), .Y(n27) );
  NAND2X1 U37 ( .A(n73), .B(n67), .Y(n28) );
  NAND2X1 U38 ( .A(n75), .B(n67), .Y(n29) );
  NAND2X1 U39 ( .A(n77), .B(n67), .Y(n30) );
  NAND2X1 U40 ( .A(n79), .B(n67), .Y(n31) );
  CLKBUFX3 U41 ( .A(n1560), .Y(n1578) );
  CLKBUFX3 U42 ( .A(n2085), .Y(n2103) );
  CLKBUFX3 U43 ( .A(n2084), .Y(n2104) );
  CLKBUFX3 U44 ( .A(n1561), .Y(n1579) );
  CLKBUFX3 U45 ( .A(n1561), .Y(n1580) );
  CLKBUFX2 U46 ( .A(rst_n), .Y(n2273) );
  CLKBUFX2 U47 ( .A(rst_n), .Y(n2272) );
  CLKBUFX2 U48 ( .A(N17), .Y(n2268) );
  CLKBUFX2 U49 ( .A(N20), .Y(n2269) );
  NOR3X1 U50 ( .A(n2453), .B(n2454), .C(n2452), .Y(n79) );
  INVXL U51 ( .A(wdata[1]), .Y(n2448) );
  INVXL U52 ( .A(wdata[5]), .Y(n2444) );
  INVXL U53 ( .A(wdata[6]), .Y(n2443) );
  INVXL U54 ( .A(wdata[2]), .Y(n2447) );
  INVXL U55 ( .A(wdata[31]), .Y(n2418) );
  INVXL U56 ( .A(wdata[12]), .Y(n2437) );
  INVXL U57 ( .A(wdata[19]), .Y(n2430) );
  INVXL U58 ( .A(wdata[27]), .Y(n2422) );
  INVXL U59 ( .A(wdata[3]), .Y(n2446) );
  INVXL U60 ( .A(wdata[7]), .Y(n2442) );
  INVXL U61 ( .A(wdata[18]), .Y(n2431) );
  INVXL U62 ( .A(wdata[0]), .Y(n2449) );
  INVXL U63 ( .A(wdata[9]), .Y(n2440) );
  INVXL U64 ( .A(wdata[11]), .Y(n2438) );
  INVXL U65 ( .A(wdata[23]), .Y(n2426) );
  INVXL U66 ( .A(wdata[24]), .Y(n2425) );
  CLKINVX1 U67 ( .A(wdata[10]), .Y(n2439) );
  INVXL U68 ( .A(wdata[21]), .Y(n2428) );
  CLKINVX1 U69 ( .A(wdata[25]), .Y(n2424) );
  INVXL U70 ( .A(wdata[4]), .Y(n2445) );
  INVXL U71 ( .A(wdata[29]), .Y(n2420) );
  INVXL U72 ( .A(wdata[15]), .Y(n2434) );
  INVXL U73 ( .A(wdata[8]), .Y(n2441) );
  INVXL U74 ( .A(wdata[13]), .Y(n2436) );
  INVXL U75 ( .A(wdata[14]), .Y(n2435) );
  INVXL U76 ( .A(wdata[17]), .Y(n2432) );
  INVXL U77 ( .A(wdata[22]), .Y(n2427) );
  INVXL U78 ( .A(wdata[26]), .Y(n2423) );
  INVXL U79 ( .A(wdata[28]), .Y(n2421) );
  INVXL U80 ( .A(wdata[30]), .Y(n2419) );
  INVXL U81 ( .A(wdata[16]), .Y(n2433) );
  INVXL U82 ( .A(wdata[20]), .Y(n2429) );
  INVX1 U83 ( .A(wsel[4]), .Y(n2450) );
  XNOR2XL U84 ( .A(n2268), .B(wsel[0]), .Y(n49) );
  XNOR2XL U85 ( .A(N12), .B(wsel[0]), .Y(n58) );
  NOR3X1 U86 ( .A(n2453), .B(wsel[0]), .C(n2452), .Y(n77) );
  INVX1 U87 ( .A(wsel[3]), .Y(n2451) );
  INVX1 U88 ( .A(wsel[2]), .Y(n2452) );
  INVX1 U89 ( .A(wsel[1]), .Y(n2453) );
  INVX1 U90 ( .A(wsel[0]), .Y(n2454) );
  CLKINVX2 U91 ( .A(wen), .Y(n2455) );
  NOR2X1 U92 ( .A(n2082), .B(n2268), .Y(n1977) );
  NOR2X1 U93 ( .A(n2082), .B(n2098), .Y(n1972) );
  NOR2X1 U94 ( .A(n2082), .B(n2102), .Y(n1962) );
  NOR2X1 U95 ( .A(n2083), .B(n2095), .Y(n1957) );
  NOR2X1 U96 ( .A(n2083), .B(n2102), .Y(n1952) );
  NOR2X1 U97 ( .A(n2083), .B(n2102), .Y(n1947) );
  NOR2X1 U98 ( .A(n2083), .B(n2102), .Y(n1942) );
  NOR2X1 U99 ( .A(n2083), .B(n2102), .Y(n1937) );
  NOR2X1 U100 ( .A(n1556), .B(n1578), .Y(n1450) );
  NOR2X1 U101 ( .A(n1556), .B(n1578), .Y(n1445) );
  NOR2X1 U102 ( .A(n1556), .B(n1578), .Y(n1435) );
  NOR2X1 U103 ( .A(n1557), .B(n1578), .Y(n1430) );
  NOR2X1 U104 ( .A(n1557), .B(n1578), .Y(n1425) );
  NOR2X1 U105 ( .A(n1557), .B(n1578), .Y(n1420) );
  NOR2X1 U106 ( .A(n1557), .B(n1578), .Y(n1415) );
  NOR2X1 U107 ( .A(n1557), .B(n1578), .Y(n1410) );
  NOR2X1 U108 ( .A(N18), .B(n2104), .Y(n2057) );
  NOR2X1 U109 ( .A(N18), .B(n2104), .Y(n2032) );
  NOR2X1 U110 ( .A(n1553), .B(n1580), .Y(n1530) );
  NOR2X1 U111 ( .A(n1553), .B(n1580), .Y(n1505) );
  NOR2X1 U112 ( .A(n2081), .B(n2104), .Y(n2052) );
  NOR2X1 U113 ( .A(n2080), .B(n2104), .Y(n2047) );
  NOR2X1 U114 ( .A(n2080), .B(n2104), .Y(n2042) );
  NOR2X1 U115 ( .A(n2080), .B(n2104), .Y(n2037) );
  NOR2X1 U116 ( .A(n2081), .B(n2104), .Y(n2027) );
  NOR2X1 U117 ( .A(n2080), .B(n2104), .Y(n2022) );
  NOR2X1 U118 ( .A(n2080), .B(n2103), .Y(n2017) );
  NOR2X1 U119 ( .A(n2080), .B(n2103), .Y(n2012) );
  NOR2X1 U120 ( .A(n2080), .B(n2103), .Y(n2007) );
  NOR2X1 U121 ( .A(n2081), .B(n2103), .Y(n2002) );
  NOR2X1 U122 ( .A(n2081), .B(n2103), .Y(n1997) );
  NOR2X1 U123 ( .A(n2081), .B(n2103), .Y(n1992) );
  NOR2X1 U124 ( .A(n2082), .B(n2103), .Y(n1987) );
  NOR2X1 U125 ( .A(n2082), .B(n2103), .Y(n1982) );
  NOR2X1 U126 ( .A(n2082), .B(n2103), .Y(n1967) );
  NOR2X1 U127 ( .A(n2083), .B(n2103), .Y(n1932) );
  NOR2X1 U128 ( .A(n1555), .B(n1580), .Y(n1525) );
  NOR2X1 U129 ( .A(n1554), .B(n1580), .Y(n1520) );
  NOR2X1 U130 ( .A(n1554), .B(n1580), .Y(n1515) );
  NOR2X1 U131 ( .A(n1554), .B(n1580), .Y(n1510) );
  NOR2X1 U132 ( .A(n1555), .B(n1580), .Y(n1500) );
  NOR2X1 U133 ( .A(n1554), .B(n1580), .Y(n1495) );
  NOR2X1 U134 ( .A(n1554), .B(n1579), .Y(n1490) );
  NOR2X1 U135 ( .A(n1554), .B(n1579), .Y(n1485) );
  NOR2X1 U136 ( .A(n1554), .B(n1579), .Y(n1480) );
  NOR2X1 U137 ( .A(n1555), .B(n1579), .Y(n1475) );
  NOR2X1 U138 ( .A(n1555), .B(n1579), .Y(n1470) );
  NOR2X1 U139 ( .A(n1555), .B(n1579), .Y(n1465) );
  NOR2X1 U140 ( .A(n1556), .B(n1579), .Y(n1460) );
  NOR2X1 U141 ( .A(n1556), .B(n1579), .Y(n1455) );
  NOR2X1 U142 ( .A(n1556), .B(n1579), .Y(n1440) );
  NOR2X1 U143 ( .A(n1557), .B(n1579), .Y(n1405) );
  CLKBUFX3 U144 ( .A(n2374), .Y(n2285) );
  CLKBUFX3 U145 ( .A(n2374), .Y(n2286) );
  CLKBUFX3 U146 ( .A(n2374), .Y(n2287) );
  CLKBUFX3 U147 ( .A(n2374), .Y(n2288) );
  CLKBUFX3 U148 ( .A(n2373), .Y(n2289) );
  CLKBUFX3 U149 ( .A(n2373), .Y(n2290) );
  CLKBUFX3 U150 ( .A(n2373), .Y(n2291) );
  CLKBUFX3 U151 ( .A(n2373), .Y(n2292) );
  CLKBUFX3 U152 ( .A(n2372), .Y(n2293) );
  CLKBUFX3 U153 ( .A(n2372), .Y(n2294) );
  CLKBUFX3 U154 ( .A(n2372), .Y(n2295) );
  CLKBUFX3 U155 ( .A(n2372), .Y(n2296) );
  CLKBUFX3 U156 ( .A(n2371), .Y(n2297) );
  CLKBUFX3 U157 ( .A(n2371), .Y(n2298) );
  CLKBUFX3 U158 ( .A(n2371), .Y(n2299) );
  CLKBUFX3 U159 ( .A(n2371), .Y(n2300) );
  CLKBUFX3 U160 ( .A(n2370), .Y(n2301) );
  CLKBUFX3 U161 ( .A(n2370), .Y(n2302) );
  CLKBUFX3 U162 ( .A(n2370), .Y(n2303) );
  CLKBUFX3 U163 ( .A(n2370), .Y(n2304) );
  CLKBUFX3 U164 ( .A(n2369), .Y(n2305) );
  CLKBUFX3 U165 ( .A(n2369), .Y(n2306) );
  CLKBUFX3 U166 ( .A(n2369), .Y(n2307) );
  CLKBUFX3 U167 ( .A(n2369), .Y(n2308) );
  CLKBUFX3 U168 ( .A(n2368), .Y(n2309) );
  CLKBUFX3 U169 ( .A(n2368), .Y(n2310) );
  CLKBUFX3 U170 ( .A(n2368), .Y(n2311) );
  CLKBUFX3 U171 ( .A(n2368), .Y(n2312) );
  CLKBUFX3 U172 ( .A(n2367), .Y(n2313) );
  CLKBUFX3 U173 ( .A(n2367), .Y(n2314) );
  CLKBUFX3 U174 ( .A(n2367), .Y(n2315) );
  CLKBUFX3 U175 ( .A(n2367), .Y(n2316) );
  CLKBUFX3 U176 ( .A(n2366), .Y(n2317) );
  CLKBUFX3 U177 ( .A(n2366), .Y(n2318) );
  CLKBUFX3 U178 ( .A(n2366), .Y(n2319) );
  CLKBUFX3 U179 ( .A(n2366), .Y(n2320) );
  CLKBUFX3 U180 ( .A(n2365), .Y(n2321) );
  CLKBUFX3 U181 ( .A(n2365), .Y(n2322) );
  CLKBUFX3 U182 ( .A(n2365), .Y(n2323) );
  CLKBUFX3 U183 ( .A(n2365), .Y(n2324) );
  CLKBUFX3 U184 ( .A(n2364), .Y(n2325) );
  CLKBUFX3 U185 ( .A(n2364), .Y(n2326) );
  CLKBUFX3 U186 ( .A(n2364), .Y(n2327) );
  CLKBUFX3 U187 ( .A(n2364), .Y(n2328) );
  CLKBUFX3 U188 ( .A(n2363), .Y(n2329) );
  CLKBUFX3 U189 ( .A(n2363), .Y(n2330) );
  CLKBUFX3 U190 ( .A(n2363), .Y(n2331) );
  CLKBUFX3 U191 ( .A(n2363), .Y(n2332) );
  CLKBUFX3 U192 ( .A(n2362), .Y(n2333) );
  CLKBUFX3 U193 ( .A(n2362), .Y(n2334) );
  CLKBUFX3 U194 ( .A(n2362), .Y(n2335) );
  CLKBUFX3 U195 ( .A(n2362), .Y(n2336) );
  CLKBUFX3 U196 ( .A(n2361), .Y(n2337) );
  CLKBUFX3 U197 ( .A(n2361), .Y(n2338) );
  CLKBUFX3 U198 ( .A(n2361), .Y(n2339) );
  CLKBUFX3 U199 ( .A(n2361), .Y(n2340) );
  CLKBUFX3 U200 ( .A(n2360), .Y(n2341) );
  CLKBUFX3 U201 ( .A(n2360), .Y(n2342) );
  CLKBUFX3 U202 ( .A(n2360), .Y(n2343) );
  CLKBUFX3 U203 ( .A(n2360), .Y(n2344) );
  CLKBUFX3 U204 ( .A(n2359), .Y(n2345) );
  CLKBUFX3 U205 ( .A(n2359), .Y(n2346) );
  CLKBUFX3 U206 ( .A(n2359), .Y(n2347) );
  CLKBUFX3 U207 ( .A(n2359), .Y(n2348) );
  CLKBUFX3 U208 ( .A(n2358), .Y(n2349) );
  CLKBUFX3 U209 ( .A(n2358), .Y(n2350) );
  CLKBUFX3 U210 ( .A(n2358), .Y(n2351) );
  CLKBUFX3 U211 ( .A(n2358), .Y(n2352) );
  CLKBUFX3 U212 ( .A(n2357), .Y(n2353) );
  CLKBUFX3 U213 ( .A(n2357), .Y(n2354) );
  CLKBUFX3 U214 ( .A(n2357), .Y(n2355) );
  CLKBUFX3 U215 ( .A(n2357), .Y(n2356) );
  CLKBUFX3 U216 ( .A(N18), .Y(n2079) );
  CLKBUFX3 U217 ( .A(n1544), .Y(n1552) );
  CLKBUFX3 U218 ( .A(n2085), .Y(n2102) );
  CLKBUFX3 U219 ( .A(n1559), .Y(n1577) );
  CLKBUFX3 U220 ( .A(n2084), .Y(n2101) );
  CLKBUFX3 U221 ( .A(n1559), .Y(n1576) );
  NOR2X1 U222 ( .A(n2083), .B(n2103), .Y(n1927) );
  NOR2X1 U223 ( .A(n2080), .B(n2103), .Y(n1922) );
  NOR2X1 U224 ( .A(n2082), .B(n2104), .Y(n1917) );
  NOR2X1 U225 ( .A(n2082), .B(n2104), .Y(n1912) );
  NOR2X1 U226 ( .A(n2083), .B(n2104), .Y(n1907) );
  NOR2X1 U227 ( .A(n2082), .B(n2104), .Y(n1902) );
  NOR2X1 U228 ( .A(n1558), .B(n1579), .Y(n1395) );
  NOR2X1 U229 ( .A(n1558), .B(n1580), .Y(n1390) );
  NOR2X1 U230 ( .A(n1558), .B(n1580), .Y(n1385) );
  NOR2X1 U231 ( .A(n1558), .B(n1580), .Y(n1380) );
  NOR2X1 U232 ( .A(n1558), .B(n1580), .Y(n1375) );
  CLKBUFX3 U233 ( .A(n2268), .Y(n2095) );
  CLKBUFX3 U234 ( .A(n2085), .Y(n2096) );
  CLKBUFX3 U235 ( .A(n2086), .Y(n2097) );
  CLKBUFX3 U236 ( .A(n2086), .Y(n2099) );
  CLKBUFX3 U237 ( .A(n2086), .Y(n2100) );
  CLKBUFX3 U238 ( .A(n2085), .Y(n2098) );
  CLKBUFX3 U239 ( .A(n2085), .Y(n2087) );
  CLKBUFX3 U240 ( .A(n2084), .Y(n2088) );
  CLKBUFX3 U241 ( .A(n2084), .Y(n2089) );
  CLKBUFX3 U242 ( .A(n2084), .Y(n2091) );
  CLKBUFX3 U243 ( .A(n2084), .Y(n2092) );
  CLKBUFX3 U244 ( .A(n2085), .Y(n2093) );
  CLKBUFX3 U245 ( .A(n2084), .Y(n2090) );
  CLKBUFX3 U246 ( .A(n2085), .Y(n2094) );
  CLKBUFX3 U247 ( .A(n1559), .Y(n1570) );
  CLKBUFX3 U248 ( .A(n1560), .Y(n1571) );
  CLKBUFX3 U249 ( .A(n1560), .Y(n1572) );
  CLKBUFX3 U250 ( .A(n1559), .Y(n1574) );
  CLKBUFX3 U251 ( .A(n1559), .Y(n1575) );
  CLKBUFX3 U252 ( .A(n1559), .Y(n1573) );
  CLKBUFX3 U253 ( .A(n1561), .Y(n1562) );
  CLKBUFX3 U254 ( .A(n1561), .Y(n1563) );
  CLKBUFX3 U255 ( .A(n1561), .Y(n1564) );
  CLKBUFX3 U256 ( .A(n1560), .Y(n1566) );
  CLKBUFX3 U257 ( .A(n1561), .Y(n1567) );
  CLKBUFX3 U258 ( .A(n1560), .Y(n1568) );
  CLKBUFX3 U259 ( .A(n1560), .Y(n1565) );
  CLKBUFX3 U260 ( .A(n1560), .Y(n1569) );
  BUFX4 U261 ( .A(n2083), .Y(n2076) );
  BUFX4 U262 ( .A(n2076), .Y(n2078) );
  BUFX4 U263 ( .A(n2081), .Y(n2077) );
  BUFX4 U264 ( .A(n2075), .Y(n2070) );
  BUFX4 U265 ( .A(n2082), .Y(n2071) );
  BUFX4 U266 ( .A(n2081), .Y(n2073) );
  BUFX4 U267 ( .A(n2083), .Y(n2075) );
  BUFX4 U268 ( .A(N18), .Y(n2072) );
  BUFX4 U269 ( .A(n2083), .Y(n2074) );
  BUFX4 U270 ( .A(n1545), .Y(n1551) );
  BUFX4 U271 ( .A(n1555), .Y(n1546) );
  BUFX4 U272 ( .A(n1545), .Y(n1548) );
  BUFX4 U273 ( .A(n1544), .Y(n1550) );
  BUFX4 U274 ( .A(n1545), .Y(n1547) );
  BUFX4 U275 ( .A(n1545), .Y(n1549) );
  CLKBUFX3 U276 ( .A(n1544), .Y(n1553) );
  CLKBUFX3 U277 ( .A(N18), .Y(n2080) );
  CLKBUFX3 U278 ( .A(n2075), .Y(n2081) );
  CLKBUFX3 U279 ( .A(n2076), .Y(n2082) );
  CLKBUFX3 U280 ( .A(N18), .Y(n2083) );
  CLKBUFX3 U281 ( .A(n1544), .Y(n1554) );
  CLKBUFX3 U282 ( .A(n1544), .Y(n1555) );
  CLKBUFX3 U283 ( .A(n1544), .Y(n1556) );
  CLKBUFX3 U284 ( .A(n1544), .Y(n1557) );
  CLKBUFX3 U285 ( .A(n2376), .Y(n2277) );
  CLKBUFX3 U286 ( .A(n2376), .Y(n2278) );
  CLKBUFX3 U287 ( .A(n2376), .Y(n2279) );
  CLKBUFX3 U288 ( .A(n2376), .Y(n2280) );
  CLKBUFX3 U289 ( .A(n2375), .Y(n2281) );
  CLKBUFX3 U290 ( .A(n2375), .Y(n2282) );
  CLKBUFX3 U291 ( .A(n2375), .Y(n2283) );
  CLKBUFX3 U292 ( .A(n2375), .Y(n2284) );
  CLKBUFX3 U293 ( .A(n2377), .Y(n2274) );
  CLKBUFX3 U294 ( .A(n2377), .Y(n2275) );
  CLKBUFX3 U295 ( .A(n2377), .Y(n2276) );
  CLKBUFX3 U296 ( .A(n2379), .Y(n2374) );
  CLKBUFX3 U297 ( .A(n2379), .Y(n2373) );
  CLKBUFX3 U298 ( .A(n2379), .Y(n2372) );
  CLKBUFX3 U299 ( .A(n2380), .Y(n2371) );
  CLKBUFX3 U300 ( .A(n2380), .Y(n2370) );
  CLKBUFX3 U301 ( .A(n2380), .Y(n2369) );
  CLKBUFX3 U302 ( .A(n2381), .Y(n2368) );
  CLKBUFX3 U303 ( .A(n2381), .Y(n2367) );
  CLKBUFX3 U304 ( .A(n2381), .Y(n2366) );
  CLKBUFX3 U305 ( .A(n2382), .Y(n2365) );
  CLKBUFX3 U306 ( .A(n2382), .Y(n2364) );
  CLKBUFX3 U307 ( .A(n2382), .Y(n2363) );
  CLKBUFX3 U308 ( .A(n2383), .Y(n2362) );
  CLKBUFX3 U309 ( .A(n2383), .Y(n2361) );
  CLKBUFX3 U310 ( .A(n2383), .Y(n2360) );
  CLKBUFX3 U311 ( .A(n2384), .Y(n2359) );
  CLKBUFX3 U312 ( .A(n2384), .Y(n2358) );
  CLKBUFX3 U313 ( .A(n2384), .Y(n2357) );
  CLKBUFX3 U314 ( .A(N20), .Y(n2062) );
  CLKBUFX3 U315 ( .A(n2269), .Y(n2063) );
  CLKBUFX3 U316 ( .A(n2269), .Y(n2064) );
  CLKBUFX3 U317 ( .A(N20), .Y(n2065) );
  CLKBUFX3 U318 ( .A(n1539), .Y(n1536) );
  CLKBUFX3 U319 ( .A(N15), .Y(n1537) );
  CLKBUFX3 U320 ( .A(n1537), .Y(n1538) );
  CLKBUFX3 U321 ( .A(N15), .Y(n1539) );
  CLKBUFX3 U322 ( .A(n1544), .Y(n1558) );
  CLKBUFX3 U323 ( .A(n2169), .Y(n2171) );
  CLKBUFX3 U324 ( .A(n8), .Y(n2170) );
  CLKBUFX3 U325 ( .A(n2069), .Y(n2066) );
  CLKBUFX3 U326 ( .A(n2068), .Y(n2067) );
  CLKBUFX3 U327 ( .A(N19), .Y(n2068) );
  CLKBUFX3 U328 ( .A(N19), .Y(n2069) );
  CLKBUFX3 U329 ( .A(n1543), .Y(n1540) );
  CLKBUFX3 U330 ( .A(N14), .Y(n1541) );
  CLKBUFX3 U331 ( .A(n1541), .Y(n1542) );
  CLKBUFX3 U332 ( .A(N14), .Y(n1543) );
  CLKBUFX3 U333 ( .A(N15), .Y(n1535) );
  CLKBUFX3 U334 ( .A(n1544), .Y(n1545) );
  CLKBUFX3 U335 ( .A(n2084), .Y(n2086) );
  CLKBUFX3 U336 ( .A(n1559), .Y(n1561) );
  CLKBUFX3 U337 ( .A(n2273), .Y(n2379) );
  CLKBUFX3 U338 ( .A(n2273), .Y(n2380) );
  CLKBUFX3 U339 ( .A(n2272), .Y(n2381) );
  CLKBUFX3 U340 ( .A(n2272), .Y(n2382) );
  CLKBUFX3 U341 ( .A(n2272), .Y(n2383) );
  CLKBUFX3 U342 ( .A(n2385), .Y(n2384) );
  CLKBUFX3 U343 ( .A(n2378), .Y(n2376) );
  CLKBUFX3 U344 ( .A(n2378), .Y(n2375) );
  CLKBUFX3 U345 ( .A(n2378), .Y(n2377) );
  CLKBUFX3 U346 ( .A(n11), .Y(n2261) );
  CLKBUFX3 U347 ( .A(n9), .Y(n2237) );
  CLKBUFX3 U348 ( .A(n10), .Y(n2213) );
  CLKBUFX3 U349 ( .A(n2187), .Y(n2189) );
  CLKBUFX3 U350 ( .A(n11), .Y(n2259) );
  CLKBUFX3 U351 ( .A(n11), .Y(n2260) );
  CLKBUFX3 U352 ( .A(n9), .Y(n2235) );
  CLKBUFX3 U353 ( .A(n9), .Y(n2236) );
  CLKBUFX3 U354 ( .A(n10), .Y(n2211) );
  CLKBUFX3 U355 ( .A(n10), .Y(n2212) );
  CLKBUFX3 U356 ( .A(n1), .Y(n2188) );
  CLKBUFX3 U357 ( .A(N21), .Y(n2061) );
  CLKBUFX3 U358 ( .A(N16), .Y(n1534) );
  CLKBUFX3 U359 ( .A(n26), .Y(n2258) );
  CLKBUFX3 U360 ( .A(n27), .Y(n2255) );
  CLKBUFX3 U361 ( .A(n28), .Y(n2252) );
  CLKBUFX3 U362 ( .A(n29), .Y(n2249) );
  CLKBUFX3 U363 ( .A(n30), .Y(n2246) );
  CLKBUFX3 U364 ( .A(n31), .Y(n2243) );
  CLKBUFX3 U365 ( .A(n12), .Y(n2240) );
  CLKBUFX3 U366 ( .A(n13), .Y(n2234) );
  CLKBUFX3 U367 ( .A(n14), .Y(n2231) );
  CLKBUFX3 U368 ( .A(n15), .Y(n2228) );
  CLKBUFX3 U369 ( .A(n16), .Y(n2225) );
  CLKBUFX3 U370 ( .A(n17), .Y(n2222) );
  CLKBUFX3 U371 ( .A(n18), .Y(n2219) );
  CLKBUFX3 U372 ( .A(n19), .Y(n2216) );
  CLKBUFX3 U373 ( .A(n20), .Y(n2210) );
  CLKBUFX3 U374 ( .A(n21), .Y(n2207) );
  CLKBUFX3 U375 ( .A(n22), .Y(n2204) );
  CLKBUFX3 U376 ( .A(n23), .Y(n2201) );
  CLKBUFX3 U377 ( .A(n24), .Y(n2198) );
  CLKBUFX3 U378 ( .A(n25), .Y(n2195) );
  CLKBUFX3 U379 ( .A(n2190), .Y(n2192) );
  CLKBUFX3 U380 ( .A(n2184), .Y(n2186) );
  CLKBUFX3 U381 ( .A(n2181), .Y(n2183) );
  CLKBUFX3 U382 ( .A(n2178), .Y(n2180) );
  CLKBUFX3 U383 ( .A(n2175), .Y(n2177) );
  CLKBUFX3 U384 ( .A(n2172), .Y(n2174) );
  CLKBUFX3 U385 ( .A(n26), .Y(n2256) );
  CLKBUFX3 U386 ( .A(n26), .Y(n2257) );
  CLKBUFX3 U387 ( .A(n27), .Y(n2253) );
  CLKBUFX3 U388 ( .A(n27), .Y(n2254) );
  CLKBUFX3 U389 ( .A(n28), .Y(n2250) );
  CLKBUFX3 U390 ( .A(n28), .Y(n2251) );
  CLKBUFX3 U391 ( .A(n29), .Y(n2247) );
  CLKBUFX3 U392 ( .A(n29), .Y(n2248) );
  CLKBUFX3 U393 ( .A(n30), .Y(n2244) );
  CLKBUFX3 U394 ( .A(n30), .Y(n2245) );
  CLKBUFX3 U395 ( .A(n31), .Y(n2241) );
  CLKBUFX3 U396 ( .A(n31), .Y(n2242) );
  CLKBUFX3 U397 ( .A(n12), .Y(n2238) );
  CLKBUFX3 U398 ( .A(n12), .Y(n2239) );
  CLKBUFX3 U399 ( .A(n13), .Y(n2232) );
  CLKBUFX3 U400 ( .A(n13), .Y(n2233) );
  CLKBUFX3 U401 ( .A(n14), .Y(n2229) );
  CLKBUFX3 U402 ( .A(n14), .Y(n2230) );
  CLKBUFX3 U403 ( .A(n15), .Y(n2226) );
  CLKBUFX3 U404 ( .A(n15), .Y(n2227) );
  CLKBUFX3 U405 ( .A(n16), .Y(n2223) );
  CLKBUFX3 U406 ( .A(n16), .Y(n2224) );
  CLKBUFX3 U407 ( .A(n17), .Y(n2220) );
  CLKBUFX3 U408 ( .A(n17), .Y(n2221) );
  CLKBUFX3 U409 ( .A(n18), .Y(n2217) );
  CLKBUFX3 U410 ( .A(n18), .Y(n2218) );
  CLKBUFX3 U411 ( .A(n19), .Y(n2214) );
  CLKBUFX3 U412 ( .A(n19), .Y(n2215) );
  CLKBUFX3 U413 ( .A(n20), .Y(n2208) );
  CLKBUFX3 U414 ( .A(n20), .Y(n2209) );
  CLKBUFX3 U415 ( .A(n21), .Y(n2205) );
  CLKBUFX3 U416 ( .A(n21), .Y(n2206) );
  CLKBUFX3 U417 ( .A(n22), .Y(n2202) );
  CLKBUFX3 U418 ( .A(n22), .Y(n2203) );
  CLKBUFX3 U419 ( .A(n23), .Y(n2199) );
  CLKBUFX3 U420 ( .A(n23), .Y(n2200) );
  CLKBUFX3 U421 ( .A(n24), .Y(n2196) );
  CLKBUFX3 U422 ( .A(n24), .Y(n2197) );
  CLKBUFX3 U423 ( .A(n25), .Y(n2193) );
  CLKBUFX3 U424 ( .A(n25), .Y(n2194) );
  CLKBUFX3 U425 ( .A(n2), .Y(n2191) );
  CLKBUFX3 U426 ( .A(n3), .Y(n2185) );
  CLKBUFX3 U427 ( .A(n4), .Y(n2182) );
  CLKBUFX3 U428 ( .A(n5), .Y(n2179) );
  CLKBUFX3 U429 ( .A(n6), .Y(n2176) );
  CLKBUFX3 U430 ( .A(n7), .Y(n2173) );
  CLKBUFX3 U431 ( .A(N17), .Y(n2084) );
  CLKBUFX3 U432 ( .A(N12), .Y(n1559) );
  CLKBUFX3 U433 ( .A(n2268), .Y(n2085) );
  CLKBUFX3 U434 ( .A(n1559), .Y(n1560) );
  CLKBUFX3 U435 ( .A(N13), .Y(n1544) );
  CLKBUFX3 U436 ( .A(n8), .Y(n2169) );
  CLKBUFX3 U437 ( .A(n2385), .Y(n2378) );
  CLKBUFX3 U438 ( .A(n2273), .Y(n2385) );
  CLKBUFX3 U439 ( .A(n1), .Y(n2187) );
  NOR4X1 U440 ( .A(n55), .B(N19), .C(n2270), .D(n2269), .Y(n52) );
  OR2X1 U441 ( .A(n2268), .B(N18), .Y(n55) );
  NOR4X1 U442 ( .A(n64), .B(N14), .C(n2271), .D(N15), .Y(n61) );
  OR2X1 U443 ( .A(N12), .B(N13), .Y(n64) );
  CLKBUFX3 U444 ( .A(n47), .Y(n2266) );
  CLKBUFX3 U445 ( .A(n47), .Y(n2267) );
  CLKBUFX3 U446 ( .A(n2449), .Y(n2167) );
  CLKBUFX3 U447 ( .A(n2448), .Y(n2166) );
  CLKBUFX3 U448 ( .A(n2445), .Y(n2160) );
  CLKBUFX3 U449 ( .A(n2444), .Y(n2157) );
  CLKBUFX3 U450 ( .A(n2443), .Y(n2156) );
  CLKBUFX3 U451 ( .A(n2437), .Y(n2144) );
  CLKBUFX3 U452 ( .A(n2430), .Y(n2130) );
  CLKBUFX3 U453 ( .A(n2427), .Y(n2124) );
  CLKBUFX3 U454 ( .A(n2426), .Y(n2122) );
  CLKBUFX3 U455 ( .A(n2425), .Y(n2120) );
  CLKBUFX3 U456 ( .A(n2422), .Y(n2114) );
  CLKBUFX3 U457 ( .A(n2448), .Y(n2165) );
  CLKBUFX3 U458 ( .A(n2445), .Y(n2159) );
  CLKBUFX3 U459 ( .A(n2443), .Y(n2155) );
  CLKBUFX3 U460 ( .A(n2437), .Y(n2143) );
  CLKBUFX3 U461 ( .A(n2430), .Y(n2129) );
  CLKBUFX3 U462 ( .A(n2427), .Y(n2123) );
  CLKBUFX3 U463 ( .A(n2426), .Y(n2121) );
  CLKBUFX3 U464 ( .A(n2425), .Y(n2119) );
  CLKBUFX3 U465 ( .A(n2422), .Y(n2113) );
  CLKBUFX3 U466 ( .A(n2447), .Y(n2164) );
  CLKBUFX3 U467 ( .A(n2446), .Y(n2162) );
  CLKBUFX3 U468 ( .A(n2434), .Y(n2138) );
  CLKBUFX3 U469 ( .A(n2420), .Y(n2110) );
  CLKBUFX3 U470 ( .A(n2418), .Y(n2106) );
  CLKBUFX3 U471 ( .A(n2447), .Y(n2163) );
  CLKBUFX3 U472 ( .A(n2446), .Y(n2161) );
  CLKBUFX3 U473 ( .A(n2434), .Y(n2137) );
  CLKBUFX3 U474 ( .A(n2420), .Y(n2109) );
  CLKBUFX3 U475 ( .A(n2418), .Y(n2105) );
  CLKBUFX3 U476 ( .A(n2442), .Y(n2153) );
  CLKBUFX3 U477 ( .A(n2441), .Y(n2151) );
  CLKBUFX3 U478 ( .A(n2440), .Y(n2149) );
  CLKBUFX3 U479 ( .A(n2439), .Y(n2147) );
  CLKBUFX3 U480 ( .A(n2438), .Y(n2146) );
  CLKBUFX3 U481 ( .A(n2436), .Y(n2142) );
  CLKBUFX3 U482 ( .A(n2435), .Y(n2140) );
  CLKBUFX3 U483 ( .A(n2433), .Y(n2136) );
  CLKBUFX3 U484 ( .A(n2432), .Y(n2134) );
  CLKBUFX3 U485 ( .A(n2431), .Y(n2132) );
  CLKBUFX3 U486 ( .A(n2429), .Y(n2128) );
  CLKBUFX3 U487 ( .A(n2428), .Y(n2126) );
  CLKBUFX3 U488 ( .A(n2424), .Y(n2118) );
  CLKBUFX3 U489 ( .A(n2423), .Y(n2116) );
  CLKBUFX3 U490 ( .A(n2421), .Y(n2112) );
  CLKBUFX3 U491 ( .A(n2419), .Y(n2108) );
  CLKBUFX3 U492 ( .A(n2438), .Y(n2145) );
  CLKBUFX3 U493 ( .A(n2436), .Y(n2141) );
  CLKBUFX3 U494 ( .A(n2435), .Y(n2139) );
  CLKBUFX3 U495 ( .A(n2433), .Y(n2135) );
  CLKBUFX3 U496 ( .A(n2432), .Y(n2133) );
  CLKBUFX3 U497 ( .A(n2431), .Y(n2131) );
  CLKBUFX3 U498 ( .A(n2429), .Y(n2127) );
  CLKBUFX3 U499 ( .A(n2428), .Y(n2125) );
  CLKBUFX3 U500 ( .A(n2424), .Y(n2117) );
  CLKBUFX3 U501 ( .A(n2423), .Y(n2115) );
  CLKBUFX3 U502 ( .A(n2421), .Y(n2111) );
  CLKBUFX3 U503 ( .A(n2419), .Y(n2107) );
  CLKBUFX3 U504 ( .A(n47), .Y(n2265) );
  CLKBUFX3 U505 ( .A(n2262), .Y(n2264) );
  CLKBUFX3 U506 ( .A(n2262), .Y(n2263) );
  CLKBUFX3 U507 ( .A(n2449), .Y(n2168) );
  CLKBUFX3 U508 ( .A(n2444), .Y(n2158) );
  CLKBUFX3 U509 ( .A(n2442), .Y(n2154) );
  CLKBUFX3 U510 ( .A(n2439), .Y(n2148) );
  CLKBUFX3 U511 ( .A(n2441), .Y(n2152) );
  CLKBUFX3 U512 ( .A(n2440), .Y(n2150) );
  CLKBUFX3 U513 ( .A(n3), .Y(n2184) );
  CLKBUFX3 U514 ( .A(n4), .Y(n2181) );
  CLKBUFX3 U515 ( .A(n5), .Y(n2178) );
  CLKBUFX3 U516 ( .A(n6), .Y(n2175) );
  CLKBUFX3 U517 ( .A(n7), .Y(n2172) );
  CLKBUFX3 U518 ( .A(n2), .Y(n2190) );
  NOR3X2 U519 ( .A(n2451), .B(n2450), .C(n2455), .Y(n100) );
  XNOR2X1 U520 ( .A(n2451), .B(n2269), .Y(n54) );
  XNOR2X1 U521 ( .A(n2451), .B(N15), .Y(n63) );
  XNOR2X1 U522 ( .A(n2450), .B(n2270), .Y(n53) );
  XNOR2X1 U523 ( .A(n2450), .B(n2271), .Y(n62) );
  CLKBUFX3 U524 ( .A(n56), .Y(n2262) );
  CLKBUFX3 U525 ( .A(N21), .Y(n2270) );
  CLKBUFX3 U526 ( .A(N16), .Y(n2271) );
  OAI2BB2XL U527 ( .B0(n2266), .B1(n2168), .A0N(N91), .A1N(n47), .Y(rdata2[0])
         );
  OAI2BB2XL U528 ( .B0(n2265), .B1(n2448), .A0N(N90), .A1N(n2266), .Y(
        rdata2[1]) );
  OAI2BB2XL U529 ( .B0(n2265), .B1(n2447), .A0N(N89), .A1N(n2267), .Y(
        rdata2[2]) );
  OAI2BB2XL U530 ( .B0(n2265), .B1(n2446), .A0N(N88), .A1N(n2267), .Y(
        rdata2[3]) );
  OAI2BB2XL U531 ( .B0(n2265), .B1(n2445), .A0N(N87), .A1N(n2267), .Y(
        rdata2[4]) );
  OAI2BB2XL U532 ( .B0(n2265), .B1(n2158), .A0N(N86), .A1N(n2267), .Y(
        rdata2[5]) );
  OAI2BB2XL U533 ( .B0(n2265), .B1(n2443), .A0N(N85), .A1N(n2267), .Y(
        rdata2[6]) );
  OAI2BB2XL U534 ( .B0(n2265), .B1(n2154), .A0N(N84), .A1N(n2266), .Y(
        rdata2[7]) );
  OAI2BB2XL U535 ( .B0(n2265), .B1(n2152), .A0N(N83), .A1N(n2266), .Y(
        rdata2[8]) );
  OAI2BB2XL U536 ( .B0(n2265), .B1(n2150), .A0N(N82), .A1N(n2266), .Y(
        rdata2[9]) );
  OAI2BB2XL U537 ( .B0(n2266), .B1(n2148), .A0N(N81), .A1N(n2265), .Y(
        rdata2[10]) );
  OAI2BB2XL U538 ( .B0(n2266), .B1(n2438), .A0N(N80), .A1N(n2267), .Y(
        rdata2[11]) );
  OAI2BB2XL U539 ( .B0(n2266), .B1(n2437), .A0N(N79), .A1N(n2267), .Y(
        rdata2[12]) );
  OAI2BB2XL U540 ( .B0(n2266), .B1(n2436), .A0N(N78), .A1N(n2267), .Y(
        rdata2[13]) );
  OAI2BB2XL U541 ( .B0(n2266), .B1(n2435), .A0N(N77), .A1N(n2267), .Y(
        rdata2[14]) );
  OAI2BB2XL U542 ( .B0(n2266), .B1(n2434), .A0N(N76), .A1N(n2267), .Y(
        rdata2[15]) );
  OAI2BB2XL U543 ( .B0(n2265), .B1(n2433), .A0N(N75), .A1N(n2267), .Y(
        rdata2[16]) );
  OAI2BB2XL U544 ( .B0(n2266), .B1(n2432), .A0N(N74), .A1N(n2266), .Y(
        rdata2[17]) );
  OAI2BB2XL U545 ( .B0(n2265), .B1(n2431), .A0N(N73), .A1N(n2267), .Y(
        rdata2[18]) );
  OAI2BB2XL U546 ( .B0(n2265), .B1(n2430), .A0N(N72), .A1N(n2266), .Y(
        rdata2[19]) );
  OAI2BB2XL U547 ( .B0(n2265), .B1(n2429), .A0N(N71), .A1N(n2266), .Y(
        rdata2[20]) );
  OAI2BB2XL U548 ( .B0(n2265), .B1(n2428), .A0N(N70), .A1N(n2266), .Y(
        rdata2[21]) );
  OAI2BB2XL U549 ( .B0(n2265), .B1(n2427), .A0N(N69), .A1N(n2266), .Y(
        rdata2[22]) );
  OAI2BB2XL U550 ( .B0(n2265), .B1(n2426), .A0N(N68), .A1N(n2267), .Y(
        rdata2[23]) );
  OAI2BB2XL U551 ( .B0(n2265), .B1(n2425), .A0N(N67), .A1N(n2266), .Y(
        rdata2[24]) );
  OAI2BB2XL U552 ( .B0(n2265), .B1(n2424), .A0N(N66), .A1N(n2267), .Y(
        rdata2[25]) );
  OAI2BB2XL U553 ( .B0(n2265), .B1(n2423), .A0N(N65), .A1N(n2267), .Y(
        rdata2[26]) );
  OAI2BB2XL U554 ( .B0(n2267), .B1(n2422), .A0N(N64), .A1N(n2267), .Y(
        rdata2[27]) );
  OAI2BB2XL U555 ( .B0(n2266), .B1(n2421), .A0N(N63), .A1N(n2267), .Y(
        rdata2[28]) );
  OAI2BB2XL U556 ( .B0(n2265), .B1(n2420), .A0N(N62), .A1N(n2267), .Y(
        rdata2[29]) );
  OAI2BB2XL U557 ( .B0(n2267), .B1(n2419), .A0N(N61), .A1N(n2267), .Y(
        rdata2[30]) );
  OAI2BB2XL U558 ( .B0(n2266), .B1(n2418), .A0N(N60), .A1N(n2267), .Y(
        rdata2[31]) );
  OAI2BB2XL U559 ( .B0(n2168), .B1(n2263), .A0N(N56), .A1N(n2263), .Y(
        rdata1[0]) );
  OAI2BB2XL U560 ( .B0(n2166), .B1(n2264), .A0N(N55), .A1N(n2262), .Y(
        rdata1[1]) );
  OAI2BB2XL U561 ( .B0(n2164), .B1(n2263), .A0N(N54), .A1N(n56), .Y(rdata1[2])
         );
  OAI2BB2XL U562 ( .B0(n2162), .B1(n2263), .A0N(N53), .A1N(n2262), .Y(
        rdata1[3]) );
  OAI2BB2XL U563 ( .B0(n2160), .B1(n2263), .A0N(N52), .A1N(n2262), .Y(
        rdata1[4]) );
  OAI2BB2XL U564 ( .B0(n2158), .B1(n2263), .A0N(N51), .A1N(n2262), .Y(
        rdata1[5]) );
  OAI2BB2XL U565 ( .B0(n2156), .B1(n2263), .A0N(N50), .A1N(n2262), .Y(
        rdata1[6]) );
  OAI2BB2XL U566 ( .B0(n2154), .B1(n2263), .A0N(N49), .A1N(n2262), .Y(
        rdata1[7]) );
  OAI2BB2XL U567 ( .B0(n2152), .B1(n2263), .A0N(N48), .A1N(n2262), .Y(
        rdata1[8]) );
  OAI2BB2XL U568 ( .B0(n2150), .B1(n2264), .A0N(N47), .A1N(n2262), .Y(
        rdata1[9]) );
  OAI2BB2XL U569 ( .B0(n2148), .B1(n2262), .A0N(N46), .A1N(n2264), .Y(
        rdata1[10]) );
  OAI2BB2XL U570 ( .B0(n2146), .B1(n2262), .A0N(N45), .A1N(n2263), .Y(
        rdata1[11]) );
  OAI2BB2XL U571 ( .B0(n2144), .B1(n2262), .A0N(N44), .A1N(n2264), .Y(
        rdata1[12]) );
  OAI2BB2XL U572 ( .B0(n2142), .B1(n2262), .A0N(N43), .A1N(n2263), .Y(
        rdata1[13]) );
  OAI2BB2XL U573 ( .B0(n2140), .B1(n2262), .A0N(N42), .A1N(n2264), .Y(
        rdata1[14]) );
  OAI2BB2XL U574 ( .B0(n2138), .B1(n2262), .A0N(N41), .A1N(n2263), .Y(
        rdata1[15]) );
  OAI2BB2XL U575 ( .B0(n2136), .B1(n2264), .A0N(N40), .A1N(n2262), .Y(
        rdata1[16]) );
  OAI2BB2XL U576 ( .B0(n2134), .B1(n2262), .A0N(N39), .A1N(n2264), .Y(
        rdata1[17]) );
  OAI2BB2XL U577 ( .B0(n2132), .B1(n2264), .A0N(N38), .A1N(n2262), .Y(
        rdata1[18]) );
  OAI2BB2XL U578 ( .B0(n2130), .B1(n2264), .A0N(N37), .A1N(n2264), .Y(
        rdata1[19]) );
  OAI2BB2XL U579 ( .B0(n2128), .B1(n2264), .A0N(N36), .A1N(n2264), .Y(
        rdata1[20]) );
  OAI2BB2XL U580 ( .B0(n2126), .B1(n2264), .A0N(N35), .A1N(n2263), .Y(
        rdata1[21]) );
  OAI2BB2XL U581 ( .B0(n2124), .B1(n2264), .A0N(N34), .A1N(n2263), .Y(
        rdata1[22]) );
  OAI2BB2XL U582 ( .B0(n2122), .B1(n2264), .A0N(N33), .A1N(n2262), .Y(
        rdata1[23]) );
  OAI2BB2XL U583 ( .B0(n2120), .B1(n2264), .A0N(N32), .A1N(n2264), .Y(
        rdata1[24]) );
  OAI2BB2XL U584 ( .B0(n2424), .B1(n2264), .A0N(N31), .A1N(n2264), .Y(
        rdata1[25]) );
  OAI2BB2XL U585 ( .B0(n2116), .B1(n2264), .A0N(N30), .A1N(n2262), .Y(
        rdata1[26]) );
  OAI2BB2XL U586 ( .B0(n2114), .B1(n2263), .A0N(N29), .A1N(n56), .Y(rdata1[27]) );
  OAI2BB2XL U587 ( .B0(n2112), .B1(n2263), .A0N(N28), .A1N(n56), .Y(rdata1[28]) );
  OAI2BB2XL U588 ( .B0(n2110), .B1(n2263), .A0N(N27), .A1N(n56), .Y(rdata1[29]) );
  OAI2BB2XL U589 ( .B0(n2108), .B1(n2263), .A0N(N26), .A1N(n56), .Y(rdata1[30]) );
  OAI2BB2XL U590 ( .B0(n2106), .B1(n2263), .A0N(N25), .A1N(n56), .Y(rdata1[31]) );
  OAI2BB2XL U591 ( .B0(n2121), .B1(n2259), .A0N(\register[1][23] ), .A1N(n2261), .Y(n131) );
  OAI2BB2XL U592 ( .B0(n2424), .B1(n11), .A0N(\register[1][25] ), .A1N(n2261), 
        .Y(n133) );
  OAI2BB2XL U593 ( .B0(n2115), .B1(n2260), .A0N(\register[1][26] ), .A1N(n2261), .Y(n134) );
  OAI2BB2XL U594 ( .B0(n2113), .B1(n2259), .A0N(\register[1][27] ), .A1N(n2261), .Y(n135) );
  OAI2BB2XL U595 ( .B0(n2111), .B1(n2260), .A0N(\register[1][28] ), .A1N(n2261), .Y(n136) );
  OAI2BB2XL U596 ( .B0(n2109), .B1(n11), .A0N(\register[1][29] ), .A1N(n2261), 
        .Y(n137) );
  OAI2BB2XL U597 ( .B0(n2107), .B1(n11), .A0N(\register[1][30] ), .A1N(n2259), 
        .Y(n138) );
  OAI2BB2XL U598 ( .B0(n2105), .B1(n11), .A0N(\register[1][31] ), .A1N(n2260), 
        .Y(n139) );
  OAI2BB2XL U599 ( .B0(n2122), .B1(n2236), .A0N(\register[9][23] ), .A1N(n2235), .Y(n387) );
  OAI2BB2XL U600 ( .B0(n2118), .B1(n2235), .A0N(\register[9][25] ), .A1N(n2237), .Y(n389) );
  OAI2BB2XL U601 ( .B0(n2116), .B1(n2236), .A0N(\register[9][26] ), .A1N(n2237), .Y(n390) );
  OAI2BB2XL U602 ( .B0(n2114), .B1(n2235), .A0N(\register[9][27] ), .A1N(n2237), .Y(n391) );
  OAI2BB2XL U603 ( .B0(n2112), .B1(n9), .A0N(\register[9][28] ), .A1N(n2237), 
        .Y(n392) );
  OAI2BB2XL U604 ( .B0(n2110), .B1(n9), .A0N(\register[9][29] ), .A1N(n2237), 
        .Y(n393) );
  OAI2BB2XL U605 ( .B0(n2108), .B1(n9), .A0N(\register[9][30] ), .A1N(n2235), 
        .Y(n394) );
  OAI2BB2XL U606 ( .B0(n2106), .B1(n9), .A0N(\register[9][31] ), .A1N(n2236), 
        .Y(n395) );
  OAI2BB2XL U607 ( .B0(n2122), .B1(n2212), .A0N(\register[17][23] ), .A1N(
        n2211), .Y(n643) );
  OAI2BB2XL U608 ( .B0(n2118), .B1(n2211), .A0N(\register[17][25] ), .A1N(
        n2213), .Y(n645) );
  OAI2BB2XL U609 ( .B0(n2116), .B1(n2212), .A0N(\register[17][26] ), .A1N(
        n2213), .Y(n646) );
  OAI2BB2XL U610 ( .B0(n2114), .B1(n2211), .A0N(\register[17][27] ), .A1N(
        n2213), .Y(n647) );
  OAI2BB2XL U611 ( .B0(n2112), .B1(n10), .A0N(\register[17][28] ), .A1N(n2213), 
        .Y(n648) );
  OAI2BB2XL U612 ( .B0(n2110), .B1(n10), .A0N(\register[17][29] ), .A1N(n2213), 
        .Y(n649) );
  OAI2BB2XL U613 ( .B0(n2108), .B1(n10), .A0N(\register[17][30] ), .A1N(n2211), 
        .Y(n650) );
  OAI2BB2XL U614 ( .B0(n2106), .B1(n10), .A0N(\register[17][31] ), .A1N(n2212), 
        .Y(n651) );
  OAI2BB2XL U615 ( .B0(n2121), .B1(n2187), .A0N(\register[25][23] ), .A1N(
        n2187), .Y(n899) );
  OAI2BB2XL U616 ( .B0(n2117), .B1(n2187), .A0N(\register[25][25] ), .A1N(
        n2189), .Y(n901) );
  OAI2BB2XL U617 ( .B0(n2115), .B1(n2187), .A0N(\register[25][26] ), .A1N(
        n2189), .Y(n902) );
  OAI2BB2XL U618 ( .B0(n2113), .B1(n2187), .A0N(\register[25][27] ), .A1N(
        n2189), .Y(n903) );
  OAI2BB2XL U619 ( .B0(n2111), .B1(n2187), .A0N(\register[25][28] ), .A1N(
        n2189), .Y(n904) );
  OAI2BB2XL U620 ( .B0(n2109), .B1(n2187), .A0N(\register[25][29] ), .A1N(
        n2189), .Y(n905) );
  OAI2BB2XL U621 ( .B0(n2107), .B1(n2187), .A0N(\register[25][30] ), .A1N(
        n2188), .Y(n906) );
  OAI2BB2XL U622 ( .B0(n2105), .B1(n2187), .A0N(\register[25][31] ), .A1N(
        n2188), .Y(n907) );
  OAI2BB2XL U623 ( .B0(n2167), .B1(n2236), .A0N(\register[9][0] ), .A1N(n2236), 
        .Y(n364) );
  OAI2BB2XL U624 ( .B0(n2166), .B1(n2235), .A0N(\register[9][1] ), .A1N(n2235), 
        .Y(n365) );
  OAI2BB2XL U625 ( .B0(n2164), .B1(n2235), .A0N(\register[9][2] ), .A1N(n2236), 
        .Y(n366) );
  OAI2BB2XL U626 ( .B0(n2162), .B1(n2235), .A0N(\register[9][3] ), .A1N(n2237), 
        .Y(n367) );
  OAI2BB2XL U627 ( .B0(n2160), .B1(n2235), .A0N(\register[9][4] ), .A1N(n2235), 
        .Y(n368) );
  OAI2BB2XL U628 ( .B0(n2157), .B1(n2235), .A0N(\register[9][5] ), .A1N(n2237), 
        .Y(n369) );
  OAI2BB2XL U629 ( .B0(n2156), .B1(n2235), .A0N(\register[9][6] ), .A1N(n2237), 
        .Y(n370) );
  OAI2BB2XL U630 ( .B0(n2153), .B1(n2235), .A0N(\register[9][7] ), .A1N(n2237), 
        .Y(n371) );
  OAI2BB2XL U631 ( .B0(n2151), .B1(n2235), .A0N(\register[9][8] ), .A1N(n2237), 
        .Y(n372) );
  OAI2BB2XL U632 ( .B0(n2149), .B1(n2235), .A0N(\register[9][9] ), .A1N(n2237), 
        .Y(n373) );
  OAI2BB2XL U633 ( .B0(n2147), .B1(n2235), .A0N(\register[9][10] ), .A1N(n2237), .Y(n374) );
  OAI2BB2XL U634 ( .B0(n2146), .B1(n2235), .A0N(\register[9][11] ), .A1N(n2237), .Y(n375) );
  OAI2BB2XL U635 ( .B0(n2144), .B1(n2235), .A0N(\register[9][12] ), .A1N(n2237), .Y(n376) );
  OAI2BB2XL U636 ( .B0(n2142), .B1(n2236), .A0N(\register[9][13] ), .A1N(n2237), .Y(n377) );
  OAI2BB2XL U637 ( .B0(n2140), .B1(n2236), .A0N(\register[9][14] ), .A1N(n2237), .Y(n378) );
  OAI2BB2XL U638 ( .B0(n2138), .B1(n2236), .A0N(\register[9][15] ), .A1N(n2237), .Y(n379) );
  OAI2BB2XL U639 ( .B0(n2136), .B1(n2236), .A0N(\register[9][16] ), .A1N(n2237), .Y(n380) );
  OAI2BB2XL U640 ( .B0(n2134), .B1(n2236), .A0N(\register[9][17] ), .A1N(n2237), .Y(n381) );
  OAI2BB2XL U641 ( .B0(n2132), .B1(n2236), .A0N(\register[9][18] ), .A1N(n2236), .Y(n382) );
  OAI2BB2XL U642 ( .B0(n2130), .B1(n2236), .A0N(\register[9][19] ), .A1N(n2235), .Y(n383) );
  OAI2BB2XL U643 ( .B0(n2128), .B1(n2236), .A0N(\register[9][20] ), .A1N(n2237), .Y(n384) );
  OAI2BB2XL U644 ( .B0(n2126), .B1(n2236), .A0N(\register[9][21] ), .A1N(n2236), .Y(n385) );
  OAI2BB2XL U645 ( .B0(n2124), .B1(n2236), .A0N(\register[9][22] ), .A1N(n2237), .Y(n386) );
  OAI2BB2XL U646 ( .B0(n2120), .B1(n2236), .A0N(\register[9][24] ), .A1N(n2237), .Y(n388) );
  OAI2BB2XL U647 ( .B0(n2167), .B1(n2212), .A0N(\register[17][0] ), .A1N(n2212), .Y(n620) );
  OAI2BB2XL U648 ( .B0(n2166), .B1(n2211), .A0N(\register[17][1] ), .A1N(n2211), .Y(n621) );
  OAI2BB2XL U649 ( .B0(n2164), .B1(n2211), .A0N(\register[17][2] ), .A1N(n2212), .Y(n622) );
  OAI2BB2XL U650 ( .B0(n2162), .B1(n2211), .A0N(\register[17][3] ), .A1N(n2213), .Y(n623) );
  OAI2BB2XL U651 ( .B0(n2160), .B1(n2211), .A0N(\register[17][4] ), .A1N(n2211), .Y(n624) );
  OAI2BB2XL U652 ( .B0(n2157), .B1(n2211), .A0N(\register[17][5] ), .A1N(n2213), .Y(n625) );
  OAI2BB2XL U653 ( .B0(n2156), .B1(n2211), .A0N(\register[17][6] ), .A1N(n2213), .Y(n626) );
  OAI2BB2XL U654 ( .B0(n2153), .B1(n2211), .A0N(\register[17][7] ), .A1N(n2213), .Y(n627) );
  OAI2BB2XL U655 ( .B0(n2151), .B1(n2211), .A0N(\register[17][8] ), .A1N(n2213), .Y(n628) );
  OAI2BB2XL U656 ( .B0(n2149), .B1(n2211), .A0N(\register[17][9] ), .A1N(n2213), .Y(n629) );
  OAI2BB2XL U657 ( .B0(n2147), .B1(n2211), .A0N(\register[17][10] ), .A1N(
        n2213), .Y(n630) );
  OAI2BB2XL U658 ( .B0(n2146), .B1(n2211), .A0N(\register[17][11] ), .A1N(
        n2213), .Y(n631) );
  OAI2BB2XL U659 ( .B0(n2144), .B1(n2211), .A0N(\register[17][12] ), .A1N(
        n2213), .Y(n632) );
  OAI2BB2XL U660 ( .B0(n2142), .B1(n2212), .A0N(\register[17][13] ), .A1N(
        n2213), .Y(n633) );
  OAI2BB2XL U661 ( .B0(n2140), .B1(n2212), .A0N(\register[17][14] ), .A1N(
        n2213), .Y(n634) );
  OAI2BB2XL U662 ( .B0(n2138), .B1(n2212), .A0N(\register[17][15] ), .A1N(
        n2213), .Y(n635) );
  OAI2BB2XL U663 ( .B0(n2136), .B1(n2212), .A0N(\register[17][16] ), .A1N(
        n2213), .Y(n636) );
  OAI2BB2XL U664 ( .B0(n2134), .B1(n2212), .A0N(\register[17][17] ), .A1N(
        n2213), .Y(n637) );
  OAI2BB2XL U665 ( .B0(n2132), .B1(n2212), .A0N(\register[17][18] ), .A1N(
        n2212), .Y(n638) );
  OAI2BB2XL U666 ( .B0(n2130), .B1(n2212), .A0N(\register[17][19] ), .A1N(
        n2211), .Y(n639) );
  OAI2BB2XL U667 ( .B0(n2128), .B1(n2212), .A0N(\register[17][20] ), .A1N(
        n2213), .Y(n640) );
  OAI2BB2XL U668 ( .B0(n2126), .B1(n2212), .A0N(\register[17][21] ), .A1N(
        n2212), .Y(n641) );
  OAI2BB2XL U669 ( .B0(n2124), .B1(n2212), .A0N(\register[17][22] ), .A1N(
        n2213), .Y(n642) );
  OAI2BB2XL U670 ( .B0(n2120), .B1(n2212), .A0N(\register[17][24] ), .A1N(
        n2213), .Y(n644) );
  OAI2BB2XL U671 ( .B0(n2167), .B1(n2188), .A0N(\register[25][0] ), .A1N(n2188), .Y(n876) );
  OAI2BB2XL U672 ( .B0(n2165), .B1(n1), .A0N(\register[25][1] ), .A1N(n2188), 
        .Y(n877) );
  OAI2BB2XL U673 ( .B0(n2163), .B1(n1), .A0N(\register[25][2] ), .A1N(n2188), 
        .Y(n878) );
  OAI2BB2XL U674 ( .B0(n2161), .B1(n1), .A0N(\register[25][3] ), .A1N(n2189), 
        .Y(n879) );
  OAI2BB2XL U675 ( .B0(n2159), .B1(n1), .A0N(\register[25][4] ), .A1N(n2188), 
        .Y(n880) );
  OAI2BB2XL U676 ( .B0(n2157), .B1(n2188), .A0N(\register[25][5] ), .A1N(n2189), .Y(n881) );
  OAI2BB2XL U677 ( .B0(n2155), .B1(n1), .A0N(\register[25][6] ), .A1N(n2189), 
        .Y(n882) );
  OAI2BB2XL U678 ( .B0(n2153), .B1(n2188), .A0N(\register[25][7] ), .A1N(n2189), .Y(n883) );
  OAI2BB2XL U679 ( .B0(n2151), .B1(n2188), .A0N(\register[25][8] ), .A1N(n2189), .Y(n884) );
  OAI2BB2XL U680 ( .B0(n2149), .B1(n2187), .A0N(\register[25][9] ), .A1N(n2189), .Y(n885) );
  OAI2BB2XL U681 ( .B0(n2147), .B1(n2187), .A0N(\register[25][10] ), .A1N(
        n2189), .Y(n886) );
  OAI2BB2XL U682 ( .B0(n2145), .B1(n2187), .A0N(\register[25][11] ), .A1N(
        n2189), .Y(n887) );
  OAI2BB2XL U683 ( .B0(n2143), .B1(n2187), .A0N(\register[25][12] ), .A1N(
        n2189), .Y(n888) );
  OAI2BB2XL U684 ( .B0(n2141), .B1(n2188), .A0N(\register[25][13] ), .A1N(
        n2189), .Y(n889) );
  OAI2BB2XL U685 ( .B0(n2139), .B1(n2188), .A0N(\register[25][14] ), .A1N(
        n2189), .Y(n890) );
  OAI2BB2XL U686 ( .B0(n2137), .B1(n2188), .A0N(\register[25][15] ), .A1N(
        n2187), .Y(n891) );
  OAI2BB2XL U687 ( .B0(n2135), .B1(n2188), .A0N(\register[25][16] ), .A1N(
        n2189), .Y(n892) );
  OAI2BB2XL U688 ( .B0(n2133), .B1(n2188), .A0N(\register[25][17] ), .A1N(
        n2187), .Y(n893) );
  OAI2BB2XL U689 ( .B0(n2131), .B1(n2188), .A0N(\register[25][18] ), .A1N(
        n2187), .Y(n894) );
  OAI2BB2XL U690 ( .B0(n2129), .B1(n2188), .A0N(\register[25][19] ), .A1N(
        n2187), .Y(n895) );
  OAI2BB2XL U691 ( .B0(n2127), .B1(n2188), .A0N(\register[25][20] ), .A1N(
        n2187), .Y(n896) );
  OAI2BB2XL U692 ( .B0(n2125), .B1(n2188), .A0N(\register[25][21] ), .A1N(
        n2187), .Y(n897) );
  OAI2BB2XL U693 ( .B0(n2123), .B1(n2188), .A0N(\register[25][22] ), .A1N(
        n2189), .Y(n898) );
  OAI2BB2XL U694 ( .B0(n2119), .B1(n2188), .A0N(\register[25][24] ), .A1N(
        n2189), .Y(n900) );
  OAI2BB2XL U695 ( .B0(n2168), .B1(n2260), .A0N(\register[1][0] ), .A1N(n2260), 
        .Y(n108) );
  OAI2BB2XL U696 ( .B0(n2165), .B1(n2259), .A0N(\register[1][1] ), .A1N(n2259), 
        .Y(n109) );
  OAI2BB2XL U697 ( .B0(n2163), .B1(n2259), .A0N(\register[1][2] ), .A1N(n2260), 
        .Y(n110) );
  OAI2BB2XL U698 ( .B0(n2161), .B1(n2259), .A0N(\register[1][3] ), .A1N(n2261), 
        .Y(n111) );
  OAI2BB2XL U699 ( .B0(n2159), .B1(n2259), .A0N(\register[1][4] ), .A1N(n2259), 
        .Y(n112) );
  OAI2BB2XL U700 ( .B0(n2158), .B1(n2259), .A0N(\register[1][5] ), .A1N(n2261), 
        .Y(n113) );
  OAI2BB2XL U701 ( .B0(n2155), .B1(n2259), .A0N(\register[1][6] ), .A1N(n2261), 
        .Y(n114) );
  OAI2BB2XL U702 ( .B0(n2154), .B1(n2259), .A0N(\register[1][7] ), .A1N(n2261), 
        .Y(n115) );
  OAI2BB2XL U703 ( .B0(n2152), .B1(n2259), .A0N(\register[1][8] ), .A1N(n2261), 
        .Y(n116) );
  OAI2BB2XL U704 ( .B0(n2150), .B1(n2259), .A0N(\register[1][9] ), .A1N(n2261), 
        .Y(n117) );
  OAI2BB2XL U705 ( .B0(n2148), .B1(n2259), .A0N(\register[1][10] ), .A1N(n2261), .Y(n118) );
  OAI2BB2XL U706 ( .B0(n2145), .B1(n2259), .A0N(\register[1][11] ), .A1N(n2261), .Y(n119) );
  OAI2BB2XL U707 ( .B0(n2143), .B1(n2259), .A0N(\register[1][12] ), .A1N(n2261), .Y(n120) );
  OAI2BB2XL U708 ( .B0(n2141), .B1(n2260), .A0N(\register[1][13] ), .A1N(n2261), .Y(n121) );
  OAI2BB2XL U709 ( .B0(n2139), .B1(n2260), .A0N(\register[1][14] ), .A1N(n2261), .Y(n122) );
  OAI2BB2XL U710 ( .B0(n2137), .B1(n2260), .A0N(\register[1][15] ), .A1N(n2261), .Y(n123) );
  OAI2BB2XL U711 ( .B0(n2135), .B1(n2260), .A0N(\register[1][16] ), .A1N(n2261), .Y(n124) );
  OAI2BB2XL U712 ( .B0(n2133), .B1(n2260), .A0N(\register[1][17] ), .A1N(n2259), .Y(n125) );
  OAI2BB2XL U713 ( .B0(n2131), .B1(n2260), .A0N(\register[1][18] ), .A1N(n2260), .Y(n126) );
  OAI2BB2XL U714 ( .B0(n2129), .B1(n2260), .A0N(\register[1][19] ), .A1N(n2261), .Y(n127) );
  OAI2BB2XL U715 ( .B0(n2127), .B1(n2260), .A0N(\register[1][20] ), .A1N(n2259), .Y(n128) );
  OAI2BB2XL U716 ( .B0(n2125), .B1(n2260), .A0N(\register[1][21] ), .A1N(n2260), .Y(n129) );
  OAI2BB2XL U717 ( .B0(n2123), .B1(n2260), .A0N(\register[1][22] ), .A1N(n2261), .Y(n130) );
  OAI2BB2XL U718 ( .B0(n2119), .B1(n2260), .A0N(\register[1][24] ), .A1N(n2261), .Y(n132) );
  NAND4X1 U719 ( .A(n48), .B(n49), .C(n50), .D(n51), .Y(n47) );
  NOR4X1 U720 ( .A(n52), .B(n2455), .C(n53), .D(n54), .Y(n51) );
  NAND4X1 U721 ( .A(n57), .B(n58), .C(n59), .D(n60), .Y(n56) );
  NOR4X1 U722 ( .A(n61), .B(n2455), .C(n62), .D(n63), .Y(n60) );
  MXI2X1 U723 ( .A(n1581), .B(n1582), .S0(N21), .Y(N91) );
  MX4X1 U724 ( .A(n1648), .B(n1646), .C(n1647), .D(n1645), .S0(n2064), .S1(
        n2067), .Y(n1582) );
  MX4X1 U725 ( .A(n1652), .B(n1650), .C(n1651), .D(n1649), .S0(n2063), .S1(
        n2069), .Y(n1581) );
  MXI4X1 U726 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n2094), .S1(n2075), .Y(
        n1648) );
  MXI2X1 U727 ( .A(n1583), .B(n1584), .S0(n2061), .Y(N90) );
  MX4X1 U728 ( .A(n1660), .B(n1658), .C(n1659), .D(n1657), .S0(N20), .S1(n2066), .Y(n1583) );
  MX4X1 U729 ( .A(n1656), .B(n1654), .C(n1655), .D(n1653), .S0(n2062), .S1(
        n2069), .Y(n1584) );
  MXI4X1 U730 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n2095), .S1(n2075), .Y(
        n1658) );
  MXI2X1 U731 ( .A(n1585), .B(n1586), .S0(n2061), .Y(N89) );
  MX4X1 U732 ( .A(n1668), .B(n1666), .C(n1667), .D(n1665), .S0(n2062), .S1(
        n2066), .Y(n1585) );
  MX4X1 U733 ( .A(n1664), .B(n1662), .C(n1663), .D(n1661), .S0(n2062), .S1(
        n2066), .Y(n1586) );
  MXI4X1 U734 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n2095), .S1(n2075), .Y(
        n1666) );
  MXI2X1 U735 ( .A(n1587), .B(n1588), .S0(n2061), .Y(N88) );
  MX4X1 U736 ( .A(n1676), .B(n1674), .C(n1675), .D(n1673), .S0(n2062), .S1(
        n2066), .Y(n1587) );
  MX4X1 U737 ( .A(n1672), .B(n1670), .C(n1671), .D(n1669), .S0(n2062), .S1(
        n2066), .Y(n1588) );
  MXI4X1 U738 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n2096), .S1(n2076), .Y(
        n1674) );
  MXI2X1 U739 ( .A(n1589), .B(n1590), .S0(N21), .Y(N87) );
  MX4X1 U740 ( .A(n1684), .B(n1682), .C(n1683), .D(n1681), .S0(n2062), .S1(
        n2066), .Y(n1589) );
  MX4X1 U741 ( .A(n1680), .B(n1678), .C(n1679), .D(n1677), .S0(n2062), .S1(
        n2066), .Y(n1590) );
  MXI4X1 U742 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n2096), .S1(n2076), .Y(
        n1682) );
  MXI2X1 U743 ( .A(n1591), .B(n1592), .S0(n2061), .Y(N86) );
  MX4X1 U744 ( .A(n1692), .B(n1690), .C(n1691), .D(n1689), .S0(n2062), .S1(
        n2066), .Y(n1591) );
  MX4X1 U745 ( .A(n1688), .B(n1686), .C(n1687), .D(n1685), .S0(n2062), .S1(
        n2066), .Y(n1592) );
  MXI4X1 U746 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n2097), .S1(n2076), .Y(
        n1690) );
  MXI2X1 U747 ( .A(n1593), .B(n1594), .S0(n2061), .Y(N85) );
  MX4X1 U748 ( .A(n1700), .B(n1698), .C(n1699), .D(n1697), .S0(n2062), .S1(
        n2066), .Y(n1593) );
  MX4X1 U749 ( .A(n1696), .B(n1694), .C(n1695), .D(n1693), .S0(n2062), .S1(
        n2066), .Y(n1594) );
  MXI4X1 U750 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n2097), .S1(n2077), .Y(
        n1698) );
  MXI2X1 U751 ( .A(n1595), .B(n1596), .S0(n2270), .Y(N84) );
  MX4X1 U752 ( .A(n1708), .B(n1706), .C(n1707), .D(n1705), .S0(n2062), .S1(
        n2066), .Y(n1595) );
  MX4X1 U753 ( .A(n1704), .B(n1702), .C(n1703), .D(n1701), .S0(n2062), .S1(
        n2066), .Y(n1596) );
  MXI4X1 U754 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n2098), .S1(n2077), .Y(
        n1706) );
  MXI2X1 U755 ( .A(n1597), .B(n1598), .S0(n2061), .Y(N83) );
  MX4X1 U756 ( .A(n1716), .B(n1714), .C(n1715), .D(n1713), .S0(n2063), .S1(
        n2067), .Y(n1597) );
  MX4X1 U757 ( .A(n1712), .B(n1710), .C(n1711), .D(n1709), .S0(n2063), .S1(
        n2067), .Y(n1598) );
  MXI4X1 U758 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n2098), .S1(n2077), .Y(
        n1714) );
  MXI2X1 U759 ( .A(n1599), .B(n1600), .S0(n2061), .Y(N82) );
  MX4X1 U760 ( .A(n1724), .B(n1722), .C(n1723), .D(n1721), .S0(n2063), .S1(
        n2067), .Y(n1599) );
  MX4X1 U761 ( .A(n1720), .B(n1718), .C(n1719), .D(n1717), .S0(n2063), .S1(
        n2067), .Y(n1600) );
  MXI4X1 U762 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n2099), .S1(n2082), .Y(
        n1722) );
  MXI2X1 U763 ( .A(n1601), .B(n1602), .S0(n2061), .Y(N81) );
  MX4X1 U764 ( .A(n1732), .B(n1730), .C(n1731), .D(n1729), .S0(n2063), .S1(
        n2067), .Y(n1601) );
  MX4X1 U765 ( .A(n1728), .B(n1726), .C(n1727), .D(n1725), .S0(n2063), .S1(
        n2067), .Y(n1602) );
  MXI4X1 U766 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n2099), .S1(n2076), 
        .Y(n1730) );
  MXI2X1 U767 ( .A(n1603), .B(n1604), .S0(n2061), .Y(N80) );
  MX4X1 U768 ( .A(n1740), .B(n1738), .C(n1739), .D(n1737), .S0(n2063), .S1(
        n2067), .Y(n1603) );
  MX4X1 U769 ( .A(n1736), .B(n1734), .C(n1735), .D(n1733), .S0(n2063), .S1(
        n2067), .Y(n1604) );
  MXI4X1 U770 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n2099), .S1(n2073), 
        .Y(n1738) );
  MXI2X1 U771 ( .A(n1605), .B(n1606), .S0(n2061), .Y(N79) );
  MX4X1 U772 ( .A(n1748), .B(n1746), .C(n1747), .D(n1745), .S0(n2063), .S1(
        n2067), .Y(n1605) );
  MX4X1 U773 ( .A(n1744), .B(n1742), .C(n1743), .D(n1741), .S0(n2063), .S1(
        n2067), .Y(n1606) );
  MXI4X1 U774 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n2100), .S1(n2078), 
        .Y(n1746) );
  MXI2X1 U775 ( .A(n1607), .B(n1608), .S0(n2061), .Y(N78) );
  MX4X1 U776 ( .A(n1756), .B(n1754), .C(n1755), .D(n1753), .S0(n2063), .S1(
        n2067), .Y(n1607) );
  MX4X1 U777 ( .A(n1752), .B(n1750), .C(n1751), .D(n1749), .S0(n2063), .S1(
        n2067), .Y(n1608) );
  MXI4X1 U778 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1754) );
  MXI2X1 U779 ( .A(n1609), .B(n1610), .S0(n2061), .Y(N77) );
  MX4X1 U780 ( .A(n1764), .B(n1762), .C(n1763), .D(n1761), .S0(n2064), .S1(
        n2068), .Y(n1609) );
  MX4X1 U781 ( .A(n1760), .B(n1758), .C(n1759), .D(n1757), .S0(n2064), .S1(
        n2068), .Y(n1610) );
  MXI4X1 U782 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n2101), .S1(n2078), 
        .Y(n1762) );
  MXI2X1 U783 ( .A(n1611), .B(n1612), .S0(n2061), .Y(N76) );
  MX4X1 U784 ( .A(n1772), .B(n1770), .C(n1771), .D(n1769), .S0(n2064), .S1(
        n2068), .Y(n1611) );
  MX4X1 U785 ( .A(n1768), .B(n1766), .C(n1767), .D(n1765), .S0(n2064), .S1(
        n2068), .Y(n1612) );
  MXI4X1 U786 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n2101), .S1(n2079), 
        .Y(n1770) );
  MXI2X1 U787 ( .A(n1613), .B(n1614), .S0(n2061), .Y(N75) );
  MX4X1 U788 ( .A(n1776), .B(n1774), .C(n1775), .D(n1773), .S0(n2064), .S1(
        n2068), .Y(n1614) );
  MX4X1 U789 ( .A(n1780), .B(n1778), .C(n1779), .D(n1777), .S0(n2064), .S1(
        n2068), .Y(n1613) );
  MXI4X1 U790 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1776) );
  MXI2X1 U791 ( .A(n1615), .B(n1616), .S0(n2061), .Y(N74) );
  MX4X1 U792 ( .A(n1784), .B(n1782), .C(n1783), .D(n1781), .S0(n2064), .S1(
        n2068), .Y(n1616) );
  MX4X1 U793 ( .A(n1788), .B(n1786), .C(n1787), .D(n1785), .S0(n2064), .S1(
        n2068), .Y(n1615) );
  MXI4X1 U794 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1784) );
  MXI2X1 U795 ( .A(n1617), .B(n1618), .S0(n2061), .Y(N73) );
  MX4X1 U796 ( .A(n1792), .B(n1790), .C(n1791), .D(n1789), .S0(n2064), .S1(
        n2068), .Y(n1618) );
  MX4X1 U797 ( .A(n1796), .B(n1794), .C(n1795), .D(n1793), .S0(n2064), .S1(
        n2068), .Y(n1617) );
  MXI4X1 U798 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n2088), .S1(n2070), 
        .Y(n1792) );
  MXI2X1 U799 ( .A(n1619), .B(n1620), .S0(n2061), .Y(N72) );
  MX4X1 U800 ( .A(n1800), .B(n1798), .C(n1799), .D(n1797), .S0(n2064), .S1(
        n2068), .Y(n1620) );
  MX4X1 U801 ( .A(n1804), .B(n1802), .C(n1803), .D(n1801), .S0(n2064), .S1(
        n2068), .Y(n1619) );
  MXI4X1 U802 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n2088), .S1(n2071), 
        .Y(n1800) );
  MXI2X1 U803 ( .A(n1621), .B(n1622), .S0(N21), .Y(N71) );
  MX4X1 U804 ( .A(n1808), .B(n1806), .C(n1807), .D(n1805), .S0(n2065), .S1(N19), .Y(n1622) );
  MX4X1 U805 ( .A(n1812), .B(n1810), .C(n1811), .D(n1809), .S0(n2065), .S1(
        n2068), .Y(n1621) );
  MXI4X1 U806 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n2089), .S1(n2071), 
        .Y(n1808) );
  MXI2X1 U807 ( .A(n1623), .B(n1624), .S0(N21), .Y(N70) );
  MX4X1 U808 ( .A(n1816), .B(n1814), .C(n1815), .D(n1813), .S0(n2065), .S1(N19), .Y(n1624) );
  MX4X1 U809 ( .A(n1820), .B(n1818), .C(n1819), .D(n1817), .S0(n2065), .S1(
        n2068), .Y(n1623) );
  MXI4X1 U810 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1816) );
  MXI2X1 U811 ( .A(n1625), .B(n1626), .S0(N21), .Y(N69) );
  MX4X1 U812 ( .A(n1824), .B(n1822), .C(n1823), .D(n1821), .S0(n2065), .S1(N19), .Y(n1626) );
  MX4X1 U813 ( .A(n1828), .B(n1826), .C(n1827), .D(n1825), .S0(n2065), .S1(
        n2068), .Y(n1625) );
  MXI4X1 U814 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n2090), .S1(n2072), 
        .Y(n1824) );
  MXI2X1 U815 ( .A(n1627), .B(n1628), .S0(N21), .Y(N68) );
  MX4X1 U816 ( .A(n1832), .B(n1830), .C(n1831), .D(n1829), .S0(n2065), .S1(N19), .Y(n1628) );
  MX4X1 U817 ( .A(n1836), .B(n1834), .C(n1835), .D(n1833), .S0(n2065), .S1(
        n2066), .Y(n1627) );
  MXI4X1 U818 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1832) );
  MXI2X1 U819 ( .A(n1629), .B(n1630), .S0(N21), .Y(N67) );
  MX4X1 U820 ( .A(n1840), .B(n1838), .C(n1839), .D(n1837), .S0(n2065), .S1(N19), .Y(n1630) );
  MX4X1 U821 ( .A(n1844), .B(n1842), .C(n1843), .D(n1841), .S0(n2065), .S1(
        n2069), .Y(n1629) );
  MXI4X1 U822 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n2091), .S1(n2072), 
        .Y(n1840) );
  MXI2X1 U823 ( .A(n1631), .B(n1632), .S0(n2270), .Y(N66) );
  MX4X1 U824 ( .A(n1848), .B(n1846), .C(n1847), .D(n1845), .S0(n2065), .S1(N19), .Y(n1632) );
  MX4X1 U825 ( .A(n1852), .B(n1850), .C(n1851), .D(n1849), .S0(n2065), .S1(N19), .Y(n1631) );
  MXI4X1 U826 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n2091), .S1(n2073), 
        .Y(n1848) );
  MXI2X1 U827 ( .A(n1633), .B(n1634), .S0(N21), .Y(N65) );
  MX4X1 U828 ( .A(n1856), .B(n1854), .C(n1855), .D(n1853), .S0(N20), .S1(n2069), .Y(n1634) );
  MX4X1 U829 ( .A(n1860), .B(n1858), .C(n1859), .D(n1857), .S0(n2065), .S1(
        n2069), .Y(n1633) );
  MXI4X1 U830 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n2091), .S1(n2073), 
        .Y(n1856) );
  MXI2X1 U831 ( .A(n1635), .B(n1636), .S0(N21), .Y(N64) );
  MX4X1 U832 ( .A(n1864), .B(n1862), .C(n1863), .D(n1861), .S0(N20), .S1(n2069), .Y(n1636) );
  MX4X1 U833 ( .A(n1868), .B(n1866), .C(n1867), .D(n1865), .S0(n2269), .S1(
        n2069), .Y(n1635) );
  MXI4X1 U834 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1864) );
  MXI2X1 U835 ( .A(n1637), .B(n1638), .S0(N21), .Y(N63) );
  MX4X1 U836 ( .A(n1872), .B(n1870), .C(n1871), .D(n1869), .S0(N20), .S1(n2069), .Y(n1638) );
  MX4X1 U837 ( .A(n1876), .B(n1874), .C(n1875), .D(n1873), .S0(N20), .S1(n2069), .Y(n1637) );
  MXI4X1 U838 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n2092), .S1(n2074), 
        .Y(n1872) );
  MXI2X1 U839 ( .A(n1639), .B(n1640), .S0(N21), .Y(N62) );
  MX4X1 U840 ( .A(n1880), .B(n1878), .C(n1879), .D(n1877), .S0(N20), .S1(n2069), .Y(n1640) );
  MX4X1 U841 ( .A(n1884), .B(n1882), .C(n1883), .D(n1881), .S0(n2269), .S1(
        n2069), .Y(n1639) );
  MXI4X1 U842 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1880) );
  MXI2X1 U843 ( .A(n1641), .B(n1642), .S0(N21), .Y(N61) );
  MX4X1 U844 ( .A(n1888), .B(n1886), .C(n1887), .D(n1885), .S0(N20), .S1(n2069), .Y(n1642) );
  MX4X1 U845 ( .A(n1892), .B(n1890), .C(n1891), .D(n1889), .S0(n2269), .S1(
        n2069), .Y(n1641) );
  MXI4X1 U846 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1888) );
  MXI2X1 U847 ( .A(n1643), .B(n1644), .S0(N21), .Y(N60) );
  MX4X1 U848 ( .A(n1896), .B(n1894), .C(n1895), .D(n1893), .S0(N20), .S1(n2069), .Y(n1644) );
  MX4X1 U849 ( .A(n1900), .B(n1898), .C(n1899), .D(n1897), .S0(N20), .S1(n2069), .Y(n1643) );
  MXI4X1 U850 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n2094), .S1(n2074), 
        .Y(n1896) );
  MXI2X1 U851 ( .A(n32), .B(n33), .S0(N16), .Y(N56) );
  MX4X1 U852 ( .A(n1121), .B(n1119), .C(n1120), .D(n1118), .S0(n1535), .S1(
        n1540), .Y(n33) );
  MX4X1 U853 ( .A(n1125), .B(n1123), .C(n1124), .D(n1122), .S0(n1535), .S1(
        n1541), .Y(n32) );
  MXI4X1 U854 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1569), .S1(n1550), .Y(
        n1121) );
  MXI2X1 U855 ( .A(n34), .B(n35), .S0(n1534), .Y(N55) );
  MX4X1 U856 ( .A(n1133), .B(n1131), .C(n1132), .D(n1130), .S0(n1535), .S1(
        n1542), .Y(n34) );
  MX4X1 U857 ( .A(n1129), .B(n1127), .C(n1128), .D(n1126), .S0(n1535), .S1(
        n1541), .Y(n35) );
  MXI4X1 U858 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1570), .S1(n1550), .Y(
        n1131) );
  MXI2X1 U859 ( .A(n36), .B(n37), .S0(N16), .Y(N54) );
  MX4X1 U860 ( .A(n1141), .B(n1139), .C(n1140), .D(n1138), .S0(n1536), .S1(
        n1540), .Y(n36) );
  MX4X1 U861 ( .A(n1137), .B(n1135), .C(n1136), .D(n1134), .S0(n1536), .S1(
        n1540), .Y(n37) );
  MXI4X1 U862 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1570), .S1(n1550), .Y(
        n1139) );
  MXI2X1 U863 ( .A(n38), .B(n39), .S0(n1534), .Y(N53) );
  MX4X1 U864 ( .A(n1149), .B(n1147), .C(n1148), .D(n1146), .S0(n1536), .S1(
        n1540), .Y(n38) );
  MX4X1 U865 ( .A(n1145), .B(n1143), .C(n1144), .D(n1142), .S0(n1536), .S1(
        n1540), .Y(n39) );
  MXI4X1 U866 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1571), .S1(n1551), .Y(
        n1147) );
  MXI2X1 U867 ( .A(n40), .B(n41), .S0(N16), .Y(N52) );
  MX4X1 U868 ( .A(n1157), .B(n1155), .C(n1156), .D(n1154), .S0(n1536), .S1(
        n1540), .Y(n40) );
  MX4X1 U869 ( .A(n1153), .B(n1151), .C(n1152), .D(n1150), .S0(n1536), .S1(
        n1540), .Y(n41) );
  MXI4X1 U870 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1571), .S1(n1551), .Y(
        n1155) );
  MXI2X1 U871 ( .A(n42), .B(n43), .S0(n1534), .Y(N51) );
  MX4X1 U872 ( .A(n1165), .B(n1163), .C(n1164), .D(n1162), .S0(n1536), .S1(
        n1540), .Y(n42) );
  MX4X1 U873 ( .A(n1161), .B(n1159), .C(n1160), .D(n1158), .S0(n1536), .S1(
        n1540), .Y(n43) );
  MXI4X1 U874 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1572), .S1(n1551), .Y(
        n1163) );
  MXI2X1 U875 ( .A(n44), .B(n45), .S0(n1534), .Y(N50) );
  MX4X1 U876 ( .A(n1173), .B(n1171), .C(n1172), .D(n1170), .S0(n1536), .S1(
        n1540), .Y(n44) );
  MX4X1 U877 ( .A(n1169), .B(n1167), .C(n1168), .D(n1166), .S0(n1536), .S1(
        n1540), .Y(n45) );
  MXI4X1 U878 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1572), .S1(n1550), .Y(
        n1171) );
  MXI2X1 U879 ( .A(n46), .B(n65), .S0(n2271), .Y(N49) );
  MX4X1 U880 ( .A(n1181), .B(n1179), .C(n1180), .D(n1178), .S0(n1536), .S1(
        n1540), .Y(n46) );
  MX4X1 U881 ( .A(n1177), .B(n1175), .C(n1176), .D(n1174), .S0(n1536), .S1(
        n1540), .Y(n65) );
  MXI4X1 U882 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1573), .S1(n1544), .Y(
        n1179) );
  MXI2X1 U883 ( .A(n68), .B(n70), .S0(n1534), .Y(N48) );
  MX4X1 U884 ( .A(n1189), .B(n1187), .C(n1188), .D(n1186), .S0(n1536), .S1(
        n1542), .Y(n68) );
  MX4X1 U885 ( .A(n1185), .B(n1183), .C(n1184), .D(n1182), .S0(N15), .S1(n1542), .Y(n70) );
  MXI4X1 U886 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1573), .S1(n1545), .Y(
        n1187) );
  MXI2X1 U887 ( .A(n72), .B(n74), .S0(n1534), .Y(N47) );
  MX4X1 U888 ( .A(n1197), .B(n1195), .C(n1196), .D(n1194), .S0(n1535), .S1(
        n1541), .Y(n72) );
  MX4X1 U889 ( .A(n1193), .B(n1191), .C(n1192), .D(n1190), .S0(n1538), .S1(
        n1540), .Y(n74) );
  MXI4X1 U890 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1574), .S1(n1544), .Y(
        n1195) );
  MXI2X1 U891 ( .A(n76), .B(n78), .S0(n1534), .Y(N46) );
  MX4X1 U892 ( .A(n1205), .B(n1203), .C(n1204), .D(n1202), .S0(n1535), .S1(
        n1543), .Y(n76) );
  MX4X1 U893 ( .A(n1201), .B(n1199), .C(n1200), .D(n1198), .S0(n1535), .S1(
        n1543), .Y(n78) );
  MXI4X1 U894 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1574), .S1(n1556), 
        .Y(n1203) );
  MXI2X1 U895 ( .A(n80), .B(n83), .S0(n1534), .Y(N45) );
  MX4X1 U896 ( .A(n1213), .B(n1211), .C(n1212), .D(n1210), .S0(n1535), .S1(
        n1543), .Y(n80) );
  MX4X1 U897 ( .A(n1209), .B(n1207), .C(n1208), .D(n1206), .S0(n1535), .S1(
        n1541), .Y(n83) );
  MXI4X1 U898 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1574), .S1(n1545), 
        .Y(n1211) );
  MXI2X1 U899 ( .A(n84), .B(n85), .S0(n1534), .Y(N44) );
  MX4X1 U900 ( .A(n1221), .B(n1219), .C(n1220), .D(n1218), .S0(n1535), .S1(
        n1543), .Y(n84) );
  MX4X1 U901 ( .A(n1217), .B(n1215), .C(n1216), .D(n1214), .S0(n1535), .S1(
        n1540), .Y(n85) );
  MXI4X1 U902 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1575), .S1(n1544), 
        .Y(n1219) );
  MXI2X1 U903 ( .A(n86), .B(n87), .S0(n1534), .Y(N43) );
  MX4X1 U904 ( .A(n1229), .B(n1227), .C(n1228), .D(n1226), .S0(n1535), .S1(
        n1542), .Y(n86) );
  MX4X1 U905 ( .A(n1225), .B(n1223), .C(n1224), .D(n1222), .S0(n1535), .S1(
        n1540), .Y(n87) );
  MXI4X1 U906 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1575), .S1(n1546), 
        .Y(n1227) );
  MXI2X1 U907 ( .A(n88), .B(n89), .S0(n1534), .Y(N42) );
  MX4X1 U908 ( .A(n1237), .B(n1235), .C(n1236), .D(n1234), .S0(n1537), .S1(
        n1541), .Y(n88) );
  MX4X1 U909 ( .A(n1233), .B(n1231), .C(n1232), .D(n1230), .S0(n1537), .S1(
        n1541), .Y(n89) );
  MXI4X1 U910 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1576), .S1(n1556), 
        .Y(n1235) );
  MXI2X1 U911 ( .A(n90), .B(n92), .S0(n1534), .Y(N41) );
  MX4X1 U912 ( .A(n1245), .B(n1243), .C(n1244), .D(n1242), .S0(n1537), .S1(
        n1541), .Y(n90) );
  MX4X1 U913 ( .A(n1241), .B(n1239), .C(n1240), .D(n1238), .S0(n1537), .S1(
        n1541), .Y(n92) );
  MXI4X1 U914 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1576), .S1(n1552), 
        .Y(n1243) );
  MXI2X1 U915 ( .A(n93), .B(n94), .S0(n1534), .Y(N40) );
  MX4X1 U916 ( .A(n1249), .B(n1247), .C(n1248), .D(n1246), .S0(n1537), .S1(
        n1541), .Y(n94) );
  MX4X1 U917 ( .A(n1253), .B(n1251), .C(n1252), .D(n1250), .S0(n1537), .S1(
        n1541), .Y(n93) );
  MXI4X1 U918 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1249) );
  MXI2X1 U919 ( .A(n95), .B(n96), .S0(n1534), .Y(N39) );
  MX4X1 U920 ( .A(n1257), .B(n1255), .C(n1256), .D(n1254), .S0(n1537), .S1(
        n1541), .Y(n96) );
  MX4X1 U921 ( .A(n1261), .B(n1259), .C(n1260), .D(n1258), .S0(n1537), .S1(
        n1541), .Y(n95) );
  MXI4X1 U922 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1257) );
  MXI2X1 U923 ( .A(n97), .B(n98), .S0(n1534), .Y(N38) );
  MX4X1 U924 ( .A(n1265), .B(n1263), .C(n1264), .D(n1262), .S0(n1537), .S1(
        n1541), .Y(n98) );
  MX4X1 U925 ( .A(n1269), .B(n1267), .C(n1268), .D(n1266), .S0(n1537), .S1(
        n1541), .Y(n97) );
  MXI4X1 U926 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1563), .S1(n1546), 
        .Y(n1265) );
  MXI2X1 U927 ( .A(n99), .B(n101), .S0(n1534), .Y(N37) );
  MX4X1 U928 ( .A(n1273), .B(n1271), .C(n1272), .D(n1270), .S0(n1537), .S1(
        n1541), .Y(n101) );
  MX4X1 U929 ( .A(n1277), .B(n1275), .C(n1276), .D(n1274), .S0(n1537), .S1(
        n1541), .Y(n99) );
  MXI4X1 U930 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1563), .S1(n1555), 
        .Y(n1273) );
  MXI2X1 U931 ( .A(n102), .B(n103), .S0(n1534), .Y(N36) );
  MX4X1 U932 ( .A(n1281), .B(n1279), .C(n1280), .D(n1278), .S0(n1538), .S1(
        n1542), .Y(n103) );
  MX4X1 U933 ( .A(n1285), .B(n1283), .C(n1284), .D(n1282), .S0(n1538), .S1(
        n1542), .Y(n102) );
  MXI4X1 U934 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1564), .S1(n1544), 
        .Y(n1281) );
  MXI2X1 U935 ( .A(n104), .B(n105), .S0(N16), .Y(N35) );
  MX4X1 U936 ( .A(n1289), .B(n1287), .C(n1288), .D(n1286), .S0(n1538), .S1(
        n1542), .Y(n105) );
  MX4X1 U937 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1538), .S1(
        n1542), .Y(n104) );
  MXI4X1 U938 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1564), .S1(n1544), 
        .Y(n1289) );
  MXI2X1 U939 ( .A(n106), .B(n107), .S0(N16), .Y(N34) );
  MX4X1 U940 ( .A(n1297), .B(n1295), .C(n1296), .D(n1294), .S0(n1538), .S1(
        n1542), .Y(n107) );
  MX4X1 U941 ( .A(n1301), .B(n1299), .C(n1300), .D(n1298), .S0(n1538), .S1(
        n1542), .Y(n106) );
  MXI4X1 U942 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1565), .S1(n1547), 
        .Y(n1297) );
  MXI2X1 U943 ( .A(n1100), .B(n1101), .S0(N16), .Y(N33) );
  MX4X1 U944 ( .A(n1305), .B(n1303), .C(n1304), .D(n1302), .S0(n1538), .S1(
        n1542), .Y(n1101) );
  MX4X1 U945 ( .A(n1309), .B(n1307), .C(n1308), .D(n1306), .S0(n1538), .S1(
        n1542), .Y(n1100) );
  MXI4X1 U946 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1305) );
  MXI2X1 U947 ( .A(n1102), .B(n1103), .S0(N16), .Y(N32) );
  MX4X1 U948 ( .A(n1313), .B(n1311), .C(n1312), .D(n1310), .S0(n1538), .S1(
        n1542), .Y(n1103) );
  MX4X1 U949 ( .A(n1317), .B(n1315), .C(n1316), .D(n1314), .S0(n1538), .S1(
        n1542), .Y(n1102) );
  MXI4X1 U950 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1566), .S1(n1547), 
        .Y(n1313) );
  MXI2X1 U951 ( .A(n1104), .B(n1105), .S0(N16), .Y(N31) );
  MX4X1 U952 ( .A(n1321), .B(n1319), .C(n1320), .D(n1318), .S0(n1538), .S1(
        n1542), .Y(n1105) );
  MX4X1 U953 ( .A(n1325), .B(n1323), .C(n1324), .D(n1322), .S0(n1538), .S1(
        n1542), .Y(n1104) );
  MXI4X1 U954 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1566), .S1(n1548), 
        .Y(n1321) );
  MXI2X1 U955 ( .A(n1106), .B(n1107), .S0(N16), .Y(N30) );
  MX4X1 U956 ( .A(n1329), .B(n1327), .C(n1328), .D(n1326), .S0(n1539), .S1(
        n1543), .Y(n1107) );
  MX4X1 U957 ( .A(n1333), .B(n1331), .C(n1332), .D(n1330), .S0(n1539), .S1(
        n1543), .Y(n1106) );
  MXI4X1 U958 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1566), .S1(n1548), 
        .Y(n1329) );
  MXI2X1 U959 ( .A(n1108), .B(n1109), .S0(N16), .Y(N29) );
  MX4X1 U960 ( .A(n1337), .B(n1335), .C(n1336), .D(n1334), .S0(n1539), .S1(
        n1543), .Y(n1109) );
  MX4X1 U961 ( .A(n1341), .B(n1339), .C(n1340), .D(n1338), .S0(n1539), .S1(
        n1543), .Y(n1108) );
  MXI4X1 U962 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1337) );
  MXI2X1 U963 ( .A(n1110), .B(n1111), .S0(N16), .Y(N28) );
  MX4X1 U964 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1539), .S1(
        n1543), .Y(n1111) );
  MX4X1 U965 ( .A(n1349), .B(n1347), .C(n1348), .D(n1346), .S0(n1539), .S1(
        n1543), .Y(n1110) );
  MXI4X1 U966 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1567), .S1(n1549), 
        .Y(n1345) );
  MXI2X1 U967 ( .A(n1112), .B(n1113), .S0(N16), .Y(N27) );
  MX4X1 U968 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1539), .S1(
        n1543), .Y(n1113) );
  MX4X1 U969 ( .A(n1357), .B(n1355), .C(n1356), .D(n1354), .S0(n1539), .S1(
        n1543), .Y(n1112) );
  MXI4X1 U970 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1353) );
  MXI2X1 U971 ( .A(n1114), .B(n1115), .S0(N16), .Y(N26) );
  MX4X1 U972 ( .A(n1361), .B(n1359), .C(n1360), .D(n1358), .S0(n1539), .S1(
        n1543), .Y(n1115) );
  MX4X1 U973 ( .A(n1365), .B(n1363), .C(n1364), .D(n1362), .S0(n1539), .S1(
        n1543), .Y(n1114) );
  MXI4X1 U974 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1361) );
  MXI2X1 U975 ( .A(n1116), .B(n1117), .S0(N16), .Y(N25) );
  MX4X1 U976 ( .A(n1369), .B(n1367), .C(n1368), .D(n1366), .S0(n1539), .S1(
        n1543), .Y(n1117) );
  MX4X1 U977 ( .A(n1373), .B(n1371), .C(n1372), .D(n1370), .S0(n1539), .S1(
        n1543), .Y(n1116) );
  MXI4X1 U978 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1569), .S1(n1549), 
        .Y(n1369) );
  OAI2BB2XL U979 ( .B0(n2121), .B1(n2256), .A0N(\register[2][23] ), .A1N(n2258), .Y(n163) );
  OAI2BB2XL U980 ( .B0(n2424), .B1(n26), .A0N(\register[2][25] ), .A1N(n2258), 
        .Y(n165) );
  OAI2BB2XL U981 ( .B0(n2115), .B1(n2257), .A0N(\register[2][26] ), .A1N(n2258), .Y(n166) );
  OAI2BB2XL U982 ( .B0(n2113), .B1(n2256), .A0N(\register[2][27] ), .A1N(n2258), .Y(n167) );
  OAI2BB2XL U983 ( .B0(n2111), .B1(n2257), .A0N(\register[2][28] ), .A1N(n2258), .Y(n168) );
  OAI2BB2XL U984 ( .B0(n2109), .B1(n26), .A0N(\register[2][29] ), .A1N(n2258), 
        .Y(n169) );
  OAI2BB2XL U985 ( .B0(n2107), .B1(n26), .A0N(\register[2][30] ), .A1N(n2256), 
        .Y(n170) );
  OAI2BB2XL U986 ( .B0(n2105), .B1(n26), .A0N(\register[2][31] ), .A1N(n2257), 
        .Y(n171) );
  OAI2BB2XL U987 ( .B0(n2121), .B1(n2253), .A0N(\register[3][23] ), .A1N(n2255), .Y(n195) );
  OAI2BB2XL U988 ( .B0(n2424), .B1(n27), .A0N(\register[3][25] ), .A1N(n2255), 
        .Y(n197) );
  OAI2BB2XL U989 ( .B0(n2115), .B1(n2254), .A0N(\register[3][26] ), .A1N(n2255), .Y(n198) );
  OAI2BB2XL U990 ( .B0(n2113), .B1(n2253), .A0N(\register[3][27] ), .A1N(n2255), .Y(n199) );
  OAI2BB2XL U991 ( .B0(n2111), .B1(n2254), .A0N(\register[3][28] ), .A1N(n2255), .Y(n200) );
  OAI2BB2XL U992 ( .B0(n2109), .B1(n27), .A0N(\register[3][29] ), .A1N(n2255), 
        .Y(n201) );
  OAI2BB2XL U993 ( .B0(n2107), .B1(n27), .A0N(\register[3][30] ), .A1N(n2253), 
        .Y(n202) );
  OAI2BB2XL U994 ( .B0(n2105), .B1(n27), .A0N(\register[3][31] ), .A1N(n2254), 
        .Y(n203) );
  OAI2BB2XL U995 ( .B0(n2121), .B1(n2250), .A0N(\register[4][23] ), .A1N(n2252), .Y(n227) );
  OAI2BB2XL U996 ( .B0(n2118), .B1(n28), .A0N(\register[4][25] ), .A1N(n2252), 
        .Y(n229) );
  OAI2BB2XL U997 ( .B0(n2115), .B1(n2251), .A0N(\register[4][26] ), .A1N(n2252), .Y(n230) );
  OAI2BB2XL U998 ( .B0(n2113), .B1(n2250), .A0N(\register[4][27] ), .A1N(n2252), .Y(n231) );
  OAI2BB2XL U999 ( .B0(n2111), .B1(n2251), .A0N(\register[4][28] ), .A1N(n2252), .Y(n232) );
  OAI2BB2XL U1000 ( .B0(n2109), .B1(n28), .A0N(\register[4][29] ), .A1N(n2252), 
        .Y(n233) );
  OAI2BB2XL U1001 ( .B0(n2107), .B1(n28), .A0N(\register[4][30] ), .A1N(n2250), 
        .Y(n234) );
  OAI2BB2XL U1002 ( .B0(n2105), .B1(n28), .A0N(\register[4][31] ), .A1N(n2251), 
        .Y(n235) );
  OAI2BB2XL U1003 ( .B0(n2121), .B1(n2247), .A0N(\register[5][23] ), .A1N(
        n2249), .Y(n259) );
  OAI2BB2XL U1004 ( .B0(n2117), .B1(n29), .A0N(\register[5][25] ), .A1N(n2249), 
        .Y(n261) );
  OAI2BB2XL U1005 ( .B0(n2115), .B1(n2248), .A0N(\register[5][26] ), .A1N(
        n2249), .Y(n262) );
  OAI2BB2XL U1006 ( .B0(n2113), .B1(n2247), .A0N(\register[5][27] ), .A1N(
        n2249), .Y(n263) );
  OAI2BB2XL U1007 ( .B0(n2111), .B1(n2248), .A0N(\register[5][28] ), .A1N(
        n2249), .Y(n264) );
  OAI2BB2XL U1008 ( .B0(n2109), .B1(n29), .A0N(\register[5][29] ), .A1N(n2249), 
        .Y(n265) );
  OAI2BB2XL U1009 ( .B0(n2107), .B1(n29), .A0N(\register[5][30] ), .A1N(n2247), 
        .Y(n266) );
  OAI2BB2XL U1010 ( .B0(n2105), .B1(n29), .A0N(\register[5][31] ), .A1N(n2248), 
        .Y(n267) );
  OAI2BB2XL U1011 ( .B0(n2121), .B1(n2244), .A0N(\register[6][23] ), .A1N(
        n2246), .Y(n291) );
  OAI2BB2XL U1012 ( .B0(n2118), .B1(n30), .A0N(\register[6][25] ), .A1N(n2246), 
        .Y(n293) );
  OAI2BB2XL U1013 ( .B0(n2115), .B1(n2245), .A0N(\register[6][26] ), .A1N(
        n2246), .Y(n294) );
  OAI2BB2XL U1014 ( .B0(n2113), .B1(n2244), .A0N(\register[6][27] ), .A1N(
        n2246), .Y(n295) );
  OAI2BB2XL U1015 ( .B0(n2111), .B1(n2245), .A0N(\register[6][28] ), .A1N(
        n2246), .Y(n296) );
  OAI2BB2XL U1016 ( .B0(n2109), .B1(n30), .A0N(\register[6][29] ), .A1N(n2246), 
        .Y(n297) );
  OAI2BB2XL U1017 ( .B0(n2107), .B1(n30), .A0N(\register[6][30] ), .A1N(n2244), 
        .Y(n298) );
  OAI2BB2XL U1018 ( .B0(n2105), .B1(n30), .A0N(\register[6][31] ), .A1N(n2245), 
        .Y(n299) );
  OAI2BB2XL U1019 ( .B0(n2121), .B1(n2241), .A0N(\register[7][23] ), .A1N(
        n2243), .Y(n323) );
  OAI2BB2XL U1020 ( .B0(n2117), .B1(n31), .A0N(\register[7][25] ), .A1N(n2243), 
        .Y(n325) );
  OAI2BB2XL U1021 ( .B0(n2115), .B1(n2242), .A0N(\register[7][26] ), .A1N(
        n2243), .Y(n326) );
  OAI2BB2XL U1022 ( .B0(n2113), .B1(n2241), .A0N(\register[7][27] ), .A1N(
        n2243), .Y(n327) );
  OAI2BB2XL U1023 ( .B0(n2111), .B1(n2242), .A0N(\register[7][28] ), .A1N(
        n2243), .Y(n328) );
  OAI2BB2XL U1024 ( .B0(n2109), .B1(n31), .A0N(\register[7][29] ), .A1N(n2243), 
        .Y(n329) );
  OAI2BB2XL U1025 ( .B0(n2107), .B1(n31), .A0N(\register[7][30] ), .A1N(n2241), 
        .Y(n330) );
  OAI2BB2XL U1026 ( .B0(n2105), .B1(n31), .A0N(\register[7][31] ), .A1N(n2242), 
        .Y(n331) );
  OAI2BB2XL U1027 ( .B0(n2122), .B1(n2239), .A0N(\register[8][23] ), .A1N(
        n2238), .Y(n355) );
  OAI2BB2XL U1028 ( .B0(n2118), .B1(n2238), .A0N(\register[8][25] ), .A1N(
        n2240), .Y(n357) );
  OAI2BB2XL U1029 ( .B0(n2116), .B1(n2239), .A0N(\register[8][26] ), .A1N(
        n2240), .Y(n358) );
  OAI2BB2XL U1030 ( .B0(n2114), .B1(n2238), .A0N(\register[8][27] ), .A1N(
        n2240), .Y(n359) );
  OAI2BB2XL U1031 ( .B0(n2112), .B1(n12), .A0N(\register[8][28] ), .A1N(n2240), 
        .Y(n360) );
  OAI2BB2XL U1032 ( .B0(n2110), .B1(n12), .A0N(\register[8][29] ), .A1N(n2240), 
        .Y(n361) );
  OAI2BB2XL U1033 ( .B0(n2108), .B1(n12), .A0N(\register[8][30] ), .A1N(n2238), 
        .Y(n362) );
  OAI2BB2XL U1034 ( .B0(n2106), .B1(n12), .A0N(\register[8][31] ), .A1N(n2239), 
        .Y(n363) );
  OAI2BB2XL U1035 ( .B0(n2122), .B1(n2233), .A0N(\register[10][23] ), .A1N(
        n2232), .Y(n419) );
  OAI2BB2XL U1036 ( .B0(n2118), .B1(n2232), .A0N(\register[10][25] ), .A1N(
        n2234), .Y(n421) );
  OAI2BB2XL U1037 ( .B0(n2116), .B1(n2233), .A0N(\register[10][26] ), .A1N(
        n2234), .Y(n422) );
  OAI2BB2XL U1038 ( .B0(n2114), .B1(n2232), .A0N(\register[10][27] ), .A1N(
        n2234), .Y(n423) );
  OAI2BB2XL U1039 ( .B0(n2112), .B1(n13), .A0N(\register[10][28] ), .A1N(n2234), .Y(n424) );
  OAI2BB2XL U1040 ( .B0(n2110), .B1(n13), .A0N(\register[10][29] ), .A1N(n2234), .Y(n425) );
  OAI2BB2XL U1041 ( .B0(n2108), .B1(n13), .A0N(\register[10][30] ), .A1N(n2232), .Y(n426) );
  OAI2BB2XL U1042 ( .B0(n2106), .B1(n13), .A0N(\register[10][31] ), .A1N(n2233), .Y(n427) );
  OAI2BB2XL U1043 ( .B0(n2122), .B1(n2230), .A0N(\register[11][23] ), .A1N(
        n2229), .Y(n451) );
  OAI2BB2XL U1044 ( .B0(n2118), .B1(n2229), .A0N(\register[11][25] ), .A1N(
        n2231), .Y(n453) );
  OAI2BB2XL U1045 ( .B0(n2116), .B1(n2230), .A0N(\register[11][26] ), .A1N(
        n2231), .Y(n454) );
  OAI2BB2XL U1046 ( .B0(n2114), .B1(n2229), .A0N(\register[11][27] ), .A1N(
        n2231), .Y(n455) );
  OAI2BB2XL U1047 ( .B0(n2112), .B1(n14), .A0N(\register[11][28] ), .A1N(n2231), .Y(n456) );
  OAI2BB2XL U1048 ( .B0(n2110), .B1(n14), .A0N(\register[11][29] ), .A1N(n2231), .Y(n457) );
  OAI2BB2XL U1049 ( .B0(n2108), .B1(n14), .A0N(\register[11][30] ), .A1N(n2229), .Y(n458) );
  OAI2BB2XL U1050 ( .B0(n2106), .B1(n14), .A0N(\register[11][31] ), .A1N(n2230), .Y(n459) );
  OAI2BB2XL U1051 ( .B0(n2122), .B1(n2227), .A0N(\register[12][23] ), .A1N(
        n2226), .Y(n483) );
  OAI2BB2XL U1052 ( .B0(n2118), .B1(n2226), .A0N(\register[12][25] ), .A1N(
        n2228), .Y(n485) );
  OAI2BB2XL U1053 ( .B0(n2116), .B1(n2227), .A0N(\register[12][26] ), .A1N(
        n2228), .Y(n486) );
  OAI2BB2XL U1054 ( .B0(n2114), .B1(n2226), .A0N(\register[12][27] ), .A1N(
        n2228), .Y(n487) );
  OAI2BB2XL U1055 ( .B0(n2112), .B1(n15), .A0N(\register[12][28] ), .A1N(n2228), .Y(n488) );
  OAI2BB2XL U1056 ( .B0(n2110), .B1(n15), .A0N(\register[12][29] ), .A1N(n2228), .Y(n489) );
  OAI2BB2XL U1057 ( .B0(n2108), .B1(n15), .A0N(\register[12][30] ), .A1N(n2226), .Y(n490) );
  OAI2BB2XL U1058 ( .B0(n2106), .B1(n15), .A0N(\register[12][31] ), .A1N(n2227), .Y(n491) );
  OAI2BB2XL U1059 ( .B0(n2122), .B1(n2224), .A0N(\register[13][23] ), .A1N(
        n2223), .Y(n515) );
  OAI2BB2XL U1060 ( .B0(n2118), .B1(n2223), .A0N(\register[13][25] ), .A1N(
        n2225), .Y(n517) );
  OAI2BB2XL U1061 ( .B0(n2116), .B1(n2224), .A0N(\register[13][26] ), .A1N(
        n2225), .Y(n518) );
  OAI2BB2XL U1062 ( .B0(n2114), .B1(n2223), .A0N(\register[13][27] ), .A1N(
        n2225), .Y(n519) );
  OAI2BB2XL U1063 ( .B0(n2112), .B1(n16), .A0N(\register[13][28] ), .A1N(n2225), .Y(n520) );
  OAI2BB2XL U1064 ( .B0(n2110), .B1(n16), .A0N(\register[13][29] ), .A1N(n2225), .Y(n521) );
  OAI2BB2XL U1065 ( .B0(n2108), .B1(n16), .A0N(\register[13][30] ), .A1N(n2223), .Y(n522) );
  OAI2BB2XL U1066 ( .B0(n2106), .B1(n16), .A0N(\register[13][31] ), .A1N(n2224), .Y(n523) );
  OAI2BB2XL U1067 ( .B0(n2122), .B1(n2221), .A0N(\register[14][23] ), .A1N(
        n2220), .Y(n547) );
  OAI2BB2XL U1068 ( .B0(n2118), .B1(n2220), .A0N(\register[14][25] ), .A1N(
        n2222), .Y(n549) );
  OAI2BB2XL U1069 ( .B0(n2116), .B1(n2221), .A0N(\register[14][26] ), .A1N(
        n2222), .Y(n550) );
  OAI2BB2XL U1070 ( .B0(n2114), .B1(n2220), .A0N(\register[14][27] ), .A1N(
        n2222), .Y(n551) );
  OAI2BB2XL U1071 ( .B0(n2112), .B1(n17), .A0N(\register[14][28] ), .A1N(n2222), .Y(n552) );
  OAI2BB2XL U1072 ( .B0(n2110), .B1(n17), .A0N(\register[14][29] ), .A1N(n2222), .Y(n553) );
  OAI2BB2XL U1073 ( .B0(n2108), .B1(n17), .A0N(\register[14][30] ), .A1N(n2220), .Y(n554) );
  OAI2BB2XL U1074 ( .B0(n2106), .B1(n17), .A0N(\register[14][31] ), .A1N(n2221), .Y(n555) );
  OAI2BB2XL U1075 ( .B0(n2122), .B1(n2218), .A0N(\register[15][23] ), .A1N(
        n2217), .Y(n579) );
  OAI2BB2XL U1076 ( .B0(n2118), .B1(n2217), .A0N(\register[15][25] ), .A1N(
        n2219), .Y(n581) );
  OAI2BB2XL U1077 ( .B0(n2116), .B1(n2218), .A0N(\register[15][26] ), .A1N(
        n2219), .Y(n582) );
  OAI2BB2XL U1078 ( .B0(n2114), .B1(n2217), .A0N(\register[15][27] ), .A1N(
        n2219), .Y(n583) );
  OAI2BB2XL U1079 ( .B0(n2112), .B1(n18), .A0N(\register[15][28] ), .A1N(n2219), .Y(n584) );
  OAI2BB2XL U1080 ( .B0(n2110), .B1(n18), .A0N(\register[15][29] ), .A1N(n2219), .Y(n585) );
  OAI2BB2XL U1081 ( .B0(n2108), .B1(n18), .A0N(\register[15][30] ), .A1N(n2217), .Y(n586) );
  OAI2BB2XL U1082 ( .B0(n2106), .B1(n18), .A0N(\register[15][31] ), .A1N(n2218), .Y(n587) );
  OAI2BB2XL U1083 ( .B0(n2122), .B1(n2215), .A0N(\register[16][23] ), .A1N(
        n2214), .Y(n611) );
  OAI2BB2XL U1084 ( .B0(n2118), .B1(n2214), .A0N(\register[16][25] ), .A1N(
        n2216), .Y(n613) );
  OAI2BB2XL U1085 ( .B0(n2116), .B1(n2215), .A0N(\register[16][26] ), .A1N(
        n2216), .Y(n614) );
  OAI2BB2XL U1086 ( .B0(n2114), .B1(n2214), .A0N(\register[16][27] ), .A1N(
        n2216), .Y(n615) );
  OAI2BB2XL U1087 ( .B0(n2112), .B1(n19), .A0N(\register[16][28] ), .A1N(n2216), .Y(n616) );
  OAI2BB2XL U1088 ( .B0(n2110), .B1(n19), .A0N(\register[16][29] ), .A1N(n2216), .Y(n617) );
  OAI2BB2XL U1089 ( .B0(n2108), .B1(n19), .A0N(\register[16][30] ), .A1N(n2214), .Y(n618) );
  OAI2BB2XL U1090 ( .B0(n2106), .B1(n19), .A0N(\register[16][31] ), .A1N(n2215), .Y(n619) );
  OAI2BB2XL U1091 ( .B0(n2122), .B1(n2209), .A0N(\register[18][23] ), .A1N(
        n2208), .Y(n675) );
  OAI2BB2XL U1092 ( .B0(n2118), .B1(n2208), .A0N(\register[18][25] ), .A1N(
        n2210), .Y(n677) );
  OAI2BB2XL U1093 ( .B0(n2116), .B1(n2209), .A0N(\register[18][26] ), .A1N(
        n2210), .Y(n678) );
  OAI2BB2XL U1094 ( .B0(n2114), .B1(n2208), .A0N(\register[18][27] ), .A1N(
        n2210), .Y(n679) );
  OAI2BB2XL U1095 ( .B0(n2112), .B1(n20), .A0N(\register[18][28] ), .A1N(n2210), .Y(n680) );
  OAI2BB2XL U1096 ( .B0(n2110), .B1(n20), .A0N(\register[18][29] ), .A1N(n2210), .Y(n681) );
  OAI2BB2XL U1097 ( .B0(n2108), .B1(n20), .A0N(\register[18][30] ), .A1N(n2208), .Y(n682) );
  OAI2BB2XL U1098 ( .B0(n2106), .B1(n20), .A0N(\register[18][31] ), .A1N(n2209), .Y(n683) );
  OAI2BB2XL U1099 ( .B0(n2122), .B1(n2206), .A0N(\register[19][23] ), .A1N(
        n2205), .Y(n707) );
  OAI2BB2XL U1100 ( .B0(n2118), .B1(n2205), .A0N(\register[19][25] ), .A1N(
        n2207), .Y(n709) );
  OAI2BB2XL U1101 ( .B0(n2116), .B1(n2206), .A0N(\register[19][26] ), .A1N(
        n2207), .Y(n710) );
  OAI2BB2XL U1102 ( .B0(n2114), .B1(n2205), .A0N(\register[19][27] ), .A1N(
        n2207), .Y(n711) );
  OAI2BB2XL U1103 ( .B0(n2112), .B1(n21), .A0N(\register[19][28] ), .A1N(n2207), .Y(n712) );
  OAI2BB2XL U1104 ( .B0(n2110), .B1(n21), .A0N(\register[19][29] ), .A1N(n2207), .Y(n713) );
  OAI2BB2XL U1105 ( .B0(n2108), .B1(n21), .A0N(\register[19][30] ), .A1N(n2205), .Y(n714) );
  OAI2BB2XL U1106 ( .B0(n2106), .B1(n21), .A0N(\register[19][31] ), .A1N(n2206), .Y(n715) );
  OAI2BB2XL U1107 ( .B0(n2121), .B1(n2203), .A0N(\register[20][23] ), .A1N(
        n2204), .Y(n739) );
  OAI2BB2XL U1108 ( .B0(n2117), .B1(n22), .A0N(\register[20][25] ), .A1N(n2204), .Y(n741) );
  OAI2BB2XL U1109 ( .B0(n2115), .B1(n2202), .A0N(\register[20][26] ), .A1N(
        n2204), .Y(n742) );
  OAI2BB2XL U1110 ( .B0(n2113), .B1(n2203), .A0N(\register[20][27] ), .A1N(
        n2204), .Y(n743) );
  OAI2BB2XL U1111 ( .B0(n2111), .B1(n2202), .A0N(\register[20][28] ), .A1N(
        n2204), .Y(n744) );
  OAI2BB2XL U1112 ( .B0(n2109), .B1(n22), .A0N(\register[20][29] ), .A1N(n2204), .Y(n745) );
  OAI2BB2XL U1113 ( .B0(n2107), .B1(n22), .A0N(\register[20][30] ), .A1N(n2202), .Y(n746) );
  OAI2BB2XL U1114 ( .B0(n2105), .B1(n22), .A0N(\register[20][31] ), .A1N(n2203), .Y(n747) );
  OAI2BB2XL U1115 ( .B0(n2121), .B1(n2200), .A0N(\register[21][23] ), .A1N(
        n2201), .Y(n771) );
  OAI2BB2XL U1116 ( .B0(n2117), .B1(n23), .A0N(\register[21][25] ), .A1N(n2201), .Y(n773) );
  OAI2BB2XL U1117 ( .B0(n2115), .B1(n2199), .A0N(\register[21][26] ), .A1N(
        n2201), .Y(n774) );
  OAI2BB2XL U1118 ( .B0(n2113), .B1(n2200), .A0N(\register[21][27] ), .A1N(
        n2201), .Y(n775) );
  OAI2BB2XL U1119 ( .B0(n2111), .B1(n2199), .A0N(\register[21][28] ), .A1N(
        n2201), .Y(n776) );
  OAI2BB2XL U1120 ( .B0(n2109), .B1(n23), .A0N(\register[21][29] ), .A1N(n2201), .Y(n777) );
  OAI2BB2XL U1121 ( .B0(n2107), .B1(n23), .A0N(\register[21][30] ), .A1N(n2199), .Y(n778) );
  OAI2BB2XL U1122 ( .B0(n2105), .B1(n23), .A0N(\register[21][31] ), .A1N(n2200), .Y(n779) );
  OAI2BB2XL U1123 ( .B0(n2121), .B1(n2197), .A0N(\register[22][23] ), .A1N(
        n2198), .Y(n803) );
  OAI2BB2XL U1124 ( .B0(n2117), .B1(n24), .A0N(\register[22][25] ), .A1N(n2198), .Y(n805) );
  OAI2BB2XL U1125 ( .B0(n2115), .B1(n2196), .A0N(\register[22][26] ), .A1N(
        n2198), .Y(n806) );
  OAI2BB2XL U1126 ( .B0(n2113), .B1(n2197), .A0N(\register[22][27] ), .A1N(
        n2198), .Y(n807) );
  OAI2BB2XL U1127 ( .B0(n2111), .B1(n2196), .A0N(\register[22][28] ), .A1N(
        n2198), .Y(n808) );
  OAI2BB2XL U1128 ( .B0(n2109), .B1(n24), .A0N(\register[22][29] ), .A1N(n2198), .Y(n809) );
  OAI2BB2XL U1129 ( .B0(n2107), .B1(n24), .A0N(\register[22][30] ), .A1N(n2196), .Y(n810) );
  OAI2BB2XL U1130 ( .B0(n2105), .B1(n24), .A0N(\register[22][31] ), .A1N(n2197), .Y(n811) );
  OAI2BB2XL U1131 ( .B0(n2121), .B1(n2194), .A0N(\register[23][23] ), .A1N(
        n2195), .Y(n835) );
  OAI2BB2XL U1132 ( .B0(n2117), .B1(n25), .A0N(\register[23][25] ), .A1N(n2195), .Y(n837) );
  OAI2BB2XL U1133 ( .B0(n2115), .B1(n2193), .A0N(\register[23][26] ), .A1N(
        n2195), .Y(n838) );
  OAI2BB2XL U1134 ( .B0(n2113), .B1(n2194), .A0N(\register[23][27] ), .A1N(
        n2195), .Y(n839) );
  OAI2BB2XL U1135 ( .B0(n2111), .B1(n2193), .A0N(\register[23][28] ), .A1N(
        n2195), .Y(n840) );
  OAI2BB2XL U1136 ( .B0(n2109), .B1(n25), .A0N(\register[23][29] ), .A1N(n2195), .Y(n841) );
  OAI2BB2XL U1137 ( .B0(n2107), .B1(n25), .A0N(\register[23][30] ), .A1N(n2193), .Y(n842) );
  OAI2BB2XL U1138 ( .B0(n2105), .B1(n25), .A0N(\register[23][31] ), .A1N(n2194), .Y(n843) );
  OAI2BB2XL U1139 ( .B0(n2121), .B1(n2190), .A0N(\register[24][23] ), .A1N(
        n2190), .Y(n867) );
  OAI2BB2XL U1140 ( .B0(n2117), .B1(n2190), .A0N(\register[24][25] ), .A1N(
        n2192), .Y(n869) );
  OAI2BB2XL U1141 ( .B0(n2115), .B1(n2190), .A0N(\register[24][26] ), .A1N(
        n2192), .Y(n870) );
  OAI2BB2XL U1142 ( .B0(n2113), .B1(n2190), .A0N(\register[24][27] ), .A1N(
        n2192), .Y(n871) );
  OAI2BB2XL U1143 ( .B0(n2111), .B1(n2190), .A0N(\register[24][28] ), .A1N(
        n2192), .Y(n872) );
  OAI2BB2XL U1144 ( .B0(n2109), .B1(n2190), .A0N(\register[24][29] ), .A1N(
        n2192), .Y(n873) );
  OAI2BB2XL U1145 ( .B0(n2107), .B1(n2190), .A0N(\register[24][30] ), .A1N(
        n2191), .Y(n874) );
  OAI2BB2XL U1146 ( .B0(n2105), .B1(n2190), .A0N(\register[24][31] ), .A1N(
        n2191), .Y(n875) );
  OAI2BB2XL U1147 ( .B0(n2121), .B1(n2184), .A0N(\register[26][23] ), .A1N(
        n2184), .Y(n931) );
  OAI2BB2XL U1148 ( .B0(n2117), .B1(n2184), .A0N(\register[26][25] ), .A1N(
        n2186), .Y(n933) );
  OAI2BB2XL U1149 ( .B0(n2115), .B1(n2184), .A0N(\register[26][26] ), .A1N(
        n2186), .Y(n934) );
  OAI2BB2XL U1150 ( .B0(n2113), .B1(n2184), .A0N(\register[26][27] ), .A1N(
        n2186), .Y(n935) );
  OAI2BB2XL U1151 ( .B0(n2111), .B1(n2184), .A0N(\register[26][28] ), .A1N(
        n2186), .Y(n936) );
  OAI2BB2XL U1152 ( .B0(n2109), .B1(n2184), .A0N(\register[26][29] ), .A1N(
        n2186), .Y(n937) );
  OAI2BB2XL U1153 ( .B0(n2107), .B1(n2184), .A0N(\register[26][30] ), .A1N(
        n2185), .Y(n938) );
  OAI2BB2XL U1154 ( .B0(n2105), .B1(n2184), .A0N(\register[26][31] ), .A1N(
        n2185), .Y(n939) );
  OAI2BB2XL U1155 ( .B0(n2121), .B1(n2181), .A0N(\register[27][23] ), .A1N(
        n2181), .Y(n963) );
  OAI2BB2XL U1156 ( .B0(n2117), .B1(n2181), .A0N(\register[27][25] ), .A1N(
        n2183), .Y(n965) );
  OAI2BB2XL U1157 ( .B0(n2115), .B1(n2181), .A0N(\register[27][26] ), .A1N(
        n2183), .Y(n966) );
  OAI2BB2XL U1158 ( .B0(n2113), .B1(n2181), .A0N(\register[27][27] ), .A1N(
        n2183), .Y(n967) );
  OAI2BB2XL U1159 ( .B0(n2111), .B1(n2181), .A0N(\register[27][28] ), .A1N(
        n2183), .Y(n968) );
  OAI2BB2XL U1160 ( .B0(n2109), .B1(n2181), .A0N(\register[27][29] ), .A1N(
        n2183), .Y(n969) );
  OAI2BB2XL U1161 ( .B0(n2107), .B1(n2181), .A0N(\register[27][30] ), .A1N(
        n2182), .Y(n970) );
  OAI2BB2XL U1162 ( .B0(n2105), .B1(n2181), .A0N(\register[27][31] ), .A1N(
        n2182), .Y(n971) );
  OAI2BB2XL U1163 ( .B0(n2121), .B1(n2178), .A0N(\register[28][23] ), .A1N(
        n2178), .Y(n995) );
  OAI2BB2XL U1164 ( .B0(n2117), .B1(n2178), .A0N(\register[28][25] ), .A1N(
        n2180), .Y(n997) );
  OAI2BB2XL U1165 ( .B0(n2115), .B1(n2178), .A0N(\register[28][26] ), .A1N(
        n2180), .Y(n998) );
  OAI2BB2XL U1166 ( .B0(n2113), .B1(n2178), .A0N(\register[28][27] ), .A1N(
        n2180), .Y(n999) );
  OAI2BB2XL U1167 ( .B0(n2111), .B1(n2178), .A0N(\register[28][28] ), .A1N(
        n2180), .Y(n1000) );
  OAI2BB2XL U1168 ( .B0(n2109), .B1(n2178), .A0N(\register[28][29] ), .A1N(
        n2180), .Y(n1001) );
  OAI2BB2XL U1169 ( .B0(n2107), .B1(n2178), .A0N(\register[28][30] ), .A1N(
        n2179), .Y(n1002) );
  OAI2BB2XL U1170 ( .B0(n2105), .B1(n2178), .A0N(\register[28][31] ), .A1N(
        n2179), .Y(n1003) );
  OAI2BB2XL U1171 ( .B0(n2121), .B1(n2175), .A0N(\register[29][23] ), .A1N(
        n2175), .Y(n1027) );
  OAI2BB2XL U1172 ( .B0(n2117), .B1(n2175), .A0N(\register[29][25] ), .A1N(
        n2177), .Y(n1029) );
  OAI2BB2XL U1173 ( .B0(n2115), .B1(n2175), .A0N(\register[29][26] ), .A1N(
        n2177), .Y(n1030) );
  OAI2BB2XL U1174 ( .B0(n2113), .B1(n2175), .A0N(\register[29][27] ), .A1N(
        n2177), .Y(n1031) );
  OAI2BB2XL U1175 ( .B0(n2111), .B1(n2175), .A0N(\register[29][28] ), .A1N(
        n2177), .Y(n1032) );
  OAI2BB2XL U1176 ( .B0(n2109), .B1(n2175), .A0N(\register[29][29] ), .A1N(
        n2177), .Y(n1033) );
  OAI2BB2XL U1177 ( .B0(n2107), .B1(n2175), .A0N(\register[29][30] ), .A1N(
        n2176), .Y(n1034) );
  OAI2BB2XL U1178 ( .B0(n2105), .B1(n2175), .A0N(\register[29][31] ), .A1N(
        n2176), .Y(n1035) );
  OAI2BB2XL U1179 ( .B0(n2121), .B1(n2172), .A0N(\register[30][23] ), .A1N(
        n2172), .Y(n1059) );
  OAI2BB2XL U1180 ( .B0(n2117), .B1(n2172), .A0N(\register[30][25] ), .A1N(
        n2174), .Y(n1061) );
  OAI2BB2XL U1181 ( .B0(n2115), .B1(n2172), .A0N(\register[30][26] ), .A1N(
        n2174), .Y(n1062) );
  OAI2BB2XL U1182 ( .B0(n2113), .B1(n2172), .A0N(\register[30][27] ), .A1N(
        n2174), .Y(n1063) );
  OAI2BB2XL U1183 ( .B0(n2111), .B1(n2172), .A0N(\register[30][28] ), .A1N(
        n2174), .Y(n1064) );
  OAI2BB2XL U1184 ( .B0(n2109), .B1(n2172), .A0N(\register[30][29] ), .A1N(
        n2174), .Y(n1065) );
  OAI2BB2XL U1185 ( .B0(n2107), .B1(n2172), .A0N(\register[30][30] ), .A1N(
        n2173), .Y(n1066) );
  OAI2BB2XL U1186 ( .B0(n2105), .B1(n2172), .A0N(\register[30][31] ), .A1N(
        n2173), .Y(n1067) );
  OAI2BB2XL U1187 ( .B0(n2121), .B1(n2169), .A0N(\register[31][23] ), .A1N(
        n2169), .Y(n1091) );
  OAI2BB2XL U1188 ( .B0(n2117), .B1(n2169), .A0N(\register[31][25] ), .A1N(
        n2171), .Y(n1093) );
  OAI2BB2XL U1189 ( .B0(n2115), .B1(n2169), .A0N(\register[31][26] ), .A1N(
        n2171), .Y(n1094) );
  OAI2BB2XL U1190 ( .B0(n2113), .B1(n2169), .A0N(\register[31][27] ), .A1N(
        n2171), .Y(n1095) );
  OAI2BB2XL U1191 ( .B0(n2111), .B1(n2169), .A0N(\register[31][28] ), .A1N(
        n2171), .Y(n1096) );
  OAI2BB2XL U1192 ( .B0(n2109), .B1(n2169), .A0N(\register[31][29] ), .A1N(
        n2171), .Y(n1097) );
  OAI2BB2XL U1193 ( .B0(n2107), .B1(n2169), .A0N(\register[31][30] ), .A1N(
        n2170), .Y(n1098) );
  OAI2BB2XL U1194 ( .B0(n2105), .B1(n2169), .A0N(\register[31][31] ), .A1N(
        n2170), .Y(n1099) );
  OAI2BB2XL U1195 ( .B0(n2167), .B1(n2239), .A0N(\register[8][0] ), .A1N(n2239), .Y(n332) );
  OAI2BB2XL U1196 ( .B0(n2166), .B1(n2238), .A0N(\register[8][1] ), .A1N(n2238), .Y(n333) );
  OAI2BB2XL U1197 ( .B0(n2164), .B1(n2238), .A0N(\register[8][2] ), .A1N(n2239), .Y(n334) );
  OAI2BB2XL U1198 ( .B0(n2162), .B1(n2238), .A0N(\register[8][3] ), .A1N(n2240), .Y(n335) );
  OAI2BB2XL U1199 ( .B0(n2160), .B1(n2238), .A0N(\register[8][4] ), .A1N(n2238), .Y(n336) );
  OAI2BB2XL U1200 ( .B0(n2157), .B1(n2238), .A0N(\register[8][5] ), .A1N(n2240), .Y(n337) );
  OAI2BB2XL U1201 ( .B0(n2156), .B1(n2238), .A0N(\register[8][6] ), .A1N(n2240), .Y(n338) );
  OAI2BB2XL U1202 ( .B0(n2153), .B1(n2238), .A0N(\register[8][7] ), .A1N(n2240), .Y(n339) );
  OAI2BB2XL U1203 ( .B0(n2151), .B1(n2238), .A0N(\register[8][8] ), .A1N(n2240), .Y(n340) );
  OAI2BB2XL U1204 ( .B0(n2149), .B1(n2238), .A0N(\register[8][9] ), .A1N(n2240), .Y(n341) );
  OAI2BB2XL U1205 ( .B0(n2147), .B1(n2238), .A0N(\register[8][10] ), .A1N(
        n2240), .Y(n342) );
  OAI2BB2XL U1206 ( .B0(n2146), .B1(n2238), .A0N(\register[8][11] ), .A1N(
        n2240), .Y(n343) );
  OAI2BB2XL U1207 ( .B0(n2144), .B1(n2238), .A0N(\register[8][12] ), .A1N(
        n2240), .Y(n344) );
  OAI2BB2XL U1208 ( .B0(n2142), .B1(n2239), .A0N(\register[8][13] ), .A1N(
        n2240), .Y(n345) );
  OAI2BB2XL U1209 ( .B0(n2140), .B1(n2239), .A0N(\register[8][14] ), .A1N(
        n2240), .Y(n346) );
  OAI2BB2XL U1210 ( .B0(n2138), .B1(n2239), .A0N(\register[8][15] ), .A1N(
        n2240), .Y(n347) );
  OAI2BB2XL U1211 ( .B0(n2136), .B1(n2239), .A0N(\register[8][16] ), .A1N(
        n2240), .Y(n348) );
  OAI2BB2XL U1212 ( .B0(n2134), .B1(n2239), .A0N(\register[8][17] ), .A1N(
        n2240), .Y(n349) );
  OAI2BB2XL U1213 ( .B0(n2132), .B1(n2239), .A0N(\register[8][18] ), .A1N(
        n2239), .Y(n350) );
  OAI2BB2XL U1214 ( .B0(n2130), .B1(n2239), .A0N(\register[8][19] ), .A1N(
        n2238), .Y(n351) );
  OAI2BB2XL U1215 ( .B0(n2128), .B1(n2239), .A0N(\register[8][20] ), .A1N(
        n2240), .Y(n352) );
  OAI2BB2XL U1216 ( .B0(n2126), .B1(n2239), .A0N(\register[8][21] ), .A1N(
        n2239), .Y(n353) );
  OAI2BB2XL U1217 ( .B0(n2124), .B1(n2239), .A0N(\register[8][22] ), .A1N(
        n2240), .Y(n354) );
  OAI2BB2XL U1218 ( .B0(n2120), .B1(n2239), .A0N(\register[8][24] ), .A1N(
        n2240), .Y(n356) );
  OAI2BB2XL U1219 ( .B0(n2167), .B1(n2233), .A0N(\register[10][0] ), .A1N(
        n2233), .Y(n396) );
  OAI2BB2XL U1220 ( .B0(n2166), .B1(n2232), .A0N(\register[10][1] ), .A1N(
        n2232), .Y(n397) );
  OAI2BB2XL U1221 ( .B0(n2164), .B1(n2232), .A0N(\register[10][2] ), .A1N(
        n2233), .Y(n398) );
  OAI2BB2XL U1222 ( .B0(n2162), .B1(n2232), .A0N(\register[10][3] ), .A1N(
        n2234), .Y(n399) );
  OAI2BB2XL U1223 ( .B0(n2160), .B1(n2232), .A0N(\register[10][4] ), .A1N(
        n2232), .Y(n400) );
  OAI2BB2XL U1224 ( .B0(n2157), .B1(n2232), .A0N(\register[10][5] ), .A1N(
        n2234), .Y(n401) );
  OAI2BB2XL U1225 ( .B0(n2156), .B1(n2232), .A0N(\register[10][6] ), .A1N(
        n2234), .Y(n402) );
  OAI2BB2XL U1226 ( .B0(n2153), .B1(n2232), .A0N(\register[10][7] ), .A1N(
        n2234), .Y(n403) );
  OAI2BB2XL U1227 ( .B0(n2151), .B1(n2232), .A0N(\register[10][8] ), .A1N(
        n2234), .Y(n404) );
  OAI2BB2XL U1228 ( .B0(n2149), .B1(n2232), .A0N(\register[10][9] ), .A1N(
        n2234), .Y(n405) );
  OAI2BB2XL U1229 ( .B0(n2147), .B1(n2232), .A0N(\register[10][10] ), .A1N(
        n2234), .Y(n406) );
  OAI2BB2XL U1230 ( .B0(n2146), .B1(n2232), .A0N(\register[10][11] ), .A1N(
        n2234), .Y(n407) );
  OAI2BB2XL U1231 ( .B0(n2144), .B1(n2232), .A0N(\register[10][12] ), .A1N(
        n2234), .Y(n408) );
  OAI2BB2XL U1232 ( .B0(n2142), .B1(n2233), .A0N(\register[10][13] ), .A1N(
        n2234), .Y(n409) );
  OAI2BB2XL U1233 ( .B0(n2140), .B1(n2233), .A0N(\register[10][14] ), .A1N(
        n2234), .Y(n410) );
  OAI2BB2XL U1234 ( .B0(n2138), .B1(n2233), .A0N(\register[10][15] ), .A1N(
        n2234), .Y(n411) );
  OAI2BB2XL U1235 ( .B0(n2136), .B1(n2233), .A0N(\register[10][16] ), .A1N(
        n2234), .Y(n412) );
  OAI2BB2XL U1236 ( .B0(n2134), .B1(n2233), .A0N(\register[10][17] ), .A1N(
        n2234), .Y(n413) );
  OAI2BB2XL U1237 ( .B0(n2132), .B1(n2233), .A0N(\register[10][18] ), .A1N(
        n2233), .Y(n414) );
  OAI2BB2XL U1238 ( .B0(n2130), .B1(n2233), .A0N(\register[10][19] ), .A1N(
        n2232), .Y(n415) );
  OAI2BB2XL U1239 ( .B0(n2128), .B1(n2233), .A0N(\register[10][20] ), .A1N(
        n2234), .Y(n416) );
  OAI2BB2XL U1240 ( .B0(n2126), .B1(n2233), .A0N(\register[10][21] ), .A1N(
        n2233), .Y(n417) );
  OAI2BB2XL U1241 ( .B0(n2124), .B1(n2233), .A0N(\register[10][22] ), .A1N(
        n2234), .Y(n418) );
  OAI2BB2XL U1242 ( .B0(n2120), .B1(n2233), .A0N(\register[10][24] ), .A1N(
        n2234), .Y(n420) );
  OAI2BB2XL U1243 ( .B0(n2167), .B1(n2230), .A0N(\register[11][0] ), .A1N(
        n2230), .Y(n428) );
  OAI2BB2XL U1244 ( .B0(n2166), .B1(n2229), .A0N(\register[11][1] ), .A1N(
        n2229), .Y(n429) );
  OAI2BB2XL U1245 ( .B0(n2164), .B1(n2229), .A0N(\register[11][2] ), .A1N(
        n2230), .Y(n430) );
  OAI2BB2XL U1246 ( .B0(n2162), .B1(n2229), .A0N(\register[11][3] ), .A1N(
        n2231), .Y(n431) );
  OAI2BB2XL U1247 ( .B0(n2160), .B1(n2229), .A0N(\register[11][4] ), .A1N(
        n2229), .Y(n432) );
  OAI2BB2XL U1248 ( .B0(n2157), .B1(n2229), .A0N(\register[11][5] ), .A1N(
        n2231), .Y(n433) );
  OAI2BB2XL U1249 ( .B0(n2156), .B1(n2229), .A0N(\register[11][6] ), .A1N(
        n2231), .Y(n434) );
  OAI2BB2XL U1250 ( .B0(n2153), .B1(n2229), .A0N(\register[11][7] ), .A1N(
        n2231), .Y(n435) );
  OAI2BB2XL U1251 ( .B0(n2151), .B1(n2229), .A0N(\register[11][8] ), .A1N(
        n2231), .Y(n436) );
  OAI2BB2XL U1252 ( .B0(n2149), .B1(n2229), .A0N(\register[11][9] ), .A1N(
        n2231), .Y(n437) );
  OAI2BB2XL U1253 ( .B0(n2147), .B1(n2229), .A0N(\register[11][10] ), .A1N(
        n2231), .Y(n438) );
  OAI2BB2XL U1254 ( .B0(n2146), .B1(n2229), .A0N(\register[11][11] ), .A1N(
        n2231), .Y(n439) );
  OAI2BB2XL U1255 ( .B0(n2144), .B1(n2229), .A0N(\register[11][12] ), .A1N(
        n2231), .Y(n440) );
  OAI2BB2XL U1256 ( .B0(n2142), .B1(n2230), .A0N(\register[11][13] ), .A1N(
        n2231), .Y(n441) );
  OAI2BB2XL U1257 ( .B0(n2140), .B1(n2230), .A0N(\register[11][14] ), .A1N(
        n2231), .Y(n442) );
  OAI2BB2XL U1258 ( .B0(n2138), .B1(n2230), .A0N(\register[11][15] ), .A1N(
        n2231), .Y(n443) );
  OAI2BB2XL U1259 ( .B0(n2136), .B1(n2230), .A0N(\register[11][16] ), .A1N(
        n2231), .Y(n444) );
  OAI2BB2XL U1260 ( .B0(n2134), .B1(n2230), .A0N(\register[11][17] ), .A1N(
        n2231), .Y(n445) );
  OAI2BB2XL U1261 ( .B0(n2132), .B1(n2230), .A0N(\register[11][18] ), .A1N(
        n2230), .Y(n446) );
  OAI2BB2XL U1262 ( .B0(n2130), .B1(n2230), .A0N(\register[11][19] ), .A1N(
        n2229), .Y(n447) );
  OAI2BB2XL U1263 ( .B0(n2128), .B1(n2230), .A0N(\register[11][20] ), .A1N(
        n2231), .Y(n448) );
  OAI2BB2XL U1264 ( .B0(n2126), .B1(n2230), .A0N(\register[11][21] ), .A1N(
        n2230), .Y(n449) );
  OAI2BB2XL U1265 ( .B0(n2124), .B1(n2230), .A0N(\register[11][22] ), .A1N(
        n2231), .Y(n450) );
  OAI2BB2XL U1266 ( .B0(n2120), .B1(n2230), .A0N(\register[11][24] ), .A1N(
        n2231), .Y(n452) );
  OAI2BB2XL U1267 ( .B0(n2167), .B1(n2227), .A0N(\register[12][0] ), .A1N(
        n2227), .Y(n460) );
  OAI2BB2XL U1268 ( .B0(n2166), .B1(n2226), .A0N(\register[12][1] ), .A1N(
        n2226), .Y(n461) );
  OAI2BB2XL U1269 ( .B0(n2164), .B1(n2226), .A0N(\register[12][2] ), .A1N(
        n2227), .Y(n462) );
  OAI2BB2XL U1270 ( .B0(n2162), .B1(n2226), .A0N(\register[12][3] ), .A1N(
        n2228), .Y(n463) );
  OAI2BB2XL U1271 ( .B0(n2160), .B1(n2226), .A0N(\register[12][4] ), .A1N(
        n2226), .Y(n464) );
  OAI2BB2XL U1272 ( .B0(n2157), .B1(n2226), .A0N(\register[12][5] ), .A1N(
        n2228), .Y(n465) );
  OAI2BB2XL U1273 ( .B0(n2156), .B1(n2226), .A0N(\register[12][6] ), .A1N(
        n2228), .Y(n466) );
  OAI2BB2XL U1274 ( .B0(n2153), .B1(n2226), .A0N(\register[12][7] ), .A1N(
        n2228), .Y(n467) );
  OAI2BB2XL U1275 ( .B0(n2151), .B1(n2226), .A0N(\register[12][8] ), .A1N(
        n2228), .Y(n468) );
  OAI2BB2XL U1276 ( .B0(n2149), .B1(n2226), .A0N(\register[12][9] ), .A1N(
        n2228), .Y(n469) );
  OAI2BB2XL U1277 ( .B0(n2147), .B1(n2226), .A0N(\register[12][10] ), .A1N(
        n2228), .Y(n470) );
  OAI2BB2XL U1278 ( .B0(n2146), .B1(n2226), .A0N(\register[12][11] ), .A1N(
        n2228), .Y(n471) );
  OAI2BB2XL U1279 ( .B0(n2144), .B1(n2226), .A0N(\register[12][12] ), .A1N(
        n2228), .Y(n472) );
  OAI2BB2XL U1280 ( .B0(n2142), .B1(n2227), .A0N(\register[12][13] ), .A1N(
        n2228), .Y(n473) );
  OAI2BB2XL U1281 ( .B0(n2140), .B1(n2227), .A0N(\register[12][14] ), .A1N(
        n2228), .Y(n474) );
  OAI2BB2XL U1282 ( .B0(n2138), .B1(n2227), .A0N(\register[12][15] ), .A1N(
        n2228), .Y(n475) );
  OAI2BB2XL U1283 ( .B0(n2136), .B1(n2227), .A0N(\register[12][16] ), .A1N(
        n2228), .Y(n476) );
  OAI2BB2XL U1284 ( .B0(n2134), .B1(n2227), .A0N(\register[12][17] ), .A1N(
        n2228), .Y(n477) );
  OAI2BB2XL U1285 ( .B0(n2132), .B1(n2227), .A0N(\register[12][18] ), .A1N(
        n2227), .Y(n478) );
  OAI2BB2XL U1286 ( .B0(n2130), .B1(n2227), .A0N(\register[12][19] ), .A1N(
        n2226), .Y(n479) );
  OAI2BB2XL U1287 ( .B0(n2128), .B1(n2227), .A0N(\register[12][20] ), .A1N(
        n2228), .Y(n480) );
  OAI2BB2XL U1288 ( .B0(n2126), .B1(n2227), .A0N(\register[12][21] ), .A1N(
        n2227), .Y(n481) );
  OAI2BB2XL U1289 ( .B0(n2124), .B1(n2227), .A0N(\register[12][22] ), .A1N(
        n2228), .Y(n482) );
  OAI2BB2XL U1290 ( .B0(n2120), .B1(n2227), .A0N(\register[12][24] ), .A1N(
        n2228), .Y(n484) );
  OAI2BB2XL U1291 ( .B0(n2167), .B1(n2224), .A0N(\register[13][0] ), .A1N(
        n2224), .Y(n492) );
  OAI2BB2XL U1292 ( .B0(n2166), .B1(n2223), .A0N(\register[13][1] ), .A1N(
        n2223), .Y(n493) );
  OAI2BB2XL U1293 ( .B0(n2164), .B1(n2223), .A0N(\register[13][2] ), .A1N(
        n2224), .Y(n494) );
  OAI2BB2XL U1294 ( .B0(n2162), .B1(n2223), .A0N(\register[13][3] ), .A1N(
        n2225), .Y(n495) );
  OAI2BB2XL U1295 ( .B0(n2160), .B1(n2223), .A0N(\register[13][4] ), .A1N(
        n2223), .Y(n496) );
  OAI2BB2XL U1296 ( .B0(n2157), .B1(n2223), .A0N(\register[13][5] ), .A1N(
        n2225), .Y(n497) );
  OAI2BB2XL U1297 ( .B0(n2156), .B1(n2223), .A0N(\register[13][6] ), .A1N(
        n2225), .Y(n498) );
  OAI2BB2XL U1298 ( .B0(n2153), .B1(n2223), .A0N(\register[13][7] ), .A1N(
        n2225), .Y(n499) );
  OAI2BB2XL U1299 ( .B0(n2151), .B1(n2223), .A0N(\register[13][8] ), .A1N(
        n2225), .Y(n500) );
  OAI2BB2XL U1300 ( .B0(n2149), .B1(n2223), .A0N(\register[13][9] ), .A1N(
        n2225), .Y(n501) );
  OAI2BB2XL U1301 ( .B0(n2147), .B1(n2223), .A0N(\register[13][10] ), .A1N(
        n2225), .Y(n502) );
  OAI2BB2XL U1302 ( .B0(n2146), .B1(n2223), .A0N(\register[13][11] ), .A1N(
        n2225), .Y(n503) );
  OAI2BB2XL U1303 ( .B0(n2144), .B1(n2223), .A0N(\register[13][12] ), .A1N(
        n2225), .Y(n504) );
  OAI2BB2XL U1304 ( .B0(n2142), .B1(n2224), .A0N(\register[13][13] ), .A1N(
        n2225), .Y(n505) );
  OAI2BB2XL U1305 ( .B0(n2140), .B1(n2224), .A0N(\register[13][14] ), .A1N(
        n2225), .Y(n506) );
  OAI2BB2XL U1306 ( .B0(n2138), .B1(n2224), .A0N(\register[13][15] ), .A1N(
        n2225), .Y(n507) );
  OAI2BB2XL U1307 ( .B0(n2136), .B1(n2224), .A0N(\register[13][16] ), .A1N(
        n2225), .Y(n508) );
  OAI2BB2XL U1308 ( .B0(n2134), .B1(n2224), .A0N(\register[13][17] ), .A1N(
        n2225), .Y(n509) );
  OAI2BB2XL U1309 ( .B0(n2132), .B1(n2224), .A0N(\register[13][18] ), .A1N(
        n2224), .Y(n510) );
  OAI2BB2XL U1310 ( .B0(n2130), .B1(n2224), .A0N(\register[13][19] ), .A1N(
        n2223), .Y(n511) );
  OAI2BB2XL U1311 ( .B0(n2128), .B1(n2224), .A0N(\register[13][20] ), .A1N(
        n2225), .Y(n512) );
  OAI2BB2XL U1312 ( .B0(n2126), .B1(n2224), .A0N(\register[13][21] ), .A1N(
        n2224), .Y(n513) );
  OAI2BB2XL U1313 ( .B0(n2124), .B1(n2224), .A0N(\register[13][22] ), .A1N(
        n2225), .Y(n514) );
  OAI2BB2XL U1314 ( .B0(n2120), .B1(n2224), .A0N(\register[13][24] ), .A1N(
        n2225), .Y(n516) );
  OAI2BB2XL U1315 ( .B0(n2167), .B1(n2221), .A0N(\register[14][0] ), .A1N(
        n2221), .Y(n524) );
  OAI2BB2XL U1316 ( .B0(n2166), .B1(n2220), .A0N(\register[14][1] ), .A1N(
        n2220), .Y(n525) );
  OAI2BB2XL U1317 ( .B0(n2164), .B1(n2220), .A0N(\register[14][2] ), .A1N(
        n2221), .Y(n526) );
  OAI2BB2XL U1318 ( .B0(n2162), .B1(n2220), .A0N(\register[14][3] ), .A1N(
        n2222), .Y(n527) );
  OAI2BB2XL U1319 ( .B0(n2160), .B1(n2220), .A0N(\register[14][4] ), .A1N(
        n2220), .Y(n528) );
  OAI2BB2XL U1320 ( .B0(n2157), .B1(n2220), .A0N(\register[14][5] ), .A1N(
        n2222), .Y(n529) );
  OAI2BB2XL U1321 ( .B0(n2156), .B1(n2220), .A0N(\register[14][6] ), .A1N(
        n2222), .Y(n530) );
  OAI2BB2XL U1322 ( .B0(n2153), .B1(n2220), .A0N(\register[14][7] ), .A1N(
        n2222), .Y(n531) );
  OAI2BB2XL U1323 ( .B0(n2151), .B1(n2220), .A0N(\register[14][8] ), .A1N(
        n2222), .Y(n532) );
  OAI2BB2XL U1324 ( .B0(n2149), .B1(n2220), .A0N(\register[14][9] ), .A1N(
        n2222), .Y(n533) );
  OAI2BB2XL U1325 ( .B0(n2147), .B1(n2220), .A0N(\register[14][10] ), .A1N(
        n2222), .Y(n534) );
  OAI2BB2XL U1326 ( .B0(n2146), .B1(n2220), .A0N(\register[14][11] ), .A1N(
        n2222), .Y(n535) );
  OAI2BB2XL U1327 ( .B0(n2144), .B1(n2220), .A0N(\register[14][12] ), .A1N(
        n2222), .Y(n536) );
  OAI2BB2XL U1328 ( .B0(n2142), .B1(n2221), .A0N(\register[14][13] ), .A1N(
        n2222), .Y(n537) );
  OAI2BB2XL U1329 ( .B0(n2140), .B1(n2221), .A0N(\register[14][14] ), .A1N(
        n2222), .Y(n538) );
  OAI2BB2XL U1330 ( .B0(n2138), .B1(n2221), .A0N(\register[14][15] ), .A1N(
        n2222), .Y(n539) );
  OAI2BB2XL U1331 ( .B0(n2136), .B1(n2221), .A0N(\register[14][16] ), .A1N(
        n2222), .Y(n540) );
  OAI2BB2XL U1332 ( .B0(n2134), .B1(n2221), .A0N(\register[14][17] ), .A1N(
        n2222), .Y(n541) );
  OAI2BB2XL U1333 ( .B0(n2132), .B1(n2221), .A0N(\register[14][18] ), .A1N(
        n2221), .Y(n542) );
  OAI2BB2XL U1334 ( .B0(n2130), .B1(n2221), .A0N(\register[14][19] ), .A1N(
        n2220), .Y(n543) );
  OAI2BB2XL U1335 ( .B0(n2128), .B1(n2221), .A0N(\register[14][20] ), .A1N(
        n2222), .Y(n544) );
  OAI2BB2XL U1336 ( .B0(n2126), .B1(n2221), .A0N(\register[14][21] ), .A1N(
        n2221), .Y(n545) );
  OAI2BB2XL U1337 ( .B0(n2124), .B1(n2221), .A0N(\register[14][22] ), .A1N(
        n2222), .Y(n546) );
  OAI2BB2XL U1338 ( .B0(n2120), .B1(n2221), .A0N(\register[14][24] ), .A1N(
        n2222), .Y(n548) );
  OAI2BB2XL U1339 ( .B0(n2167), .B1(n2218), .A0N(\register[15][0] ), .A1N(
        n2218), .Y(n556) );
  OAI2BB2XL U1340 ( .B0(n2166), .B1(n2217), .A0N(\register[15][1] ), .A1N(
        n2217), .Y(n557) );
  OAI2BB2XL U1341 ( .B0(n2164), .B1(n2217), .A0N(\register[15][2] ), .A1N(
        n2218), .Y(n558) );
  OAI2BB2XL U1342 ( .B0(n2162), .B1(n2217), .A0N(\register[15][3] ), .A1N(
        n2219), .Y(n559) );
  OAI2BB2XL U1343 ( .B0(n2160), .B1(n2217), .A0N(\register[15][4] ), .A1N(
        n2217), .Y(n560) );
  OAI2BB2XL U1344 ( .B0(n2157), .B1(n2217), .A0N(\register[15][5] ), .A1N(
        n2219), .Y(n561) );
  OAI2BB2XL U1345 ( .B0(n2156), .B1(n2217), .A0N(\register[15][6] ), .A1N(
        n2219), .Y(n562) );
  OAI2BB2XL U1346 ( .B0(n2153), .B1(n2217), .A0N(\register[15][7] ), .A1N(
        n2219), .Y(n563) );
  OAI2BB2XL U1347 ( .B0(n2151), .B1(n2217), .A0N(\register[15][8] ), .A1N(
        n2219), .Y(n564) );
  OAI2BB2XL U1348 ( .B0(n2149), .B1(n2217), .A0N(\register[15][9] ), .A1N(
        n2219), .Y(n565) );
  OAI2BB2XL U1349 ( .B0(n2147), .B1(n2217), .A0N(\register[15][10] ), .A1N(
        n2219), .Y(n566) );
  OAI2BB2XL U1350 ( .B0(n2146), .B1(n2217), .A0N(\register[15][11] ), .A1N(
        n2219), .Y(n567) );
  OAI2BB2XL U1351 ( .B0(n2144), .B1(n2217), .A0N(\register[15][12] ), .A1N(
        n2219), .Y(n568) );
  OAI2BB2XL U1352 ( .B0(n2142), .B1(n2218), .A0N(\register[15][13] ), .A1N(
        n2219), .Y(n569) );
  OAI2BB2XL U1353 ( .B0(n2140), .B1(n2218), .A0N(\register[15][14] ), .A1N(
        n2219), .Y(n570) );
  OAI2BB2XL U1354 ( .B0(n2138), .B1(n2218), .A0N(\register[15][15] ), .A1N(
        n2219), .Y(n571) );
  OAI2BB2XL U1355 ( .B0(n2136), .B1(n2218), .A0N(\register[15][16] ), .A1N(
        n2219), .Y(n572) );
  OAI2BB2XL U1356 ( .B0(n2134), .B1(n2218), .A0N(\register[15][17] ), .A1N(
        n2219), .Y(n573) );
  OAI2BB2XL U1357 ( .B0(n2132), .B1(n2218), .A0N(\register[15][18] ), .A1N(
        n2218), .Y(n574) );
  OAI2BB2XL U1358 ( .B0(n2130), .B1(n2218), .A0N(\register[15][19] ), .A1N(
        n2217), .Y(n575) );
  OAI2BB2XL U1359 ( .B0(n2128), .B1(n2218), .A0N(\register[15][20] ), .A1N(
        n2219), .Y(n576) );
  OAI2BB2XL U1360 ( .B0(n2126), .B1(n2218), .A0N(\register[15][21] ), .A1N(
        n2218), .Y(n577) );
  OAI2BB2XL U1361 ( .B0(n2124), .B1(n2218), .A0N(\register[15][22] ), .A1N(
        n2219), .Y(n578) );
  OAI2BB2XL U1362 ( .B0(n2120), .B1(n2218), .A0N(\register[15][24] ), .A1N(
        n2219), .Y(n580) );
  OAI2BB2XL U1363 ( .B0(n2167), .B1(n2215), .A0N(\register[16][0] ), .A1N(
        n2215), .Y(n588) );
  OAI2BB2XL U1364 ( .B0(n2166), .B1(n2214), .A0N(\register[16][1] ), .A1N(
        n2214), .Y(n589) );
  OAI2BB2XL U1365 ( .B0(n2164), .B1(n2214), .A0N(\register[16][2] ), .A1N(
        n2215), .Y(n590) );
  OAI2BB2XL U1366 ( .B0(n2162), .B1(n2214), .A0N(\register[16][3] ), .A1N(
        n2216), .Y(n591) );
  OAI2BB2XL U1367 ( .B0(n2160), .B1(n2214), .A0N(\register[16][4] ), .A1N(
        n2214), .Y(n592) );
  OAI2BB2XL U1368 ( .B0(n2157), .B1(n2214), .A0N(\register[16][5] ), .A1N(
        n2216), .Y(n593) );
  OAI2BB2XL U1369 ( .B0(n2156), .B1(n2214), .A0N(\register[16][6] ), .A1N(
        n2216), .Y(n594) );
  OAI2BB2XL U1370 ( .B0(n2153), .B1(n2214), .A0N(\register[16][7] ), .A1N(
        n2216), .Y(n595) );
  OAI2BB2XL U1371 ( .B0(n2151), .B1(n2214), .A0N(\register[16][8] ), .A1N(
        n2216), .Y(n596) );
  OAI2BB2XL U1372 ( .B0(n2149), .B1(n2214), .A0N(\register[16][9] ), .A1N(
        n2216), .Y(n597) );
  OAI2BB2XL U1373 ( .B0(n2147), .B1(n2214), .A0N(\register[16][10] ), .A1N(
        n2216), .Y(n598) );
  OAI2BB2XL U1374 ( .B0(n2146), .B1(n2214), .A0N(\register[16][11] ), .A1N(
        n2216), .Y(n599) );
  OAI2BB2XL U1375 ( .B0(n2144), .B1(n2214), .A0N(\register[16][12] ), .A1N(
        n2216), .Y(n600) );
  OAI2BB2XL U1376 ( .B0(n2142), .B1(n2215), .A0N(\register[16][13] ), .A1N(
        n2216), .Y(n601) );
  OAI2BB2XL U1377 ( .B0(n2140), .B1(n2215), .A0N(\register[16][14] ), .A1N(
        n2216), .Y(n602) );
  OAI2BB2XL U1378 ( .B0(n2138), .B1(n2215), .A0N(\register[16][15] ), .A1N(
        n2216), .Y(n603) );
  OAI2BB2XL U1379 ( .B0(n2136), .B1(n2215), .A0N(\register[16][16] ), .A1N(
        n2216), .Y(n604) );
  OAI2BB2XL U1380 ( .B0(n2134), .B1(n2215), .A0N(\register[16][17] ), .A1N(
        n2216), .Y(n605) );
  OAI2BB2XL U1381 ( .B0(n2132), .B1(n2215), .A0N(\register[16][18] ), .A1N(
        n2215), .Y(n606) );
  OAI2BB2XL U1382 ( .B0(n2130), .B1(n2215), .A0N(\register[16][19] ), .A1N(
        n2214), .Y(n607) );
  OAI2BB2XL U1383 ( .B0(n2128), .B1(n2215), .A0N(\register[16][20] ), .A1N(
        n2216), .Y(n608) );
  OAI2BB2XL U1384 ( .B0(n2126), .B1(n2215), .A0N(\register[16][21] ), .A1N(
        n2215), .Y(n609) );
  OAI2BB2XL U1385 ( .B0(n2124), .B1(n2215), .A0N(\register[16][22] ), .A1N(
        n2216), .Y(n610) );
  OAI2BB2XL U1386 ( .B0(n2120), .B1(n2215), .A0N(\register[16][24] ), .A1N(
        n2216), .Y(n612) );
  OAI2BB2XL U1387 ( .B0(n2167), .B1(n2209), .A0N(\register[18][0] ), .A1N(
        n2209), .Y(n652) );
  OAI2BB2XL U1388 ( .B0(n2166), .B1(n2208), .A0N(\register[18][1] ), .A1N(
        n2208), .Y(n653) );
  OAI2BB2XL U1389 ( .B0(n2164), .B1(n2208), .A0N(\register[18][2] ), .A1N(
        n2209), .Y(n654) );
  OAI2BB2XL U1390 ( .B0(n2162), .B1(n2208), .A0N(\register[18][3] ), .A1N(
        n2210), .Y(n655) );
  OAI2BB2XL U1391 ( .B0(n2160), .B1(n2208), .A0N(\register[18][4] ), .A1N(
        n2208), .Y(n656) );
  OAI2BB2XL U1392 ( .B0(n2157), .B1(n2208), .A0N(\register[18][5] ), .A1N(
        n2210), .Y(n657) );
  OAI2BB2XL U1393 ( .B0(n2156), .B1(n2208), .A0N(\register[18][6] ), .A1N(
        n2210), .Y(n658) );
  OAI2BB2XL U1394 ( .B0(n2153), .B1(n2208), .A0N(\register[18][7] ), .A1N(
        n2210), .Y(n659) );
  OAI2BB2XL U1395 ( .B0(n2151), .B1(n2208), .A0N(\register[18][8] ), .A1N(
        n2210), .Y(n660) );
  OAI2BB2XL U1396 ( .B0(n2149), .B1(n2208), .A0N(\register[18][9] ), .A1N(
        n2210), .Y(n661) );
  OAI2BB2XL U1397 ( .B0(n2147), .B1(n2208), .A0N(\register[18][10] ), .A1N(
        n2210), .Y(n662) );
  OAI2BB2XL U1398 ( .B0(n2146), .B1(n2208), .A0N(\register[18][11] ), .A1N(
        n2210), .Y(n663) );
  OAI2BB2XL U1399 ( .B0(n2144), .B1(n2208), .A0N(\register[18][12] ), .A1N(
        n2210), .Y(n664) );
  OAI2BB2XL U1400 ( .B0(n2142), .B1(n2209), .A0N(\register[18][13] ), .A1N(
        n2210), .Y(n665) );
  OAI2BB2XL U1401 ( .B0(n2140), .B1(n2209), .A0N(\register[18][14] ), .A1N(
        n2210), .Y(n666) );
  OAI2BB2XL U1402 ( .B0(n2138), .B1(n2209), .A0N(\register[18][15] ), .A1N(
        n2210), .Y(n667) );
  OAI2BB2XL U1403 ( .B0(n2136), .B1(n2209), .A0N(\register[18][16] ), .A1N(
        n2210), .Y(n668) );
  OAI2BB2XL U1404 ( .B0(n2134), .B1(n2209), .A0N(\register[18][17] ), .A1N(
        n2210), .Y(n669) );
  OAI2BB2XL U1405 ( .B0(n2132), .B1(n2209), .A0N(\register[18][18] ), .A1N(
        n2209), .Y(n670) );
  OAI2BB2XL U1406 ( .B0(n2130), .B1(n2209), .A0N(\register[18][19] ), .A1N(
        n2208), .Y(n671) );
  OAI2BB2XL U1407 ( .B0(n2128), .B1(n2209), .A0N(\register[18][20] ), .A1N(
        n2210), .Y(n672) );
  OAI2BB2XL U1408 ( .B0(n2126), .B1(n2209), .A0N(\register[18][21] ), .A1N(
        n2209), .Y(n673) );
  OAI2BB2XL U1409 ( .B0(n2124), .B1(n2209), .A0N(\register[18][22] ), .A1N(
        n2210), .Y(n674) );
  OAI2BB2XL U1410 ( .B0(n2120), .B1(n2209), .A0N(\register[18][24] ), .A1N(
        n2210), .Y(n676) );
  OAI2BB2XL U1411 ( .B0(n2167), .B1(n2206), .A0N(\register[19][0] ), .A1N(
        n2206), .Y(n684) );
  OAI2BB2XL U1412 ( .B0(n2166), .B1(n2205), .A0N(\register[19][1] ), .A1N(
        n2205), .Y(n685) );
  OAI2BB2XL U1413 ( .B0(n2164), .B1(n2205), .A0N(\register[19][2] ), .A1N(
        n2206), .Y(n686) );
  OAI2BB2XL U1414 ( .B0(n2162), .B1(n2205), .A0N(\register[19][3] ), .A1N(
        n2207), .Y(n687) );
  OAI2BB2XL U1415 ( .B0(n2160), .B1(n2205), .A0N(\register[19][4] ), .A1N(
        n2205), .Y(n688) );
  OAI2BB2XL U1416 ( .B0(n2157), .B1(n2205), .A0N(\register[19][5] ), .A1N(
        n2207), .Y(n689) );
  OAI2BB2XL U1417 ( .B0(n2156), .B1(n2205), .A0N(\register[19][6] ), .A1N(
        n2207), .Y(n690) );
  OAI2BB2XL U1418 ( .B0(n2153), .B1(n2205), .A0N(\register[19][7] ), .A1N(
        n2207), .Y(n691) );
  OAI2BB2XL U1419 ( .B0(n2151), .B1(n2205), .A0N(\register[19][8] ), .A1N(
        n2207), .Y(n692) );
  OAI2BB2XL U1420 ( .B0(n2149), .B1(n2205), .A0N(\register[19][9] ), .A1N(
        n2207), .Y(n693) );
  OAI2BB2XL U1421 ( .B0(n2147), .B1(n2205), .A0N(\register[19][10] ), .A1N(
        n2207), .Y(n694) );
  OAI2BB2XL U1422 ( .B0(n2146), .B1(n2205), .A0N(\register[19][11] ), .A1N(
        n2207), .Y(n695) );
  OAI2BB2XL U1423 ( .B0(n2144), .B1(n2205), .A0N(\register[19][12] ), .A1N(
        n2207), .Y(n696) );
  OAI2BB2XL U1424 ( .B0(n2142), .B1(n2206), .A0N(\register[19][13] ), .A1N(
        n2207), .Y(n697) );
  OAI2BB2XL U1425 ( .B0(n2140), .B1(n2206), .A0N(\register[19][14] ), .A1N(
        n2207), .Y(n698) );
  OAI2BB2XL U1426 ( .B0(n2138), .B1(n2206), .A0N(\register[19][15] ), .A1N(
        n2207), .Y(n699) );
  OAI2BB2XL U1427 ( .B0(n2136), .B1(n2206), .A0N(\register[19][16] ), .A1N(
        n2207), .Y(n700) );
  OAI2BB2XL U1428 ( .B0(n2134), .B1(n2206), .A0N(\register[19][17] ), .A1N(
        n2207), .Y(n701) );
  OAI2BB2XL U1429 ( .B0(n2132), .B1(n2206), .A0N(\register[19][18] ), .A1N(
        n2206), .Y(n702) );
  OAI2BB2XL U1430 ( .B0(n2130), .B1(n2206), .A0N(\register[19][19] ), .A1N(
        n2205), .Y(n703) );
  OAI2BB2XL U1431 ( .B0(n2128), .B1(n2206), .A0N(\register[19][20] ), .A1N(
        n2207), .Y(n704) );
  OAI2BB2XL U1432 ( .B0(n2126), .B1(n2206), .A0N(\register[19][21] ), .A1N(
        n2206), .Y(n705) );
  OAI2BB2XL U1433 ( .B0(n2124), .B1(n2206), .A0N(\register[19][22] ), .A1N(
        n2207), .Y(n706) );
  OAI2BB2XL U1434 ( .B0(n2120), .B1(n2206), .A0N(\register[19][24] ), .A1N(
        n2207), .Y(n708) );
  OAI2BB2XL U1435 ( .B0(n2167), .B1(n2203), .A0N(\register[20][0] ), .A1N(
        n2203), .Y(n716) );
  OAI2BB2XL U1436 ( .B0(n2165), .B1(n2202), .A0N(\register[20][1] ), .A1N(
        n2202), .Y(n717) );
  OAI2BB2XL U1437 ( .B0(n2163), .B1(n2202), .A0N(\register[20][2] ), .A1N(
        n2203), .Y(n718) );
  OAI2BB2XL U1438 ( .B0(n2161), .B1(n2202), .A0N(\register[20][3] ), .A1N(
        n2204), .Y(n719) );
  OAI2BB2XL U1439 ( .B0(n2159), .B1(n2202), .A0N(\register[20][4] ), .A1N(
        n2202), .Y(n720) );
  OAI2BB2XL U1440 ( .B0(n2157), .B1(n2202), .A0N(\register[20][5] ), .A1N(
        n2204), .Y(n721) );
  OAI2BB2XL U1441 ( .B0(n2155), .B1(n2202), .A0N(\register[20][6] ), .A1N(
        n2204), .Y(n722) );
  OAI2BB2XL U1442 ( .B0(n2153), .B1(n2202), .A0N(\register[20][7] ), .A1N(
        n2204), .Y(n723) );
  OAI2BB2XL U1443 ( .B0(n2151), .B1(n2202), .A0N(\register[20][8] ), .A1N(
        n2204), .Y(n724) );
  OAI2BB2XL U1444 ( .B0(n2149), .B1(n2202), .A0N(\register[20][9] ), .A1N(
        n2204), .Y(n725) );
  OAI2BB2XL U1445 ( .B0(n2147), .B1(n2202), .A0N(\register[20][10] ), .A1N(
        n2204), .Y(n726) );
  OAI2BB2XL U1446 ( .B0(n2145), .B1(n2202), .A0N(\register[20][11] ), .A1N(
        n2204), .Y(n727) );
  OAI2BB2XL U1447 ( .B0(n2143), .B1(n2202), .A0N(\register[20][12] ), .A1N(
        n2204), .Y(n728) );
  OAI2BB2XL U1448 ( .B0(n2141), .B1(n2203), .A0N(\register[20][13] ), .A1N(
        n2204), .Y(n729) );
  OAI2BB2XL U1449 ( .B0(n2139), .B1(n2203), .A0N(\register[20][14] ), .A1N(
        n2204), .Y(n730) );
  OAI2BB2XL U1450 ( .B0(n2137), .B1(n2203), .A0N(\register[20][15] ), .A1N(
        n2204), .Y(n731) );
  OAI2BB2XL U1451 ( .B0(n2135), .B1(n2203), .A0N(\register[20][16] ), .A1N(
        n2204), .Y(n732) );
  OAI2BB2XL U1452 ( .B0(n2133), .B1(n2203), .A0N(\register[20][17] ), .A1N(
        n2203), .Y(n733) );
  OAI2BB2XL U1453 ( .B0(n2131), .B1(n2203), .A0N(\register[20][18] ), .A1N(
        n2202), .Y(n734) );
  OAI2BB2XL U1454 ( .B0(n2129), .B1(n2203), .A0N(\register[20][19] ), .A1N(
        n2204), .Y(n735) );
  OAI2BB2XL U1455 ( .B0(n2127), .B1(n2203), .A0N(\register[20][20] ), .A1N(
        n2203), .Y(n736) );
  OAI2BB2XL U1456 ( .B0(n2125), .B1(n2203), .A0N(\register[20][21] ), .A1N(
        n2202), .Y(n737) );
  OAI2BB2XL U1457 ( .B0(n2123), .B1(n2203), .A0N(\register[20][22] ), .A1N(
        n2204), .Y(n738) );
  OAI2BB2XL U1458 ( .B0(n2119), .B1(n2203), .A0N(\register[20][24] ), .A1N(
        n2204), .Y(n740) );
  OAI2BB2XL U1459 ( .B0(n2167), .B1(n2200), .A0N(\register[21][0] ), .A1N(
        n2200), .Y(n748) );
  OAI2BB2XL U1460 ( .B0(n2165), .B1(n2199), .A0N(\register[21][1] ), .A1N(
        n2199), .Y(n749) );
  OAI2BB2XL U1461 ( .B0(n2163), .B1(n2199), .A0N(\register[21][2] ), .A1N(
        n2200), .Y(n750) );
  OAI2BB2XL U1462 ( .B0(n2161), .B1(n2199), .A0N(\register[21][3] ), .A1N(
        n2201), .Y(n751) );
  OAI2BB2XL U1463 ( .B0(n2159), .B1(n2199), .A0N(\register[21][4] ), .A1N(
        n2199), .Y(n752) );
  OAI2BB2XL U1464 ( .B0(n2157), .B1(n2199), .A0N(\register[21][5] ), .A1N(
        n2201), .Y(n753) );
  OAI2BB2XL U1465 ( .B0(n2155), .B1(n2199), .A0N(\register[21][6] ), .A1N(
        n2201), .Y(n754) );
  OAI2BB2XL U1466 ( .B0(n2153), .B1(n2199), .A0N(\register[21][7] ), .A1N(
        n2201), .Y(n755) );
  OAI2BB2XL U1467 ( .B0(n2151), .B1(n2199), .A0N(\register[21][8] ), .A1N(
        n2201), .Y(n756) );
  OAI2BB2XL U1468 ( .B0(n2149), .B1(n2199), .A0N(\register[21][9] ), .A1N(
        n2201), .Y(n757) );
  OAI2BB2XL U1469 ( .B0(n2147), .B1(n2199), .A0N(\register[21][10] ), .A1N(
        n2201), .Y(n758) );
  OAI2BB2XL U1470 ( .B0(n2145), .B1(n2199), .A0N(\register[21][11] ), .A1N(
        n2201), .Y(n759) );
  OAI2BB2XL U1471 ( .B0(n2143), .B1(n2199), .A0N(\register[21][12] ), .A1N(
        n2201), .Y(n760) );
  OAI2BB2XL U1472 ( .B0(n2141), .B1(n2200), .A0N(\register[21][13] ), .A1N(
        n2201), .Y(n761) );
  OAI2BB2XL U1473 ( .B0(n2139), .B1(n2200), .A0N(\register[21][14] ), .A1N(
        n2201), .Y(n762) );
  OAI2BB2XL U1474 ( .B0(n2137), .B1(n2200), .A0N(\register[21][15] ), .A1N(
        n2201), .Y(n763) );
  OAI2BB2XL U1475 ( .B0(n2135), .B1(n2200), .A0N(\register[21][16] ), .A1N(
        n2201), .Y(n764) );
  OAI2BB2XL U1476 ( .B0(n2133), .B1(n2200), .A0N(\register[21][17] ), .A1N(
        n2200), .Y(n765) );
  OAI2BB2XL U1477 ( .B0(n2131), .B1(n2200), .A0N(\register[21][18] ), .A1N(
        n2199), .Y(n766) );
  OAI2BB2XL U1478 ( .B0(n2129), .B1(n2200), .A0N(\register[21][19] ), .A1N(
        n2201), .Y(n767) );
  OAI2BB2XL U1479 ( .B0(n2127), .B1(n2200), .A0N(\register[21][20] ), .A1N(
        n2200), .Y(n768) );
  OAI2BB2XL U1480 ( .B0(n2125), .B1(n2200), .A0N(\register[21][21] ), .A1N(
        n2199), .Y(n769) );
  OAI2BB2XL U1481 ( .B0(n2123), .B1(n2200), .A0N(\register[21][22] ), .A1N(
        n2201), .Y(n770) );
  OAI2BB2XL U1482 ( .B0(n2119), .B1(n2200), .A0N(\register[21][24] ), .A1N(
        n2201), .Y(n772) );
  OAI2BB2XL U1483 ( .B0(n2167), .B1(n2197), .A0N(\register[22][0] ), .A1N(
        n2197), .Y(n780) );
  OAI2BB2XL U1484 ( .B0(n2165), .B1(n2196), .A0N(\register[22][1] ), .A1N(
        n2196), .Y(n781) );
  OAI2BB2XL U1485 ( .B0(n2163), .B1(n2196), .A0N(\register[22][2] ), .A1N(
        n2197), .Y(n782) );
  OAI2BB2XL U1486 ( .B0(n2161), .B1(n2196), .A0N(\register[22][3] ), .A1N(
        n2198), .Y(n783) );
  OAI2BB2XL U1487 ( .B0(n2159), .B1(n2196), .A0N(\register[22][4] ), .A1N(
        n2196), .Y(n784) );
  OAI2BB2XL U1488 ( .B0(n2157), .B1(n2196), .A0N(\register[22][5] ), .A1N(
        n2198), .Y(n785) );
  OAI2BB2XL U1489 ( .B0(n2155), .B1(n2196), .A0N(\register[22][6] ), .A1N(
        n2198), .Y(n786) );
  OAI2BB2XL U1490 ( .B0(n2153), .B1(n2196), .A0N(\register[22][7] ), .A1N(
        n2198), .Y(n787) );
  OAI2BB2XL U1491 ( .B0(n2151), .B1(n2196), .A0N(\register[22][8] ), .A1N(
        n2198), .Y(n788) );
  OAI2BB2XL U1492 ( .B0(n2149), .B1(n2196), .A0N(\register[22][9] ), .A1N(
        n2198), .Y(n789) );
  OAI2BB2XL U1493 ( .B0(n2147), .B1(n2196), .A0N(\register[22][10] ), .A1N(
        n2198), .Y(n790) );
  OAI2BB2XL U1494 ( .B0(n2145), .B1(n2196), .A0N(\register[22][11] ), .A1N(
        n2198), .Y(n791) );
  OAI2BB2XL U1495 ( .B0(n2143), .B1(n2196), .A0N(\register[22][12] ), .A1N(
        n2198), .Y(n792) );
  OAI2BB2XL U1496 ( .B0(n2141), .B1(n2197), .A0N(\register[22][13] ), .A1N(
        n2198), .Y(n793) );
  OAI2BB2XL U1497 ( .B0(n2139), .B1(n2197), .A0N(\register[22][14] ), .A1N(
        n2198), .Y(n794) );
  OAI2BB2XL U1498 ( .B0(n2137), .B1(n2197), .A0N(\register[22][15] ), .A1N(
        n2198), .Y(n795) );
  OAI2BB2XL U1499 ( .B0(n2135), .B1(n2197), .A0N(\register[22][16] ), .A1N(
        n2198), .Y(n796) );
  OAI2BB2XL U1500 ( .B0(n2133), .B1(n2197), .A0N(\register[22][17] ), .A1N(
        n2197), .Y(n797) );
  OAI2BB2XL U1501 ( .B0(n2131), .B1(n2197), .A0N(\register[22][18] ), .A1N(
        n2196), .Y(n798) );
  OAI2BB2XL U1502 ( .B0(n2129), .B1(n2197), .A0N(\register[22][19] ), .A1N(
        n2198), .Y(n799) );
  OAI2BB2XL U1503 ( .B0(n2127), .B1(n2197), .A0N(\register[22][20] ), .A1N(
        n2197), .Y(n800) );
  OAI2BB2XL U1504 ( .B0(n2125), .B1(n2197), .A0N(\register[22][21] ), .A1N(
        n2196), .Y(n801) );
  OAI2BB2XL U1505 ( .B0(n2123), .B1(n2197), .A0N(\register[22][22] ), .A1N(
        n2198), .Y(n802) );
  OAI2BB2XL U1506 ( .B0(n2119), .B1(n2197), .A0N(\register[22][24] ), .A1N(
        n2198), .Y(n804) );
  OAI2BB2XL U1507 ( .B0(n2167), .B1(n2194), .A0N(\register[23][0] ), .A1N(
        n2194), .Y(n812) );
  OAI2BB2XL U1508 ( .B0(n2165), .B1(n2193), .A0N(\register[23][1] ), .A1N(
        n2193), .Y(n813) );
  OAI2BB2XL U1509 ( .B0(n2163), .B1(n2193), .A0N(\register[23][2] ), .A1N(
        n2194), .Y(n814) );
  OAI2BB2XL U1510 ( .B0(n2161), .B1(n2193), .A0N(\register[23][3] ), .A1N(
        n2195), .Y(n815) );
  OAI2BB2XL U1511 ( .B0(n2159), .B1(n2193), .A0N(\register[23][4] ), .A1N(
        n2193), .Y(n816) );
  OAI2BB2XL U1512 ( .B0(n2157), .B1(n2193), .A0N(\register[23][5] ), .A1N(
        n2195), .Y(n817) );
  OAI2BB2XL U1513 ( .B0(n2155), .B1(n2193), .A0N(\register[23][6] ), .A1N(
        n2195), .Y(n818) );
  OAI2BB2XL U1514 ( .B0(n2153), .B1(n2193), .A0N(\register[23][7] ), .A1N(
        n2195), .Y(n819) );
  OAI2BB2XL U1515 ( .B0(n2151), .B1(n2193), .A0N(\register[23][8] ), .A1N(
        n2195), .Y(n820) );
  OAI2BB2XL U1516 ( .B0(n2149), .B1(n2193), .A0N(\register[23][9] ), .A1N(
        n2195), .Y(n821) );
  OAI2BB2XL U1517 ( .B0(n2147), .B1(n2193), .A0N(\register[23][10] ), .A1N(
        n2195), .Y(n822) );
  OAI2BB2XL U1518 ( .B0(n2145), .B1(n2193), .A0N(\register[23][11] ), .A1N(
        n2195), .Y(n823) );
  OAI2BB2XL U1519 ( .B0(n2143), .B1(n2193), .A0N(\register[23][12] ), .A1N(
        n2195), .Y(n824) );
  OAI2BB2XL U1520 ( .B0(n2141), .B1(n2194), .A0N(\register[23][13] ), .A1N(
        n2195), .Y(n825) );
  OAI2BB2XL U1521 ( .B0(n2139), .B1(n2194), .A0N(\register[23][14] ), .A1N(
        n2195), .Y(n826) );
  OAI2BB2XL U1522 ( .B0(n2137), .B1(n2194), .A0N(\register[23][15] ), .A1N(
        n2195), .Y(n827) );
  OAI2BB2XL U1523 ( .B0(n2135), .B1(n2194), .A0N(\register[23][16] ), .A1N(
        n2195), .Y(n828) );
  OAI2BB2XL U1524 ( .B0(n2133), .B1(n2194), .A0N(\register[23][17] ), .A1N(
        n2194), .Y(n829) );
  OAI2BB2XL U1525 ( .B0(n2131), .B1(n2194), .A0N(\register[23][18] ), .A1N(
        n2193), .Y(n830) );
  OAI2BB2XL U1526 ( .B0(n2129), .B1(n2194), .A0N(\register[23][19] ), .A1N(
        n2195), .Y(n831) );
  OAI2BB2XL U1527 ( .B0(n2127), .B1(n2194), .A0N(\register[23][20] ), .A1N(
        n2194), .Y(n832) );
  OAI2BB2XL U1528 ( .B0(n2125), .B1(n2194), .A0N(\register[23][21] ), .A1N(
        n2193), .Y(n833) );
  OAI2BB2XL U1529 ( .B0(n2123), .B1(n2194), .A0N(\register[23][22] ), .A1N(
        n2195), .Y(n834) );
  OAI2BB2XL U1530 ( .B0(n2119), .B1(n2194), .A0N(\register[23][24] ), .A1N(
        n2195), .Y(n836) );
  OAI2BB2XL U1531 ( .B0(n2167), .B1(n2191), .A0N(\register[24][0] ), .A1N(
        n2191), .Y(n844) );
  OAI2BB2XL U1532 ( .B0(n2165), .B1(n2), .A0N(\register[24][1] ), .A1N(n2191), 
        .Y(n845) );
  OAI2BB2XL U1533 ( .B0(n2163), .B1(n2), .A0N(\register[24][2] ), .A1N(n2191), 
        .Y(n846) );
  OAI2BB2XL U1534 ( .B0(n2161), .B1(n2), .A0N(\register[24][3] ), .A1N(n2192), 
        .Y(n847) );
  OAI2BB2XL U1535 ( .B0(n2159), .B1(n2), .A0N(\register[24][4] ), .A1N(n2191), 
        .Y(n848) );
  OAI2BB2XL U1536 ( .B0(n2157), .B1(n2191), .A0N(\register[24][5] ), .A1N(
        n2192), .Y(n849) );
  OAI2BB2XL U1537 ( .B0(n2155), .B1(n2), .A0N(\register[24][6] ), .A1N(n2192), 
        .Y(n850) );
  OAI2BB2XL U1538 ( .B0(n2153), .B1(n2191), .A0N(\register[24][7] ), .A1N(
        n2192), .Y(n851) );
  OAI2BB2XL U1539 ( .B0(n2151), .B1(n2191), .A0N(\register[24][8] ), .A1N(
        n2192), .Y(n852) );
  OAI2BB2XL U1540 ( .B0(n2149), .B1(n2190), .A0N(\register[24][9] ), .A1N(
        n2192), .Y(n853) );
  OAI2BB2XL U1541 ( .B0(n2147), .B1(n2190), .A0N(\register[24][10] ), .A1N(
        n2192), .Y(n854) );
  OAI2BB2XL U1542 ( .B0(n2145), .B1(n2190), .A0N(\register[24][11] ), .A1N(
        n2192), .Y(n855) );
  OAI2BB2XL U1543 ( .B0(n2143), .B1(n2190), .A0N(\register[24][12] ), .A1N(
        n2192), .Y(n856) );
  OAI2BB2XL U1544 ( .B0(n2141), .B1(n2191), .A0N(\register[24][13] ), .A1N(
        n2192), .Y(n857) );
  OAI2BB2XL U1545 ( .B0(n2139), .B1(n2191), .A0N(\register[24][14] ), .A1N(
        n2192), .Y(n858) );
  OAI2BB2XL U1546 ( .B0(n2137), .B1(n2191), .A0N(\register[24][15] ), .A1N(
        n2190), .Y(n859) );
  OAI2BB2XL U1547 ( .B0(n2135), .B1(n2191), .A0N(\register[24][16] ), .A1N(
        n2192), .Y(n860) );
  OAI2BB2XL U1548 ( .B0(n2133), .B1(n2191), .A0N(\register[24][17] ), .A1N(
        n2190), .Y(n861) );
  OAI2BB2XL U1549 ( .B0(n2131), .B1(n2191), .A0N(\register[24][18] ), .A1N(
        n2190), .Y(n862) );
  OAI2BB2XL U1550 ( .B0(n2129), .B1(n2191), .A0N(\register[24][19] ), .A1N(
        n2190), .Y(n863) );
  OAI2BB2XL U1551 ( .B0(n2127), .B1(n2191), .A0N(\register[24][20] ), .A1N(
        n2190), .Y(n864) );
  OAI2BB2XL U1552 ( .B0(n2125), .B1(n2191), .A0N(\register[24][21] ), .A1N(
        n2190), .Y(n865) );
  OAI2BB2XL U1553 ( .B0(n2123), .B1(n2191), .A0N(\register[24][22] ), .A1N(
        n2192), .Y(n866) );
  OAI2BB2XL U1554 ( .B0(n2119), .B1(n2191), .A0N(\register[24][24] ), .A1N(
        n2192), .Y(n868) );
  OAI2BB2XL U1555 ( .B0(n2167), .B1(n2185), .A0N(\register[26][0] ), .A1N(
        n2185), .Y(n908) );
  OAI2BB2XL U1556 ( .B0(n2165), .B1(n3), .A0N(\register[26][1] ), .A1N(n2185), 
        .Y(n909) );
  OAI2BB2XL U1557 ( .B0(n2163), .B1(n3), .A0N(\register[26][2] ), .A1N(n2185), 
        .Y(n910) );
  OAI2BB2XL U1558 ( .B0(n2161), .B1(n3), .A0N(\register[26][3] ), .A1N(n2186), 
        .Y(n911) );
  OAI2BB2XL U1559 ( .B0(n2159), .B1(n3), .A0N(\register[26][4] ), .A1N(n2185), 
        .Y(n912) );
  OAI2BB2XL U1560 ( .B0(n2157), .B1(n2185), .A0N(\register[26][5] ), .A1N(
        n2186), .Y(n913) );
  OAI2BB2XL U1561 ( .B0(n2155), .B1(n3), .A0N(\register[26][6] ), .A1N(n2186), 
        .Y(n914) );
  OAI2BB2XL U1562 ( .B0(n2153), .B1(n2185), .A0N(\register[26][7] ), .A1N(
        n2186), .Y(n915) );
  OAI2BB2XL U1563 ( .B0(n2151), .B1(n2185), .A0N(\register[26][8] ), .A1N(
        n2186), .Y(n916) );
  OAI2BB2XL U1564 ( .B0(n2149), .B1(n2184), .A0N(\register[26][9] ), .A1N(
        n2186), .Y(n917) );
  OAI2BB2XL U1565 ( .B0(n2147), .B1(n2184), .A0N(\register[26][10] ), .A1N(
        n2186), .Y(n918) );
  OAI2BB2XL U1566 ( .B0(n2145), .B1(n2184), .A0N(\register[26][11] ), .A1N(
        n2186), .Y(n919) );
  OAI2BB2XL U1567 ( .B0(n2143), .B1(n2184), .A0N(\register[26][12] ), .A1N(
        n2186), .Y(n920) );
  OAI2BB2XL U1568 ( .B0(n2141), .B1(n2185), .A0N(\register[26][13] ), .A1N(
        n2186), .Y(n921) );
  OAI2BB2XL U1569 ( .B0(n2139), .B1(n2185), .A0N(\register[26][14] ), .A1N(
        n2186), .Y(n922) );
  OAI2BB2XL U1570 ( .B0(n2137), .B1(n2185), .A0N(\register[26][15] ), .A1N(
        n2184), .Y(n923) );
  OAI2BB2XL U1571 ( .B0(n2135), .B1(n2185), .A0N(\register[26][16] ), .A1N(
        n2186), .Y(n924) );
  OAI2BB2XL U1572 ( .B0(n2133), .B1(n2185), .A0N(\register[26][17] ), .A1N(
        n2184), .Y(n925) );
  OAI2BB2XL U1573 ( .B0(n2131), .B1(n2185), .A0N(\register[26][18] ), .A1N(
        n2184), .Y(n926) );
  OAI2BB2XL U1574 ( .B0(n2129), .B1(n2185), .A0N(\register[26][19] ), .A1N(
        n2184), .Y(n927) );
  OAI2BB2XL U1575 ( .B0(n2127), .B1(n2185), .A0N(\register[26][20] ), .A1N(
        n2184), .Y(n928) );
  OAI2BB2XL U1576 ( .B0(n2125), .B1(n2185), .A0N(\register[26][21] ), .A1N(
        n2184), .Y(n929) );
  OAI2BB2XL U1577 ( .B0(n2123), .B1(n2185), .A0N(\register[26][22] ), .A1N(
        n2186), .Y(n930) );
  OAI2BB2XL U1578 ( .B0(n2119), .B1(n2185), .A0N(\register[26][24] ), .A1N(
        n2186), .Y(n932) );
  OAI2BB2XL U1579 ( .B0(n2167), .B1(n2182), .A0N(\register[27][0] ), .A1N(
        n2182), .Y(n940) );
  OAI2BB2XL U1580 ( .B0(n2165), .B1(n4), .A0N(\register[27][1] ), .A1N(n2182), 
        .Y(n941) );
  OAI2BB2XL U1581 ( .B0(n2163), .B1(n4), .A0N(\register[27][2] ), .A1N(n2182), 
        .Y(n942) );
  OAI2BB2XL U1582 ( .B0(n2161), .B1(n4), .A0N(\register[27][3] ), .A1N(n2183), 
        .Y(n943) );
  OAI2BB2XL U1583 ( .B0(n2159), .B1(n4), .A0N(\register[27][4] ), .A1N(n2182), 
        .Y(n944) );
  OAI2BB2XL U1584 ( .B0(n2157), .B1(n2182), .A0N(\register[27][5] ), .A1N(
        n2183), .Y(n945) );
  OAI2BB2XL U1585 ( .B0(n2155), .B1(n4), .A0N(\register[27][6] ), .A1N(n2183), 
        .Y(n946) );
  OAI2BB2XL U1586 ( .B0(n2153), .B1(n2182), .A0N(\register[27][7] ), .A1N(
        n2183), .Y(n947) );
  OAI2BB2XL U1587 ( .B0(n2151), .B1(n2182), .A0N(\register[27][8] ), .A1N(
        n2183), .Y(n948) );
  OAI2BB2XL U1588 ( .B0(n2149), .B1(n2181), .A0N(\register[27][9] ), .A1N(
        n2183), .Y(n949) );
  OAI2BB2XL U1589 ( .B0(n2147), .B1(n2181), .A0N(\register[27][10] ), .A1N(
        n2183), .Y(n950) );
  OAI2BB2XL U1590 ( .B0(n2145), .B1(n2181), .A0N(\register[27][11] ), .A1N(
        n2183), .Y(n951) );
  OAI2BB2XL U1591 ( .B0(n2143), .B1(n2181), .A0N(\register[27][12] ), .A1N(
        n2183), .Y(n952) );
  OAI2BB2XL U1592 ( .B0(n2141), .B1(n2182), .A0N(\register[27][13] ), .A1N(
        n2183), .Y(n953) );
  OAI2BB2XL U1593 ( .B0(n2139), .B1(n2182), .A0N(\register[27][14] ), .A1N(
        n2183), .Y(n954) );
  OAI2BB2XL U1594 ( .B0(n2137), .B1(n2182), .A0N(\register[27][15] ), .A1N(
        n2181), .Y(n955) );
  OAI2BB2XL U1595 ( .B0(n2135), .B1(n2182), .A0N(\register[27][16] ), .A1N(
        n2183), .Y(n956) );
  OAI2BB2XL U1596 ( .B0(n2133), .B1(n2182), .A0N(\register[27][17] ), .A1N(
        n2181), .Y(n957) );
  OAI2BB2XL U1597 ( .B0(n2131), .B1(n2182), .A0N(\register[27][18] ), .A1N(
        n2181), .Y(n958) );
  OAI2BB2XL U1598 ( .B0(n2129), .B1(n2182), .A0N(\register[27][19] ), .A1N(
        n2181), .Y(n959) );
  OAI2BB2XL U1599 ( .B0(n2127), .B1(n2182), .A0N(\register[27][20] ), .A1N(
        n2181), .Y(n960) );
  OAI2BB2XL U1600 ( .B0(n2125), .B1(n2182), .A0N(\register[27][21] ), .A1N(
        n2181), .Y(n961) );
  OAI2BB2XL U1601 ( .B0(n2123), .B1(n2182), .A0N(\register[27][22] ), .A1N(
        n2183), .Y(n962) );
  OAI2BB2XL U1602 ( .B0(n2119), .B1(n2182), .A0N(\register[27][24] ), .A1N(
        n2183), .Y(n964) );
  OAI2BB2XL U1603 ( .B0(n2167), .B1(n2179), .A0N(\register[28][0] ), .A1N(
        n2179), .Y(n972) );
  OAI2BB2XL U1604 ( .B0(n2165), .B1(n5), .A0N(\register[28][1] ), .A1N(n2179), 
        .Y(n973) );
  OAI2BB2XL U1605 ( .B0(n2163), .B1(n5), .A0N(\register[28][2] ), .A1N(n2179), 
        .Y(n974) );
  OAI2BB2XL U1606 ( .B0(n2161), .B1(n5), .A0N(\register[28][3] ), .A1N(n2180), 
        .Y(n975) );
  OAI2BB2XL U1607 ( .B0(n2159), .B1(n5), .A0N(\register[28][4] ), .A1N(n2179), 
        .Y(n976) );
  OAI2BB2XL U1608 ( .B0(n2157), .B1(n2179), .A0N(\register[28][5] ), .A1N(
        n2180), .Y(n977) );
  OAI2BB2XL U1609 ( .B0(n2155), .B1(n5), .A0N(\register[28][6] ), .A1N(n2180), 
        .Y(n978) );
  OAI2BB2XL U1610 ( .B0(n2153), .B1(n2179), .A0N(\register[28][7] ), .A1N(
        n2180), .Y(n979) );
  OAI2BB2XL U1611 ( .B0(n2151), .B1(n2179), .A0N(\register[28][8] ), .A1N(
        n2180), .Y(n980) );
  OAI2BB2XL U1612 ( .B0(n2149), .B1(n2178), .A0N(\register[28][9] ), .A1N(
        n2180), .Y(n981) );
  OAI2BB2XL U1613 ( .B0(n2147), .B1(n2178), .A0N(\register[28][10] ), .A1N(
        n2180), .Y(n982) );
  OAI2BB2XL U1614 ( .B0(n2145), .B1(n2178), .A0N(\register[28][11] ), .A1N(
        n2180), .Y(n983) );
  OAI2BB2XL U1615 ( .B0(n2143), .B1(n2178), .A0N(\register[28][12] ), .A1N(
        n2180), .Y(n984) );
  OAI2BB2XL U1616 ( .B0(n2141), .B1(n2179), .A0N(\register[28][13] ), .A1N(
        n2180), .Y(n985) );
  OAI2BB2XL U1617 ( .B0(n2139), .B1(n2179), .A0N(\register[28][14] ), .A1N(
        n2180), .Y(n986) );
  OAI2BB2XL U1618 ( .B0(n2137), .B1(n2179), .A0N(\register[28][15] ), .A1N(
        n2178), .Y(n987) );
  OAI2BB2XL U1619 ( .B0(n2135), .B1(n2179), .A0N(\register[28][16] ), .A1N(
        n2180), .Y(n988) );
  OAI2BB2XL U1620 ( .B0(n2133), .B1(n2179), .A0N(\register[28][17] ), .A1N(
        n2178), .Y(n989) );
  OAI2BB2XL U1621 ( .B0(n2131), .B1(n2179), .A0N(\register[28][18] ), .A1N(
        n2178), .Y(n990) );
  OAI2BB2XL U1622 ( .B0(n2129), .B1(n2179), .A0N(\register[28][19] ), .A1N(
        n2178), .Y(n991) );
  OAI2BB2XL U1623 ( .B0(n2127), .B1(n2179), .A0N(\register[28][20] ), .A1N(
        n2178), .Y(n992) );
  OAI2BB2XL U1624 ( .B0(n2125), .B1(n2179), .A0N(\register[28][21] ), .A1N(
        n2178), .Y(n993) );
  OAI2BB2XL U1625 ( .B0(n2123), .B1(n2179), .A0N(\register[28][22] ), .A1N(
        n2180), .Y(n994) );
  OAI2BB2XL U1626 ( .B0(n2119), .B1(n2179), .A0N(\register[28][24] ), .A1N(
        n2180), .Y(n996) );
  OAI2BB2XL U1627 ( .B0(n2168), .B1(n2176), .A0N(\register[29][0] ), .A1N(
        n2176), .Y(n1004) );
  OAI2BB2XL U1628 ( .B0(n2165), .B1(n2176), .A0N(\register[29][1] ), .A1N(
        n2176), .Y(n1005) );
  OAI2BB2XL U1629 ( .B0(n2163), .B1(n2176), .A0N(\register[29][2] ), .A1N(
        n2176), .Y(n1006) );
  OAI2BB2XL U1630 ( .B0(n2161), .B1(n2176), .A0N(\register[29][3] ), .A1N(
        n2177), .Y(n1007) );
  OAI2BB2XL U1631 ( .B0(n2159), .B1(n2175), .A0N(\register[29][4] ), .A1N(
        n2176), .Y(n1008) );
  OAI2BB2XL U1632 ( .B0(n2158), .B1(n6), .A0N(\register[29][5] ), .A1N(n2177), 
        .Y(n1009) );
  OAI2BB2XL U1633 ( .B0(n2155), .B1(n2175), .A0N(\register[29][6] ), .A1N(
        n2177), .Y(n1010) );
  OAI2BB2XL U1634 ( .B0(n2154), .B1(n6), .A0N(\register[29][7] ), .A1N(n2177), 
        .Y(n1011) );
  OAI2BB2XL U1635 ( .B0(n2152), .B1(n6), .A0N(\register[29][8] ), .A1N(n2177), 
        .Y(n1012) );
  OAI2BB2XL U1636 ( .B0(n2150), .B1(n2175), .A0N(\register[29][9] ), .A1N(
        n2177), .Y(n1013) );
  OAI2BB2XL U1637 ( .B0(n2148), .B1(n2175), .A0N(\register[29][10] ), .A1N(
        n2177), .Y(n1014) );
  OAI2BB2XL U1638 ( .B0(n2145), .B1(n6), .A0N(\register[29][11] ), .A1N(n2177), 
        .Y(n1015) );
  OAI2BB2XL U1639 ( .B0(n2143), .B1(n6), .A0N(\register[29][12] ), .A1N(n2177), 
        .Y(n1016) );
  OAI2BB2XL U1640 ( .B0(n2141), .B1(n2176), .A0N(\register[29][13] ), .A1N(
        n2177), .Y(n1017) );
  OAI2BB2XL U1641 ( .B0(n2139), .B1(n2176), .A0N(\register[29][14] ), .A1N(
        n2177), .Y(n1018) );
  OAI2BB2XL U1642 ( .B0(n2137), .B1(n2176), .A0N(\register[29][15] ), .A1N(
        n2175), .Y(n1019) );
  OAI2BB2XL U1643 ( .B0(n2135), .B1(n2176), .A0N(\register[29][16] ), .A1N(
        n2177), .Y(n1020) );
  OAI2BB2XL U1644 ( .B0(n2133), .B1(n2176), .A0N(\register[29][17] ), .A1N(
        n2175), .Y(n1021) );
  OAI2BB2XL U1645 ( .B0(n2131), .B1(n2176), .A0N(\register[29][18] ), .A1N(
        n2175), .Y(n1022) );
  OAI2BB2XL U1646 ( .B0(n2129), .B1(n2176), .A0N(\register[29][19] ), .A1N(
        n2175), .Y(n1023) );
  OAI2BB2XL U1647 ( .B0(n2127), .B1(n2176), .A0N(\register[29][20] ), .A1N(
        n2175), .Y(n1024) );
  OAI2BB2XL U1648 ( .B0(n2125), .B1(n2176), .A0N(\register[29][21] ), .A1N(
        n2175), .Y(n1025) );
  OAI2BB2XL U1649 ( .B0(n2123), .B1(n2176), .A0N(\register[29][22] ), .A1N(
        n2177), .Y(n1026) );
  OAI2BB2XL U1650 ( .B0(n2119), .B1(n2176), .A0N(\register[29][24] ), .A1N(
        n2177), .Y(n1028) );
  OAI2BB2XL U1651 ( .B0(n2168), .B1(n2173), .A0N(\register[30][0] ), .A1N(
        n2173), .Y(n1036) );
  OAI2BB2XL U1652 ( .B0(n2165), .B1(n2173), .A0N(\register[30][1] ), .A1N(
        n2173), .Y(n1037) );
  OAI2BB2XL U1653 ( .B0(n2163), .B1(n2173), .A0N(\register[30][2] ), .A1N(
        n2173), .Y(n1038) );
  OAI2BB2XL U1654 ( .B0(n2161), .B1(n2173), .A0N(\register[30][3] ), .A1N(
        n2174), .Y(n1039) );
  OAI2BB2XL U1655 ( .B0(n2159), .B1(n2172), .A0N(\register[30][4] ), .A1N(
        n2173), .Y(n1040) );
  OAI2BB2XL U1656 ( .B0(n2158), .B1(n7), .A0N(\register[30][5] ), .A1N(n2174), 
        .Y(n1041) );
  OAI2BB2XL U1657 ( .B0(n2155), .B1(n2172), .A0N(\register[30][6] ), .A1N(
        n2174), .Y(n1042) );
  OAI2BB2XL U1658 ( .B0(n2154), .B1(n7), .A0N(\register[30][7] ), .A1N(n2174), 
        .Y(n1043) );
  OAI2BB2XL U1659 ( .B0(n2152), .B1(n7), .A0N(\register[30][8] ), .A1N(n2174), 
        .Y(n1044) );
  OAI2BB2XL U1660 ( .B0(n2150), .B1(n2172), .A0N(\register[30][9] ), .A1N(
        n2174), .Y(n1045) );
  OAI2BB2XL U1661 ( .B0(n2148), .B1(n2172), .A0N(\register[30][10] ), .A1N(
        n2174), .Y(n1046) );
  OAI2BB2XL U1662 ( .B0(n2145), .B1(n7), .A0N(\register[30][11] ), .A1N(n2174), 
        .Y(n1047) );
  OAI2BB2XL U1663 ( .B0(n2143), .B1(n7), .A0N(\register[30][12] ), .A1N(n2174), 
        .Y(n1048) );
  OAI2BB2XL U1664 ( .B0(n2141), .B1(n2173), .A0N(\register[30][13] ), .A1N(
        n2174), .Y(n1049) );
  OAI2BB2XL U1665 ( .B0(n2139), .B1(n2173), .A0N(\register[30][14] ), .A1N(
        n2174), .Y(n1050) );
  OAI2BB2XL U1666 ( .B0(n2137), .B1(n2173), .A0N(\register[30][15] ), .A1N(
        n2172), .Y(n1051) );
  OAI2BB2XL U1667 ( .B0(n2135), .B1(n2173), .A0N(\register[30][16] ), .A1N(
        n2174), .Y(n1052) );
  OAI2BB2XL U1668 ( .B0(n2133), .B1(n2173), .A0N(\register[30][17] ), .A1N(
        n2172), .Y(n1053) );
  OAI2BB2XL U1669 ( .B0(n2131), .B1(n2173), .A0N(\register[30][18] ), .A1N(
        n2172), .Y(n1054) );
  OAI2BB2XL U1670 ( .B0(n2129), .B1(n2173), .A0N(\register[30][19] ), .A1N(
        n2172), .Y(n1055) );
  OAI2BB2XL U1671 ( .B0(n2127), .B1(n2173), .A0N(\register[30][20] ), .A1N(
        n2172), .Y(n1056) );
  OAI2BB2XL U1672 ( .B0(n2125), .B1(n2173), .A0N(\register[30][21] ), .A1N(
        n2172), .Y(n1057) );
  OAI2BB2XL U1673 ( .B0(n2123), .B1(n2173), .A0N(\register[30][22] ), .A1N(
        n2174), .Y(n1058) );
  OAI2BB2XL U1674 ( .B0(n2119), .B1(n2173), .A0N(\register[30][24] ), .A1N(
        n2174), .Y(n1060) );
  OAI2BB2XL U1675 ( .B0(n2168), .B1(n2170), .A0N(\register[31][0] ), .A1N(
        n2170), .Y(n1068) );
  OAI2BB2XL U1676 ( .B0(n2165), .B1(n2170), .A0N(\register[31][1] ), .A1N(
        n2170), .Y(n1069) );
  OAI2BB2XL U1677 ( .B0(n2163), .B1(n2170), .A0N(\register[31][2] ), .A1N(
        n2170), .Y(n1070) );
  OAI2BB2XL U1678 ( .B0(n2161), .B1(n2170), .A0N(\register[31][3] ), .A1N(
        n2171), .Y(n1071) );
  OAI2BB2XL U1679 ( .B0(n2159), .B1(n2169), .A0N(\register[31][4] ), .A1N(
        n2170), .Y(n1072) );
  OAI2BB2XL U1680 ( .B0(n2158), .B1(n8), .A0N(\register[31][5] ), .A1N(n2171), 
        .Y(n1073) );
  OAI2BB2XL U1681 ( .B0(n2155), .B1(n2169), .A0N(\register[31][6] ), .A1N(
        n2171), .Y(n1074) );
  OAI2BB2XL U1682 ( .B0(n2154), .B1(n8), .A0N(\register[31][7] ), .A1N(n2171), 
        .Y(n1075) );
  OAI2BB2XL U1683 ( .B0(n2152), .B1(n8), .A0N(\register[31][8] ), .A1N(n2171), 
        .Y(n1076) );
  OAI2BB2XL U1684 ( .B0(n2150), .B1(n2169), .A0N(\register[31][9] ), .A1N(
        n2171), .Y(n1077) );
  OAI2BB2XL U1685 ( .B0(n2439), .B1(n2169), .A0N(\register[31][10] ), .A1N(
        n2171), .Y(n1078) );
  OAI2BB2XL U1686 ( .B0(n2145), .B1(n8), .A0N(\register[31][11] ), .A1N(n2171), 
        .Y(n1079) );
  OAI2BB2XL U1687 ( .B0(n2143), .B1(n8), .A0N(\register[31][12] ), .A1N(n2171), 
        .Y(n1080) );
  OAI2BB2XL U1688 ( .B0(n2141), .B1(n2170), .A0N(\register[31][13] ), .A1N(
        n2171), .Y(n1081) );
  OAI2BB2XL U1689 ( .B0(n2139), .B1(n2170), .A0N(\register[31][14] ), .A1N(
        n2171), .Y(n1082) );
  OAI2BB2XL U1690 ( .B0(n2137), .B1(n2170), .A0N(\register[31][15] ), .A1N(
        n2169), .Y(n1083) );
  OAI2BB2XL U1691 ( .B0(n2135), .B1(n2170), .A0N(\register[31][16] ), .A1N(
        n2171), .Y(n1084) );
  OAI2BB2XL U1692 ( .B0(n2133), .B1(n2170), .A0N(\register[31][17] ), .A1N(
        n2169), .Y(n1085) );
  OAI2BB2XL U1693 ( .B0(n2131), .B1(n2170), .A0N(\register[31][18] ), .A1N(
        n2169), .Y(n1086) );
  OAI2BB2XL U1694 ( .B0(n2129), .B1(n2170), .A0N(\register[31][19] ), .A1N(
        n2169), .Y(n1087) );
  OAI2BB2XL U1695 ( .B0(n2127), .B1(n2170), .A0N(\register[31][20] ), .A1N(
        n2169), .Y(n1088) );
  OAI2BB2XL U1696 ( .B0(n2125), .B1(n2170), .A0N(\register[31][21] ), .A1N(
        n2169), .Y(n1089) );
  OAI2BB2XL U1697 ( .B0(n2123), .B1(n2170), .A0N(\register[31][22] ), .A1N(
        n2171), .Y(n1090) );
  OAI2BB2XL U1698 ( .B0(n2119), .B1(n2170), .A0N(\register[31][24] ), .A1N(
        n2171), .Y(n1092) );
  OAI2BB2XL U1699 ( .B0(n2168), .B1(n2257), .A0N(\register[2][0] ), .A1N(n2257), .Y(n140) );
  OAI2BB2XL U1700 ( .B0(n2165), .B1(n2256), .A0N(\register[2][1] ), .A1N(n2256), .Y(n141) );
  OAI2BB2XL U1701 ( .B0(n2163), .B1(n2256), .A0N(\register[2][2] ), .A1N(n2257), .Y(n142) );
  OAI2BB2XL U1702 ( .B0(n2161), .B1(n2256), .A0N(\register[2][3] ), .A1N(n2258), .Y(n143) );
  OAI2BB2XL U1703 ( .B0(n2159), .B1(n2256), .A0N(\register[2][4] ), .A1N(n2256), .Y(n144) );
  OAI2BB2XL U1704 ( .B0(n2158), .B1(n2256), .A0N(\register[2][5] ), .A1N(n2258), .Y(n145) );
  OAI2BB2XL U1705 ( .B0(n2155), .B1(n2256), .A0N(\register[2][6] ), .A1N(n2258), .Y(n146) );
  OAI2BB2XL U1706 ( .B0(n2154), .B1(n2256), .A0N(\register[2][7] ), .A1N(n2258), .Y(n147) );
  OAI2BB2XL U1707 ( .B0(n2152), .B1(n2256), .A0N(\register[2][8] ), .A1N(n2258), .Y(n148) );
  OAI2BB2XL U1708 ( .B0(n2150), .B1(n2256), .A0N(\register[2][9] ), .A1N(n2258), .Y(n149) );
  OAI2BB2XL U1709 ( .B0(n2148), .B1(n2256), .A0N(\register[2][10] ), .A1N(
        n2258), .Y(n150) );
  OAI2BB2XL U1710 ( .B0(n2145), .B1(n2256), .A0N(\register[2][11] ), .A1N(
        n2258), .Y(n151) );
  OAI2BB2XL U1711 ( .B0(n2143), .B1(n2256), .A0N(\register[2][12] ), .A1N(
        n2258), .Y(n152) );
  OAI2BB2XL U1712 ( .B0(n2141), .B1(n2257), .A0N(\register[2][13] ), .A1N(
        n2258), .Y(n153) );
  OAI2BB2XL U1713 ( .B0(n2139), .B1(n2257), .A0N(\register[2][14] ), .A1N(
        n2258), .Y(n154) );
  OAI2BB2XL U1714 ( .B0(n2137), .B1(n2257), .A0N(\register[2][15] ), .A1N(
        n2258), .Y(n155) );
  OAI2BB2XL U1715 ( .B0(n2135), .B1(n2257), .A0N(\register[2][16] ), .A1N(
        n2258), .Y(n156) );
  OAI2BB2XL U1716 ( .B0(n2133), .B1(n2257), .A0N(\register[2][17] ), .A1N(
        n2256), .Y(n157) );
  OAI2BB2XL U1717 ( .B0(n2131), .B1(n2257), .A0N(\register[2][18] ), .A1N(
        n2257), .Y(n158) );
  OAI2BB2XL U1718 ( .B0(n2129), .B1(n2257), .A0N(\register[2][19] ), .A1N(
        n2258), .Y(n159) );
  OAI2BB2XL U1719 ( .B0(n2127), .B1(n2257), .A0N(\register[2][20] ), .A1N(
        n2256), .Y(n160) );
  OAI2BB2XL U1720 ( .B0(n2125), .B1(n2257), .A0N(\register[2][21] ), .A1N(
        n2257), .Y(n161) );
  OAI2BB2XL U1721 ( .B0(n2123), .B1(n2257), .A0N(\register[2][22] ), .A1N(
        n2258), .Y(n162) );
  OAI2BB2XL U1722 ( .B0(n2119), .B1(n2257), .A0N(\register[2][24] ), .A1N(
        n2258), .Y(n164) );
  OAI2BB2XL U1723 ( .B0(n2168), .B1(n2254), .A0N(\register[3][0] ), .A1N(n2254), .Y(n172) );
  OAI2BB2XL U1724 ( .B0(n2165), .B1(n2253), .A0N(\register[3][1] ), .A1N(n2253), .Y(n173) );
  OAI2BB2XL U1725 ( .B0(n2163), .B1(n2253), .A0N(\register[3][2] ), .A1N(n2254), .Y(n174) );
  OAI2BB2XL U1726 ( .B0(n2161), .B1(n2253), .A0N(\register[3][3] ), .A1N(n2255), .Y(n175) );
  OAI2BB2XL U1727 ( .B0(n2159), .B1(n2253), .A0N(\register[3][4] ), .A1N(n2253), .Y(n176) );
  OAI2BB2XL U1728 ( .B0(n2158), .B1(n2253), .A0N(\register[3][5] ), .A1N(n2255), .Y(n177) );
  OAI2BB2XL U1729 ( .B0(n2155), .B1(n2253), .A0N(\register[3][6] ), .A1N(n2255), .Y(n178) );
  OAI2BB2XL U1730 ( .B0(n2154), .B1(n2253), .A0N(\register[3][7] ), .A1N(n2255), .Y(n179) );
  OAI2BB2XL U1731 ( .B0(n2152), .B1(n2253), .A0N(\register[3][8] ), .A1N(n2255), .Y(n180) );
  OAI2BB2XL U1732 ( .B0(n2150), .B1(n2253), .A0N(\register[3][9] ), .A1N(n2255), .Y(n181) );
  OAI2BB2XL U1733 ( .B0(n2148), .B1(n2253), .A0N(\register[3][10] ), .A1N(
        n2255), .Y(n182) );
  OAI2BB2XL U1734 ( .B0(n2145), .B1(n2253), .A0N(\register[3][11] ), .A1N(
        n2255), .Y(n183) );
  OAI2BB2XL U1735 ( .B0(n2143), .B1(n2253), .A0N(\register[3][12] ), .A1N(
        n2255), .Y(n184) );
  OAI2BB2XL U1736 ( .B0(n2141), .B1(n2254), .A0N(\register[3][13] ), .A1N(
        n2255), .Y(n185) );
  OAI2BB2XL U1737 ( .B0(n2139), .B1(n2254), .A0N(\register[3][14] ), .A1N(
        n2255), .Y(n186) );
  OAI2BB2XL U1738 ( .B0(n2137), .B1(n2254), .A0N(\register[3][15] ), .A1N(
        n2255), .Y(n187) );
  OAI2BB2XL U1739 ( .B0(n2135), .B1(n2254), .A0N(\register[3][16] ), .A1N(
        n2255), .Y(n188) );
  OAI2BB2XL U1740 ( .B0(n2133), .B1(n2254), .A0N(\register[3][17] ), .A1N(
        n2253), .Y(n189) );
  OAI2BB2XL U1741 ( .B0(n2131), .B1(n2254), .A0N(\register[3][18] ), .A1N(
        n2254), .Y(n190) );
  OAI2BB2XL U1742 ( .B0(n2129), .B1(n2254), .A0N(\register[3][19] ), .A1N(
        n2255), .Y(n191) );
  OAI2BB2XL U1743 ( .B0(n2127), .B1(n2254), .A0N(\register[3][20] ), .A1N(
        n2253), .Y(n192) );
  OAI2BB2XL U1744 ( .B0(n2125), .B1(n2254), .A0N(\register[3][21] ), .A1N(
        n2254), .Y(n193) );
  OAI2BB2XL U1745 ( .B0(n2123), .B1(n2254), .A0N(\register[3][22] ), .A1N(
        n2255), .Y(n194) );
  OAI2BB2XL U1746 ( .B0(n2119), .B1(n2254), .A0N(\register[3][24] ), .A1N(
        n2255), .Y(n196) );
  OAI2BB2XL U1747 ( .B0(n2168), .B1(n2251), .A0N(\register[4][0] ), .A1N(n2251), .Y(n204) );
  OAI2BB2XL U1748 ( .B0(n2165), .B1(n2250), .A0N(\register[4][1] ), .A1N(n2250), .Y(n205) );
  OAI2BB2XL U1749 ( .B0(n2163), .B1(n2250), .A0N(\register[4][2] ), .A1N(n2251), .Y(n206) );
  OAI2BB2XL U1750 ( .B0(n2161), .B1(n2250), .A0N(\register[4][3] ), .A1N(n2252), .Y(n207) );
  OAI2BB2XL U1751 ( .B0(n2159), .B1(n2250), .A0N(\register[4][4] ), .A1N(n2250), .Y(n208) );
  OAI2BB2XL U1752 ( .B0(n2158), .B1(n2250), .A0N(\register[4][5] ), .A1N(n2252), .Y(n209) );
  OAI2BB2XL U1753 ( .B0(n2155), .B1(n2250), .A0N(\register[4][6] ), .A1N(n2252), .Y(n210) );
  OAI2BB2XL U1754 ( .B0(n2154), .B1(n2250), .A0N(\register[4][7] ), .A1N(n2252), .Y(n211) );
  OAI2BB2XL U1755 ( .B0(n2152), .B1(n2250), .A0N(\register[4][8] ), .A1N(n2252), .Y(n212) );
  OAI2BB2XL U1756 ( .B0(n2150), .B1(n2250), .A0N(\register[4][9] ), .A1N(n2252), .Y(n213) );
  OAI2BB2XL U1757 ( .B0(n2148), .B1(n2250), .A0N(\register[4][10] ), .A1N(
        n2252), .Y(n214) );
  OAI2BB2XL U1758 ( .B0(n2145), .B1(n2250), .A0N(\register[4][11] ), .A1N(
        n2252), .Y(n215) );
  OAI2BB2XL U1759 ( .B0(n2143), .B1(n2250), .A0N(\register[4][12] ), .A1N(
        n2252), .Y(n216) );
  OAI2BB2XL U1760 ( .B0(n2141), .B1(n2251), .A0N(\register[4][13] ), .A1N(
        n2252), .Y(n217) );
  OAI2BB2XL U1761 ( .B0(n2139), .B1(n2251), .A0N(\register[4][14] ), .A1N(
        n2252), .Y(n218) );
  OAI2BB2XL U1762 ( .B0(n2137), .B1(n2251), .A0N(\register[4][15] ), .A1N(
        n2252), .Y(n219) );
  OAI2BB2XL U1763 ( .B0(n2135), .B1(n2251), .A0N(\register[4][16] ), .A1N(
        n2252), .Y(n220) );
  OAI2BB2XL U1764 ( .B0(n2133), .B1(n2251), .A0N(\register[4][17] ), .A1N(
        n2250), .Y(n221) );
  OAI2BB2XL U1765 ( .B0(n2131), .B1(n2251), .A0N(\register[4][18] ), .A1N(
        n2251), .Y(n222) );
  OAI2BB2XL U1766 ( .B0(n2129), .B1(n2251), .A0N(\register[4][19] ), .A1N(
        n2252), .Y(n223) );
  OAI2BB2XL U1767 ( .B0(n2127), .B1(n2251), .A0N(\register[4][20] ), .A1N(
        n2250), .Y(n224) );
  OAI2BB2XL U1768 ( .B0(n2125), .B1(n2251), .A0N(\register[4][21] ), .A1N(
        n2251), .Y(n225) );
  OAI2BB2XL U1769 ( .B0(n2123), .B1(n2251), .A0N(\register[4][22] ), .A1N(
        n2252), .Y(n226) );
  OAI2BB2XL U1770 ( .B0(n2119), .B1(n2251), .A0N(\register[4][24] ), .A1N(
        n2252), .Y(n228) );
  OAI2BB2XL U1771 ( .B0(n2168), .B1(n2248), .A0N(\register[5][0] ), .A1N(n2248), .Y(n236) );
  OAI2BB2XL U1772 ( .B0(n2165), .B1(n2247), .A0N(\register[5][1] ), .A1N(n2247), .Y(n237) );
  OAI2BB2XL U1773 ( .B0(n2163), .B1(n2247), .A0N(\register[5][2] ), .A1N(n2248), .Y(n238) );
  OAI2BB2XL U1774 ( .B0(n2161), .B1(n2247), .A0N(\register[5][3] ), .A1N(n2249), .Y(n239) );
  OAI2BB2XL U1775 ( .B0(n2159), .B1(n2247), .A0N(\register[5][4] ), .A1N(n2247), .Y(n240) );
  OAI2BB2XL U1776 ( .B0(n2158), .B1(n2247), .A0N(\register[5][5] ), .A1N(n2249), .Y(n241) );
  OAI2BB2XL U1777 ( .B0(n2155), .B1(n2247), .A0N(\register[5][6] ), .A1N(n2249), .Y(n242) );
  OAI2BB2XL U1778 ( .B0(n2154), .B1(n2247), .A0N(\register[5][7] ), .A1N(n2249), .Y(n243) );
  OAI2BB2XL U1779 ( .B0(n2152), .B1(n2247), .A0N(\register[5][8] ), .A1N(n2249), .Y(n244) );
  OAI2BB2XL U1780 ( .B0(n2150), .B1(n2247), .A0N(\register[5][9] ), .A1N(n2249), .Y(n245) );
  OAI2BB2XL U1781 ( .B0(n2148), .B1(n2247), .A0N(\register[5][10] ), .A1N(
        n2249), .Y(n246) );
  OAI2BB2XL U1782 ( .B0(n2145), .B1(n2247), .A0N(\register[5][11] ), .A1N(
        n2249), .Y(n247) );
  OAI2BB2XL U1783 ( .B0(n2143), .B1(n2247), .A0N(\register[5][12] ), .A1N(
        n2249), .Y(n248) );
  OAI2BB2XL U1784 ( .B0(n2141), .B1(n2248), .A0N(\register[5][13] ), .A1N(
        n2249), .Y(n249) );
  OAI2BB2XL U1785 ( .B0(n2139), .B1(n2248), .A0N(\register[5][14] ), .A1N(
        n2249), .Y(n250) );
  OAI2BB2XL U1786 ( .B0(n2137), .B1(n2248), .A0N(\register[5][15] ), .A1N(
        n2249), .Y(n251) );
  OAI2BB2XL U1787 ( .B0(n2135), .B1(n2248), .A0N(\register[5][16] ), .A1N(
        n2249), .Y(n252) );
  OAI2BB2XL U1788 ( .B0(n2133), .B1(n2248), .A0N(\register[5][17] ), .A1N(
        n2247), .Y(n253) );
  OAI2BB2XL U1789 ( .B0(n2131), .B1(n2248), .A0N(\register[5][18] ), .A1N(
        n2248), .Y(n254) );
  OAI2BB2XL U1790 ( .B0(n2129), .B1(n2248), .A0N(\register[5][19] ), .A1N(
        n2249), .Y(n255) );
  OAI2BB2XL U1791 ( .B0(n2127), .B1(n2248), .A0N(\register[5][20] ), .A1N(
        n2247), .Y(n256) );
  OAI2BB2XL U1792 ( .B0(n2125), .B1(n2248), .A0N(\register[5][21] ), .A1N(
        n2248), .Y(n257) );
  OAI2BB2XL U1793 ( .B0(n2123), .B1(n2248), .A0N(\register[5][22] ), .A1N(
        n2249), .Y(n258) );
  OAI2BB2XL U1794 ( .B0(n2119), .B1(n2248), .A0N(\register[5][24] ), .A1N(
        n2249), .Y(n260) );
  OAI2BB2XL U1795 ( .B0(n2168), .B1(n2245), .A0N(\register[6][0] ), .A1N(n2245), .Y(n268) );
  OAI2BB2XL U1796 ( .B0(n2165), .B1(n2244), .A0N(\register[6][1] ), .A1N(n2244), .Y(n269) );
  OAI2BB2XL U1797 ( .B0(n2163), .B1(n2244), .A0N(\register[6][2] ), .A1N(n2245), .Y(n270) );
  OAI2BB2XL U1798 ( .B0(n2161), .B1(n2244), .A0N(\register[6][3] ), .A1N(n2246), .Y(n271) );
  OAI2BB2XL U1799 ( .B0(n2159), .B1(n2244), .A0N(\register[6][4] ), .A1N(n2244), .Y(n272) );
  OAI2BB2XL U1800 ( .B0(n2158), .B1(n2244), .A0N(\register[6][5] ), .A1N(n2246), .Y(n273) );
  OAI2BB2XL U1801 ( .B0(n2155), .B1(n2244), .A0N(\register[6][6] ), .A1N(n2246), .Y(n274) );
  OAI2BB2XL U1802 ( .B0(n2154), .B1(n2244), .A0N(\register[6][7] ), .A1N(n2246), .Y(n275) );
  OAI2BB2XL U1803 ( .B0(n2152), .B1(n2244), .A0N(\register[6][8] ), .A1N(n2246), .Y(n276) );
  OAI2BB2XL U1804 ( .B0(n2150), .B1(n2244), .A0N(\register[6][9] ), .A1N(n2246), .Y(n277) );
  OAI2BB2XL U1805 ( .B0(n2148), .B1(n2244), .A0N(\register[6][10] ), .A1N(
        n2246), .Y(n278) );
  OAI2BB2XL U1806 ( .B0(n2145), .B1(n2244), .A0N(\register[6][11] ), .A1N(
        n2246), .Y(n279) );
  OAI2BB2XL U1807 ( .B0(n2143), .B1(n2244), .A0N(\register[6][12] ), .A1N(
        n2246), .Y(n280) );
  OAI2BB2XL U1808 ( .B0(n2141), .B1(n2245), .A0N(\register[6][13] ), .A1N(
        n2246), .Y(n281) );
  OAI2BB2XL U1809 ( .B0(n2139), .B1(n2245), .A0N(\register[6][14] ), .A1N(
        n2246), .Y(n282) );
  OAI2BB2XL U1810 ( .B0(n2137), .B1(n2245), .A0N(\register[6][15] ), .A1N(
        n2246), .Y(n283) );
  OAI2BB2XL U1811 ( .B0(n2135), .B1(n2245), .A0N(\register[6][16] ), .A1N(
        n2246), .Y(n284) );
  OAI2BB2XL U1812 ( .B0(n2133), .B1(n2245), .A0N(\register[6][17] ), .A1N(
        n2244), .Y(n285) );
  OAI2BB2XL U1813 ( .B0(n2131), .B1(n2245), .A0N(\register[6][18] ), .A1N(
        n2245), .Y(n286) );
  OAI2BB2XL U1814 ( .B0(n2129), .B1(n2245), .A0N(\register[6][19] ), .A1N(
        n2246), .Y(n287) );
  OAI2BB2XL U1815 ( .B0(n2127), .B1(n2245), .A0N(\register[6][20] ), .A1N(
        n2244), .Y(n288) );
  OAI2BB2XL U1816 ( .B0(n2125), .B1(n2245), .A0N(\register[6][21] ), .A1N(
        n2245), .Y(n289) );
  OAI2BB2XL U1817 ( .B0(n2123), .B1(n2245), .A0N(\register[6][22] ), .A1N(
        n2246), .Y(n290) );
  OAI2BB2XL U1818 ( .B0(n2119), .B1(n2245), .A0N(\register[6][24] ), .A1N(
        n2246), .Y(n292) );
  OAI2BB2XL U1819 ( .B0(n2168), .B1(n2242), .A0N(\register[7][0] ), .A1N(n2242), .Y(n300) );
  OAI2BB2XL U1820 ( .B0(n2165), .B1(n2241), .A0N(\register[7][1] ), .A1N(n2241), .Y(n301) );
  OAI2BB2XL U1821 ( .B0(n2163), .B1(n2241), .A0N(\register[7][2] ), .A1N(n2242), .Y(n302) );
  OAI2BB2XL U1822 ( .B0(n2161), .B1(n2241), .A0N(\register[7][3] ), .A1N(n2243), .Y(n303) );
  OAI2BB2XL U1823 ( .B0(n2159), .B1(n2241), .A0N(\register[7][4] ), .A1N(n2241), .Y(n304) );
  OAI2BB2XL U1824 ( .B0(n2158), .B1(n2241), .A0N(\register[7][5] ), .A1N(n2243), .Y(n305) );
  OAI2BB2XL U1825 ( .B0(n2155), .B1(n2241), .A0N(\register[7][6] ), .A1N(n2243), .Y(n306) );
  OAI2BB2XL U1826 ( .B0(n2154), .B1(n2241), .A0N(\register[7][7] ), .A1N(n2243), .Y(n307) );
  OAI2BB2XL U1827 ( .B0(n2152), .B1(n2241), .A0N(\register[7][8] ), .A1N(n2243), .Y(n308) );
  OAI2BB2XL U1828 ( .B0(n2150), .B1(n2241), .A0N(\register[7][9] ), .A1N(n2243), .Y(n309) );
  OAI2BB2XL U1829 ( .B0(n2148), .B1(n2241), .A0N(\register[7][10] ), .A1N(
        n2243), .Y(n310) );
  OAI2BB2XL U1830 ( .B0(n2145), .B1(n2241), .A0N(\register[7][11] ), .A1N(
        n2243), .Y(n311) );
  OAI2BB2XL U1831 ( .B0(n2143), .B1(n2241), .A0N(\register[7][12] ), .A1N(
        n2243), .Y(n312) );
  OAI2BB2XL U1832 ( .B0(n2141), .B1(n2242), .A0N(\register[7][13] ), .A1N(
        n2243), .Y(n313) );
  OAI2BB2XL U1833 ( .B0(n2139), .B1(n2242), .A0N(\register[7][14] ), .A1N(
        n2243), .Y(n314) );
  OAI2BB2XL U1834 ( .B0(n2137), .B1(n2242), .A0N(\register[7][15] ), .A1N(
        n2243), .Y(n315) );
  OAI2BB2XL U1835 ( .B0(n2135), .B1(n2242), .A0N(\register[7][16] ), .A1N(
        n2243), .Y(n316) );
  OAI2BB2XL U1836 ( .B0(n2133), .B1(n2242), .A0N(\register[7][17] ), .A1N(
        n2241), .Y(n317) );
  OAI2BB2XL U1837 ( .B0(n2131), .B1(n2242), .A0N(\register[7][18] ), .A1N(
        n2242), .Y(n318) );
  OAI2BB2XL U1838 ( .B0(n2129), .B1(n2242), .A0N(\register[7][19] ), .A1N(
        n2243), .Y(n319) );
  OAI2BB2XL U1839 ( .B0(n2127), .B1(n2242), .A0N(\register[7][20] ), .A1N(
        n2241), .Y(n320) );
  OAI2BB2XL U1840 ( .B0(n2125), .B1(n2242), .A0N(\register[7][21] ), .A1N(
        n2242), .Y(n321) );
  OAI2BB2XL U1841 ( .B0(n2123), .B1(n2242), .A0N(\register[7][22] ), .A1N(
        n2243), .Y(n322) );
  OAI2BB2XL U1842 ( .B0(n2119), .B1(n2242), .A0N(\register[7][24] ), .A1N(
        n2243), .Y(n324) );
  NOR2BX1 U1843 ( .AN(N18), .B(\register[3][0] ), .Y(n2056) );
  NOR2BX1 U1844 ( .AN(n2074), .B(\register[3][1] ), .Y(n2051) );
  NOR2BX1 U1845 ( .AN(n2080), .B(\register[3][2] ), .Y(n2046) );
  NOR2BX1 U1846 ( .AN(n2080), .B(\register[3][3] ), .Y(n2041) );
  NOR2BX1 U1847 ( .AN(n2080), .B(\register[3][4] ), .Y(n2036) );
  NOR2BX1 U1848 ( .AN(n2079), .B(\register[3][5] ), .Y(n2031) );
  NOR2BX1 U1849 ( .AN(N18), .B(\register[3][6] ), .Y(n2026) );
  NOR2BX1 U1850 ( .AN(n2079), .B(\register[3][7] ), .Y(n2021) );
  NOR2BX1 U1851 ( .AN(n2079), .B(\register[3][8] ), .Y(n2016) );
  NOR2BX1 U1852 ( .AN(n2079), .B(\register[3][9] ), .Y(n2011) );
  NOR2BX1 U1853 ( .AN(n2079), .B(\register[3][10] ), .Y(n2006) );
  NOR2BX1 U1854 ( .AN(n2079), .B(\register[3][11] ), .Y(n2001) );
  NOR2BX1 U1855 ( .AN(N18), .B(\register[3][12] ), .Y(n1996) );
  NOR2BX1 U1856 ( .AN(n2079), .B(\register[3][13] ), .Y(n1991) );
  NOR2BX1 U1857 ( .AN(n2079), .B(\register[3][14] ), .Y(n1986) );
  NOR2BX1 U1858 ( .AN(n2079), .B(\register[3][15] ), .Y(n1981) );
  NOR2BX1 U1859 ( .AN(n2079), .B(\register[3][16] ), .Y(n1976) );
  NOR2BX1 U1860 ( .AN(n2079), .B(\register[3][17] ), .Y(n1971) );
  NOR2BX1 U1861 ( .AN(n2079), .B(\register[3][18] ), .Y(n1966) );
  NOR2BX1 U1862 ( .AN(n2079), .B(\register[3][19] ), .Y(n1961) );
  NOR2BX1 U1863 ( .AN(n2079), .B(\register[3][20] ), .Y(n1956) );
  NOR2BX1 U1864 ( .AN(n2079), .B(\register[3][21] ), .Y(n1951) );
  NOR2BX1 U1865 ( .AN(n2079), .B(\register[3][22] ), .Y(n1946) );
  NOR2BX1 U1866 ( .AN(n2079), .B(\register[3][23] ), .Y(n1941) );
  NOR2BX1 U1867 ( .AN(n2079), .B(\register[3][24] ), .Y(n1936) );
  NOR2BX1 U1868 ( .AN(n2083), .B(\register[3][25] ), .Y(n1931) );
  NOR2BX1 U1869 ( .AN(n2074), .B(\register[3][26] ), .Y(n1926) );
  NOR2BX1 U1870 ( .AN(N18), .B(\register[3][27] ), .Y(n1921) );
  NOR2BX1 U1871 ( .AN(N18), .B(\register[3][28] ), .Y(n1916) );
  NOR2BX1 U1872 ( .AN(N18), .B(\register[3][29] ), .Y(n1911) );
  NOR2BX1 U1873 ( .AN(N18), .B(\register[3][30] ), .Y(n1906) );
  NOR2BX1 U1874 ( .AN(n2074), .B(\register[3][31] ), .Y(n1901) );
  NOR2BX1 U1875 ( .AN(n1553), .B(\register[3][0] ), .Y(n1529) );
  NOR2BX1 U1876 ( .AN(n1553), .B(\register[3][1] ), .Y(n1524) );
  NOR2BX1 U1877 ( .AN(n1553), .B(\register[3][2] ), .Y(n1519) );
  NOR2BX1 U1878 ( .AN(n1553), .B(\register[3][3] ), .Y(n1514) );
  NOR2BX1 U1879 ( .AN(n1553), .B(\register[3][4] ), .Y(n1509) );
  NOR2BX1 U1880 ( .AN(n1552), .B(\register[3][5] ), .Y(n1504) );
  NOR2BX1 U1881 ( .AN(n1553), .B(\register[3][6] ), .Y(n1499) );
  NOR2BX1 U1882 ( .AN(n1552), .B(\register[3][7] ), .Y(n1494) );
  NOR2BX1 U1883 ( .AN(n1552), .B(\register[3][8] ), .Y(n1489) );
  NOR2BX1 U1884 ( .AN(n1552), .B(\register[3][9] ), .Y(n1484) );
  NOR2BX1 U1885 ( .AN(n1552), .B(\register[3][10] ), .Y(n1479) );
  NOR2BX1 U1886 ( .AN(n1552), .B(\register[3][11] ), .Y(n1474) );
  NOR2BX1 U1887 ( .AN(n1553), .B(\register[3][12] ), .Y(n1469) );
  NOR2BX1 U1888 ( .AN(n1552), .B(\register[3][13] ), .Y(n1464) );
  NOR2BX1 U1889 ( .AN(n1552), .B(\register[3][14] ), .Y(n1459) );
  NOR2BX1 U1890 ( .AN(n1552), .B(\register[3][15] ), .Y(n1454) );
  NOR2BX1 U1891 ( .AN(n1552), .B(\register[3][16] ), .Y(n1449) );
  NOR2BX1 U1892 ( .AN(n1552), .B(\register[3][17] ), .Y(n1444) );
  NOR2BX1 U1893 ( .AN(n1552), .B(\register[3][18] ), .Y(n1439) );
  NOR2BX1 U1894 ( .AN(n1552), .B(\register[3][19] ), .Y(n1434) );
  NOR2BX1 U1895 ( .AN(n1552), .B(\register[3][20] ), .Y(n1429) );
  NOR2BX1 U1896 ( .AN(n1552), .B(\register[3][21] ), .Y(n1424) );
  NOR2BX1 U1897 ( .AN(n1552), .B(\register[3][22] ), .Y(n1419) );
  NOR2BX1 U1898 ( .AN(n1552), .B(\register[3][23] ), .Y(n1414) );
  NOR2BX1 U1899 ( .AN(n1552), .B(\register[3][24] ), .Y(n1409) );
  NOR2BX1 U1900 ( .AN(n1553), .B(\register[3][25] ), .Y(n1404) );
  NOR2BX1 U1901 ( .AN(n1553), .B(\register[3][26] ), .Y(n1399) );
  NOR2BX1 U1902 ( .AN(n1553), .B(\register[3][27] ), .Y(n1394) );
  NOR2BX1 U1903 ( .AN(n1553), .B(\register[3][28] ), .Y(n1389) );
  NOR2BX1 U1904 ( .AN(n1553), .B(\register[3][29] ), .Y(n1384) );
  NOR2BX1 U1905 ( .AN(n1553), .B(\register[3][30] ), .Y(n1379) );
  NOR2BX1 U1906 ( .AN(n1553), .B(\register[3][31] ), .Y(n1374) );
  NOR2X1 U1907 ( .A(n1557), .B(\register[1][26] ), .Y(n1401) );
  NAND2X1 U1908 ( .A(n2055), .B(n2054), .Y(n1660) );
  NOR2X1 U1909 ( .A(n2053), .B(n2052), .Y(n2055) );
  MXI2X1 U1910 ( .A(n2387), .B(n2051), .S0(n2101), .Y(n2054) );
  NOR2X1 U1911 ( .A(n2081), .B(\register[1][1] ), .Y(n2053) );
  NAND2X1 U1912 ( .A(n1528), .B(n1527), .Y(n1133) );
  NOR2X1 U1913 ( .A(n1526), .B(n1525), .Y(n1528) );
  MXI2X1 U1914 ( .A(n2387), .B(n1524), .S0(n1576), .Y(n1527) );
  NOR2X1 U1915 ( .A(n1555), .B(\register[1][1] ), .Y(n1526) );
  NAND2X1 U1916 ( .A(n2050), .B(n2049), .Y(n1668) );
  NOR2X1 U1917 ( .A(n2048), .B(n2047), .Y(n2050) );
  MXI2X1 U1918 ( .A(n2388), .B(n2046), .S0(n2087), .Y(n2049) );
  NOR2X1 U1919 ( .A(n2081), .B(\register[1][2] ), .Y(n2048) );
  NAND2X1 U1920 ( .A(n2045), .B(n2044), .Y(n1676) );
  NOR2X1 U1921 ( .A(n2043), .B(n2042), .Y(n2045) );
  MXI2X1 U1922 ( .A(n2389), .B(n2041), .S0(n2088), .Y(n2044) );
  NOR2X1 U1923 ( .A(n2080), .B(\register[1][3] ), .Y(n2043) );
  NAND2X1 U1924 ( .A(n2040), .B(n2039), .Y(n1684) );
  NOR2X1 U1925 ( .A(n2038), .B(n2037), .Y(n2040) );
  MXI2X1 U1926 ( .A(n2390), .B(n2036), .S0(n2101), .Y(n2039) );
  NOR2X1 U1927 ( .A(N18), .B(\register[1][4] ), .Y(n2038) );
  NAND2X1 U1928 ( .A(n2035), .B(n2034), .Y(n1692) );
  NOR2X1 U1929 ( .A(n2033), .B(n2032), .Y(n2035) );
  MXI2X1 U1930 ( .A(n2391), .B(n2031), .S0(n2091), .Y(n2034) );
  NOR2X1 U1931 ( .A(n2080), .B(\register[1][5] ), .Y(n2033) );
  NAND2X1 U1932 ( .A(n2030), .B(n2029), .Y(n1700) );
  NOR2X1 U1933 ( .A(n2028), .B(n2027), .Y(n2030) );
  MXI2X1 U1934 ( .A(n2392), .B(n2026), .S0(n2092), .Y(n2029) );
  NOR2X1 U1935 ( .A(N18), .B(\register[1][6] ), .Y(n2028) );
  NAND2X1 U1936 ( .A(n2025), .B(n2024), .Y(n1708) );
  NOR2X1 U1937 ( .A(n2023), .B(n2022), .Y(n2025) );
  MXI2X1 U1938 ( .A(n2393), .B(n2021), .S0(n2084), .Y(n2024) );
  NOR2X1 U1939 ( .A(n2080), .B(\register[1][7] ), .Y(n2023) );
  NAND2X1 U1940 ( .A(n2020), .B(n2019), .Y(n1716) );
  NOR2X1 U1941 ( .A(n2018), .B(n2017), .Y(n2020) );
  MXI2X1 U1942 ( .A(n2394), .B(n2016), .S0(n2089), .Y(n2019) );
  NOR2X1 U1943 ( .A(n2081), .B(\register[1][8] ), .Y(n2018) );
  NAND2X1 U1944 ( .A(n2015), .B(n2014), .Y(n1724) );
  NOR2X1 U1945 ( .A(n2013), .B(n2012), .Y(n2015) );
  MXI2X1 U1946 ( .A(n2395), .B(n2011), .S0(n2090), .Y(n2014) );
  NOR2X1 U1947 ( .A(n2080), .B(\register[1][9] ), .Y(n2013) );
  NAND2X1 U1948 ( .A(n2010), .B(n2009), .Y(n1732) );
  NOR2X1 U1949 ( .A(n2008), .B(n2007), .Y(n2010) );
  MXI2X1 U1950 ( .A(n2396), .B(n2006), .S0(n2084), .Y(n2009) );
  NOR2X1 U1951 ( .A(n2080), .B(\register[1][10] ), .Y(n2008) );
  NAND2X1 U1952 ( .A(n2005), .B(n2004), .Y(n1740) );
  NOR2X1 U1953 ( .A(n2003), .B(n2002), .Y(n2005) );
  MXI2X1 U1954 ( .A(n2397), .B(n2001), .S0(n2084), .Y(n2004) );
  NOR2X1 U1955 ( .A(n2081), .B(\register[1][11] ), .Y(n2003) );
  NAND2X1 U1956 ( .A(n2000), .B(n1999), .Y(n1748) );
  NOR2X1 U1957 ( .A(n1998), .B(n1997), .Y(n2000) );
  MXI2X1 U1958 ( .A(n2398), .B(n1996), .S0(n2084), .Y(n1999) );
  NOR2X1 U1959 ( .A(n2081), .B(\register[1][12] ), .Y(n1998) );
  NAND2X1 U1960 ( .A(n1995), .B(n1994), .Y(n1756) );
  NOR2X1 U1961 ( .A(n1993), .B(n1992), .Y(n1995) );
  MXI2X1 U1962 ( .A(n2399), .B(n1991), .S0(n2084), .Y(n1994) );
  NOR2X1 U1963 ( .A(n2081), .B(\register[1][13] ), .Y(n1993) );
  NAND2X1 U1964 ( .A(n1990), .B(n1989), .Y(n1764) );
  NOR2X1 U1965 ( .A(n1988), .B(n1987), .Y(n1990) );
  MXI2X1 U1966 ( .A(n2400), .B(n1986), .S0(n2084), .Y(n1989) );
  NOR2X1 U1967 ( .A(n2081), .B(\register[1][14] ), .Y(n1988) );
  NAND2X1 U1968 ( .A(n1985), .B(n1984), .Y(n1772) );
  NOR2X1 U1969 ( .A(n1983), .B(n1982), .Y(n1985) );
  MXI2X1 U1970 ( .A(n2401), .B(n1981), .S0(n2102), .Y(n1984) );
  NOR2X1 U1971 ( .A(n2082), .B(\register[1][15] ), .Y(n1983) );
  NAND2X1 U1972 ( .A(n1980), .B(n1979), .Y(n1780) );
  NOR2X1 U1973 ( .A(n1978), .B(n1977), .Y(n1980) );
  MXI2X1 U1974 ( .A(n2402), .B(n1976), .S0(n2102), .Y(n1979) );
  NOR2X1 U1975 ( .A(n2082), .B(\register[1][16] ), .Y(n1978) );
  NAND2X1 U1976 ( .A(n1975), .B(n1974), .Y(n1788) );
  NOR2X1 U1977 ( .A(n1973), .B(n1972), .Y(n1975) );
  MXI2X1 U1978 ( .A(n2403), .B(n1971), .S0(n2102), .Y(n1974) );
  NOR2X1 U1979 ( .A(n2082), .B(\register[1][17] ), .Y(n1973) );
  NAND2X1 U1980 ( .A(n1970), .B(n1969), .Y(n1796) );
  NOR2X1 U1981 ( .A(n1968), .B(n1967), .Y(n1970) );
  MXI2X1 U1982 ( .A(n2404), .B(n1966), .S0(n2102), .Y(n1969) );
  NOR2X1 U1983 ( .A(n2082), .B(\register[1][18] ), .Y(n1968) );
  NAND2X1 U1984 ( .A(n1965), .B(n1964), .Y(n1804) );
  NOR2X1 U1985 ( .A(n1963), .B(n1962), .Y(n1965) );
  MXI2X1 U1986 ( .A(n2405), .B(n1961), .S0(n2102), .Y(n1964) );
  NOR2X1 U1987 ( .A(n2082), .B(\register[1][19] ), .Y(n1963) );
  NAND2X1 U1988 ( .A(n1960), .B(n1959), .Y(n1812) );
  NOR2X1 U1989 ( .A(n1958), .B(n1957), .Y(n1960) );
  MXI2X1 U1990 ( .A(n2406), .B(n1956), .S0(n2102), .Y(n1959) );
  NOR2X1 U1991 ( .A(n2082), .B(\register[1][20] ), .Y(n1958) );
  NAND2X1 U1992 ( .A(n1955), .B(n1954), .Y(n1820) );
  NOR2X1 U1993 ( .A(n1953), .B(n1952), .Y(n1955) );
  MXI2X1 U1994 ( .A(n2407), .B(n1951), .S0(n2102), .Y(n1954) );
  NOR2X1 U1995 ( .A(n2083), .B(\register[1][21] ), .Y(n1953) );
  NAND2X1 U1996 ( .A(n1950), .B(n1949), .Y(n1828) );
  NOR2X1 U1997 ( .A(n1948), .B(n1947), .Y(n1950) );
  MXI2X1 U1998 ( .A(n2408), .B(n1946), .S0(n2102), .Y(n1949) );
  NOR2X1 U1999 ( .A(n2083), .B(\register[1][22] ), .Y(n1948) );
  NAND2X1 U2000 ( .A(n1945), .B(n1944), .Y(n1836) );
  NOR2X1 U2001 ( .A(n1943), .B(n1942), .Y(n1945) );
  MXI2X1 U2002 ( .A(n2409), .B(n1941), .S0(n2102), .Y(n1944) );
  NOR2X1 U2003 ( .A(n2083), .B(\register[1][23] ), .Y(n1943) );
  NAND2X1 U2004 ( .A(n1940), .B(n1939), .Y(n1844) );
  NOR2X1 U2005 ( .A(n1938), .B(n1937), .Y(n1940) );
  MXI2X1 U2006 ( .A(n2410), .B(n1936), .S0(n2102), .Y(n1939) );
  NOR2X1 U2007 ( .A(n2083), .B(\register[1][24] ), .Y(n1938) );
  NAND2X1 U2008 ( .A(n1930), .B(n1929), .Y(n1860) );
  NOR2X1 U2009 ( .A(n1928), .B(n1927), .Y(n1930) );
  MXI2X1 U2010 ( .A(n2412), .B(n1926), .S0(n2102), .Y(n1929) );
  NOR2X1 U2011 ( .A(n2083), .B(\register[1][26] ), .Y(n1928) );
  NAND2X1 U2012 ( .A(n1915), .B(n1914), .Y(n1884) );
  NOR2X1 U2013 ( .A(n1913), .B(n1912), .Y(n1915) );
  MXI2X1 U2014 ( .A(n2415), .B(n1911), .S0(n2102), .Y(n1914) );
  NOR2X1 U2015 ( .A(N18), .B(\register[1][29] ), .Y(n1913) );
  NAND2X1 U2016 ( .A(n1905), .B(n1904), .Y(n1900) );
  NOR2X1 U2017 ( .A(n1903), .B(n1902), .Y(n1905) );
  MXI2X1 U2018 ( .A(n2417), .B(n1901), .S0(n2102), .Y(n1904) );
  NOR2X1 U2019 ( .A(n2081), .B(\register[1][31] ), .Y(n1903) );
  NAND2X1 U2020 ( .A(n1523), .B(n1522), .Y(n1141) );
  NOR2X1 U2021 ( .A(n1521), .B(n1520), .Y(n1523) );
  MXI2X1 U2022 ( .A(n2388), .B(n1519), .S0(n1562), .Y(n1522) );
  NOR2X1 U2023 ( .A(n1555), .B(\register[1][2] ), .Y(n1521) );
  NAND2X1 U2024 ( .A(n1518), .B(n1517), .Y(n1149) );
  NOR2X1 U2025 ( .A(n1516), .B(n1515), .Y(n1518) );
  MXI2X1 U2026 ( .A(n2389), .B(n1514), .S0(n1559), .Y(n1517) );
  NOR2X1 U2027 ( .A(n1554), .B(\register[1][3] ), .Y(n1516) );
  NAND2X1 U2028 ( .A(n1513), .B(n1512), .Y(n1157) );
  NOR2X1 U2029 ( .A(n1511), .B(n1510), .Y(n1513) );
  MXI2X1 U2030 ( .A(n2390), .B(n1509), .S0(n1559), .Y(n1512) );
  NOR2X1 U2031 ( .A(n1553), .B(\register[1][4] ), .Y(n1511) );
  NAND2X1 U2032 ( .A(n1508), .B(n1507), .Y(n1165) );
  NOR2X1 U2033 ( .A(n1506), .B(n1505), .Y(n1508) );
  MXI2X1 U2034 ( .A(n2391), .B(n1504), .S0(n1559), .Y(n1507) );
  NOR2X1 U2035 ( .A(n1554), .B(\register[1][5] ), .Y(n1506) );
  NAND2X1 U2036 ( .A(n1503), .B(n1502), .Y(n1173) );
  NOR2X1 U2037 ( .A(n1501), .B(n1500), .Y(n1503) );
  MXI2X1 U2038 ( .A(n2392), .B(n1499), .S0(n1559), .Y(n1502) );
  NOR2X1 U2039 ( .A(n1553), .B(\register[1][6] ), .Y(n1501) );
  NAND2X1 U2040 ( .A(n1498), .B(n1497), .Y(n1181) );
  NOR2X1 U2041 ( .A(n1496), .B(n1495), .Y(n1498) );
  MXI2X1 U2042 ( .A(n2393), .B(n1494), .S0(n1559), .Y(n1497) );
  NOR2X1 U2043 ( .A(n1554), .B(\register[1][7] ), .Y(n1496) );
  NAND2X1 U2044 ( .A(n1493), .B(n1492), .Y(n1189) );
  NOR2X1 U2045 ( .A(n1491), .B(n1490), .Y(n1493) );
  MXI2X1 U2046 ( .A(n2394), .B(n1489), .S0(n1559), .Y(n1492) );
  NOR2X1 U2047 ( .A(n1555), .B(\register[1][8] ), .Y(n1491) );
  NAND2X1 U2048 ( .A(n1488), .B(n1487), .Y(n1197) );
  NOR2X1 U2049 ( .A(n1486), .B(n1485), .Y(n1488) );
  MXI2X1 U2050 ( .A(n2395), .B(n1484), .S0(n1563), .Y(n1487) );
  NOR2X1 U2051 ( .A(n1554), .B(\register[1][9] ), .Y(n1486) );
  NAND2X1 U2052 ( .A(n1483), .B(n1482), .Y(n1205) );
  NOR2X1 U2053 ( .A(n1481), .B(n1480), .Y(n1483) );
  MXI2X1 U2054 ( .A(n2396), .B(n1479), .S0(n1567), .Y(n1482) );
  NOR2X1 U2055 ( .A(n1554), .B(\register[1][10] ), .Y(n1481) );
  NAND2X1 U2056 ( .A(n1478), .B(n1477), .Y(n1213) );
  NOR2X1 U2057 ( .A(n1476), .B(n1475), .Y(n1478) );
  MXI2X1 U2058 ( .A(n2397), .B(n1474), .S0(n1565), .Y(n1477) );
  NOR2X1 U2059 ( .A(n1555), .B(\register[1][11] ), .Y(n1476) );
  NAND2X1 U2060 ( .A(n1473), .B(n1472), .Y(n1221) );
  NOR2X1 U2061 ( .A(n1471), .B(n1470), .Y(n1473) );
  MXI2X1 U2062 ( .A(n2398), .B(n1469), .S0(n1564), .Y(n1472) );
  NOR2X1 U2063 ( .A(n1555), .B(\register[1][12] ), .Y(n1471) );
  NAND2X1 U2064 ( .A(n1468), .B(n1467), .Y(n1229) );
  NOR2X1 U2065 ( .A(n1466), .B(n1465), .Y(n1468) );
  MXI2X1 U2066 ( .A(n2399), .B(n1464), .S0(n1566), .Y(n1467) );
  NOR2X1 U2067 ( .A(n1555), .B(\register[1][13] ), .Y(n1466) );
  NAND2X1 U2068 ( .A(n1463), .B(n1462), .Y(n1237) );
  NOR2X1 U2069 ( .A(n1461), .B(n1460), .Y(n1463) );
  MXI2X1 U2070 ( .A(n2400), .B(n1459), .S0(n1576), .Y(n1462) );
  NOR2X1 U2071 ( .A(n1555), .B(\register[1][14] ), .Y(n1461) );
  NAND2X1 U2072 ( .A(n1458), .B(n1457), .Y(n1245) );
  NOR2X1 U2073 ( .A(n1456), .B(n1455), .Y(n1458) );
  MXI2X1 U2074 ( .A(n2401), .B(n1454), .S0(n1577), .Y(n1457) );
  NOR2X1 U2075 ( .A(n1556), .B(\register[1][15] ), .Y(n1456) );
  NAND2X1 U2076 ( .A(n1453), .B(n1452), .Y(n1253) );
  NOR2X1 U2077 ( .A(n1451), .B(n1450), .Y(n1453) );
  MXI2X1 U2078 ( .A(n2402), .B(n1449), .S0(n1577), .Y(n1452) );
  NOR2X1 U2079 ( .A(n1556), .B(\register[1][16] ), .Y(n1451) );
  NAND2X1 U2080 ( .A(n1448), .B(n1447), .Y(n1261) );
  NOR2X1 U2081 ( .A(n1446), .B(n1445), .Y(n1448) );
  MXI2X1 U2082 ( .A(n2403), .B(n1444), .S0(n1577), .Y(n1447) );
  NOR2X1 U2083 ( .A(n1556), .B(\register[1][17] ), .Y(n1446) );
  NAND2X1 U2084 ( .A(n1443), .B(n1442), .Y(n1269) );
  NOR2X1 U2085 ( .A(n1441), .B(n1440), .Y(n1443) );
  MXI2X1 U2086 ( .A(n2404), .B(n1439), .S0(n1577), .Y(n1442) );
  NOR2X1 U2087 ( .A(n1556), .B(\register[1][18] ), .Y(n1441) );
  NAND2X1 U2088 ( .A(n1438), .B(n1437), .Y(n1277) );
  NOR2X1 U2089 ( .A(n1436), .B(n1435), .Y(n1438) );
  MXI2X1 U2090 ( .A(n2405), .B(n1434), .S0(n1577), .Y(n1437) );
  NOR2X1 U2091 ( .A(n1556), .B(\register[1][19] ), .Y(n1436) );
  NAND2X1 U2092 ( .A(n1433), .B(n1432), .Y(n1285) );
  NOR2X1 U2093 ( .A(n1431), .B(n1430), .Y(n1433) );
  MXI2X1 U2094 ( .A(n2406), .B(n1429), .S0(n1577), .Y(n1432) );
  NOR2X1 U2095 ( .A(n1556), .B(\register[1][20] ), .Y(n1431) );
  NAND2X1 U2096 ( .A(n1428), .B(n1427), .Y(n1293) );
  NOR2X1 U2097 ( .A(n1426), .B(n1425), .Y(n1428) );
  MXI2X1 U2098 ( .A(n2407), .B(n1424), .S0(n1577), .Y(n1427) );
  NOR2X1 U2099 ( .A(n1557), .B(\register[1][21] ), .Y(n1426) );
  NAND2X1 U2100 ( .A(n1423), .B(n1422), .Y(n1301) );
  NOR2X1 U2101 ( .A(n1421), .B(n1420), .Y(n1423) );
  MXI2X1 U2102 ( .A(n2408), .B(n1419), .S0(n1577), .Y(n1422) );
  NOR2X1 U2103 ( .A(n1557), .B(\register[1][22] ), .Y(n1421) );
  NAND2X1 U2104 ( .A(n1418), .B(n1417), .Y(n1309) );
  NOR2X1 U2105 ( .A(n1416), .B(n1415), .Y(n1418) );
  MXI2X1 U2106 ( .A(n2409), .B(n1414), .S0(n1577), .Y(n1417) );
  NOR2X1 U2107 ( .A(n1557), .B(\register[1][23] ), .Y(n1416) );
  NAND2X1 U2108 ( .A(n1413), .B(n1412), .Y(n1317) );
  NOR2X1 U2109 ( .A(n1411), .B(n1410), .Y(n1413) );
  MXI2X1 U2110 ( .A(n2410), .B(n1409), .S0(n1577), .Y(n1412) );
  NOR2X1 U2111 ( .A(n1557), .B(\register[1][24] ), .Y(n1411) );
  NAND2X1 U2112 ( .A(n1403), .B(n1402), .Y(n1333) );
  NOR2X1 U2113 ( .A(n1401), .B(n1400), .Y(n1403) );
  MXI2X1 U2114 ( .A(n2412), .B(n1399), .S0(n1577), .Y(n1402) );
  NOR2X1 U2115 ( .A(n1558), .B(n1579), .Y(n1400) );
  NAND2X1 U2116 ( .A(n1388), .B(n1387), .Y(n1357) );
  NOR2X1 U2117 ( .A(n1386), .B(n1385), .Y(n1388) );
  MXI2X1 U2118 ( .A(n2415), .B(n1384), .S0(n1577), .Y(n1387) );
  NOR2X1 U2119 ( .A(n1558), .B(\register[1][29] ), .Y(n1386) );
  NAND2X1 U2120 ( .A(n1378), .B(n1377), .Y(n1373) );
  NOR2X1 U2121 ( .A(n1376), .B(n1375), .Y(n1378) );
  MXI2X1 U2122 ( .A(n2417), .B(n1374), .S0(n1577), .Y(n1377) );
  NOR2X1 U2123 ( .A(n1558), .B(\register[1][31] ), .Y(n1376) );
  NAND2X1 U2124 ( .A(n2060), .B(n2059), .Y(n1652) );
  NOR2X1 U2125 ( .A(n2058), .B(n2057), .Y(n2060) );
  MXI2X1 U2126 ( .A(n2386), .B(n2056), .S0(n2085), .Y(n2059) );
  NOR2X1 U2127 ( .A(n2082), .B(\register[1][0] ), .Y(n2058) );
  NAND2X1 U2128 ( .A(n1935), .B(n1934), .Y(n1852) );
  NOR2X1 U2129 ( .A(n1933), .B(n1932), .Y(n1935) );
  MXI2X1 U2130 ( .A(n2411), .B(n1931), .S0(n2268), .Y(n1934) );
  NOR2X1 U2131 ( .A(n2083), .B(\register[1][25] ), .Y(n1933) );
  NAND2X1 U2132 ( .A(n1925), .B(n1924), .Y(n1868) );
  NOR2X1 U2133 ( .A(n1923), .B(n1922), .Y(n1925) );
  MXI2X1 U2134 ( .A(n2413), .B(n1921), .S0(n2093), .Y(n1924) );
  NOR2X1 U2135 ( .A(n2083), .B(\register[1][27] ), .Y(n1923) );
  NAND2X1 U2136 ( .A(n1920), .B(n1919), .Y(n1876) );
  NOR2X1 U2137 ( .A(n1918), .B(n1917), .Y(n1920) );
  MXI2X1 U2138 ( .A(n2414), .B(n1916), .S0(n2096), .Y(n1919) );
  NOR2X1 U2139 ( .A(n2081), .B(\register[1][28] ), .Y(n1918) );
  NAND2X1 U2140 ( .A(n1910), .B(n1909), .Y(n1892) );
  NOR2X1 U2141 ( .A(n1908), .B(n1907), .Y(n1910) );
  MXI2X1 U2142 ( .A(n2416), .B(n1906), .S0(n2094), .Y(n1909) );
  NOR2X1 U2143 ( .A(n2081), .B(\register[1][30] ), .Y(n1908) );
  NAND2X1 U2144 ( .A(n1533), .B(n1532), .Y(n1125) );
  NOR2X1 U2145 ( .A(n1531), .B(n1530), .Y(n1533) );
  MXI2X1 U2146 ( .A(n2386), .B(n1529), .S0(n1578), .Y(n1532) );
  NOR2X1 U2147 ( .A(n1558), .B(\register[1][0] ), .Y(n1531) );
  NAND2X1 U2148 ( .A(n1408), .B(n1407), .Y(n1325) );
  NOR2X1 U2149 ( .A(n1406), .B(n1405), .Y(n1408) );
  MXI2X1 U2150 ( .A(n2411), .B(n1404), .S0(n1578), .Y(n1407) );
  NOR2X1 U2151 ( .A(n1557), .B(\register[1][25] ), .Y(n1406) );
  NAND2X1 U2152 ( .A(n1398), .B(n1397), .Y(n1341) );
  NOR2X1 U2153 ( .A(n1396), .B(n1395), .Y(n1398) );
  MXI2X1 U2154 ( .A(n2413), .B(n1394), .S0(n1578), .Y(n1397) );
  NOR2X1 U2155 ( .A(n1558), .B(\register[1][27] ), .Y(n1396) );
  NAND2X1 U2156 ( .A(n1393), .B(n1392), .Y(n1349) );
  NOR2X1 U2157 ( .A(n1391), .B(n1390), .Y(n1393) );
  MXI2X1 U2158 ( .A(n2414), .B(n1389), .S0(n1578), .Y(n1392) );
  NOR2X1 U2159 ( .A(n1558), .B(\register[1][28] ), .Y(n1391) );
  NAND2X1 U2160 ( .A(n1383), .B(n1382), .Y(n1365) );
  NOR2X1 U2161 ( .A(n1381), .B(n1380), .Y(n1383) );
  MXI2X1 U2162 ( .A(n2416), .B(n1379), .S0(n1578), .Y(n1382) );
  NOR2X1 U2163 ( .A(n1558), .B(\register[1][30] ), .Y(n1381) );
  MXI4X1 U2164 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n2094), .S1(n2075), .Y(
        n1651) );
  MXI4X1 U2165 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n2094), .S1(n2075), .Y(
        n1647) );
  MXI4X1 U2166 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n2095), .S1(n2075), .Y(
        n1655) );
  MXI4X1 U2167 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n2095), .S1(n2075), .Y(
        n1659) );
  MXI4X1 U2168 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n2095), .S1(n2075), .Y(
        n1663) );
  MXI4X1 U2169 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n2095), .S1(n2075), .Y(
        n1667) );
  MXI4X1 U2170 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n2095), .S1(n2076), .Y(
        n1671) );
  MXI4X1 U2171 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n2096), .S1(n2076), .Y(
        n1675) );
  MXI4X1 U2172 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n2096), .S1(n2076), .Y(
        n1679) );
  MXI4X1 U2173 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n2096), .S1(n2076), .Y(
        n1683) );
  MXI4X1 U2174 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n2096), .S1(n2076), .Y(
        n1687) );
  MXI4X1 U2175 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n2097), .S1(n2076), .Y(
        n1691) );
  MXI4X1 U2176 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n2097), .S1(n2077), .Y(
        n1695) );
  MXI4X1 U2177 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n2097), .S1(n2077), .Y(
        n1699) );
  MXI4X1 U2178 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n2097), .S1(n2077), .Y(
        n1703) );
  MXI4X1 U2179 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n2098), .S1(n2077), .Y(
        n1707) );
  MXI4X1 U2180 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n2098), .S1(n2077), .Y(
        n1711) );
  MXI4X1 U2181 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n2098), .S1(n2077), .Y(
        n1715) );
  MXI4X1 U2182 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n2098), .S1(n2080), .Y(
        n1719) );
  MXI4X1 U2183 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n2099), .S1(n2080), .Y(
        n1723) );
  MXI4X1 U2184 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n2099), .S1(n2076), 
        .Y(n1727) );
  MXI4X1 U2185 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n2099), .S1(n2080), .Y(
        n1731) );
  MXI4X1 U2186 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n2099), .S1(n2081), 
        .Y(n1735) );
  MXI4X1 U2187 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n2100), .S1(n2081), .Y(
        n1739) );
  MXI4X1 U2188 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n2100), .S1(n2078), 
        .Y(n1743) );
  MXI4X1 U2189 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n2098), .S1(n2077), .Y(
        n1747) );
  MXI4X1 U2190 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1751) );
  MXI4X1 U2191 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n2100), .S1(n2078), .Y(
        n1755) );
  MXI4X1 U2192 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n2101), .S1(n2078), 
        .Y(n1759) );
  MXI4X1 U2193 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n2101), .S1(n2078), .Y(
        n1763) );
  MXI4X1 U2194 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n2101), .S1(n2078), 
        .Y(n1767) );
  MXI4X1 U2195 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n2098), .S1(n2077), .Y(
        n1771) );
  MXI4X1 U2196 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n2087), .S1(n2070), .Y(
        n1779) );
  MXI4X1 U2197 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1775) );
  MXI4X1 U2198 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n2087), .S1(n2070), .Y(
        n1787) );
  MXI4X1 U2199 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1783) );
  MXI4X1 U2200 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n2088), .S1(n2070), .Y(
        n1795) );
  MXI4X1 U2201 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n2088), .S1(n2070), 
        .Y(n1791) );
  MXI4X1 U2202 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n2088), .S1(n2071), .Y(
        n1803) );
  MXI4X1 U2203 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n2088), .S1(n2071), 
        .Y(n1799) );
  MXI4X1 U2204 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n2089), .S1(n2071), .Y(
        n1811) );
  MXI4X1 U2205 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n2089), .S1(n2071), 
        .Y(n1807) );
  MXI4X1 U2206 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n2089), .S1(n2071), .Y(
        n1819) );
  MXI4X1 U2207 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1815) );
  MXI4X1 U2208 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n2090), .S1(n2072), .Y(
        n1827) );
  MXI4X1 U2209 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n2089), .S1(n2072), 
        .Y(n1823) );
  MXI4X1 U2210 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n2090), .S1(n2072), .Y(
        n1835) );
  MXI4X1 U2211 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1831) );
  MXI4X1 U2212 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n2091), .S1(n2072), .Y(
        n1843) );
  MXI4X1 U2213 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n2090), .S1(n2072), 
        .Y(n1839) );
  MXI4X1 U2214 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n2091), .S1(n2073), .Y(
        n1851) );
  MXI4X1 U2215 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n2091), .S1(n2073), 
        .Y(n1847) );
  MXI4X1 U2216 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n2092), .S1(n2073), .Y(
        n1859) );
  MXI4X1 U2217 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n2091), .S1(n2073), 
        .Y(n1855) );
  MXI4X1 U2218 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n2092), .S1(n2073), .Y(
        n1867) );
  MXI4X1 U2219 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1863) );
  MXI4X1 U2220 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n2093), .S1(n2074), .Y(
        n1875) );
  MXI4X1 U2221 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n2092), .S1(n2073), 
        .Y(n1871) );
  MXI4X1 U2222 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n2093), .S1(n2074), .Y(
        n1883) );
  MXI4X1 U2223 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1879) );
  MXI4X1 U2224 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n2094), .S1(n2074), .Y(
        n1891) );
  MXI4X1 U2225 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1887) );
  MXI4X1 U2226 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n2101), .S1(n2079), .Y(
        n1899) );
  MXI4X1 U2227 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n2094), .S1(n2074), 
        .Y(n1895) );
  MXI4X1 U2228 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n1569), .S1(n1550), .Y(
        n1124) );
  MXI4X1 U2229 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1569), .S1(n1550), .Y(
        n1120) );
  MXI4X1 U2230 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1570), .S1(n1550), .Y(
        n1128) );
  MXI4X1 U2231 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n1570), .S1(n1550), .Y(
        n1132) );
  MXI4X1 U2232 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1570), .S1(n1550), .Y(
        n1136) );
  MXI4X1 U2233 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n1570), .S1(n1550), .Y(
        n1140) );
  MXI4X1 U2234 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1570), .S1(n1551), .Y(
        n1144) );
  MXI4X1 U2235 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n1571), .S1(n1551), .Y(
        n1148) );
  MXI4X1 U2236 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1571), .S1(n1551), .Y(
        n1152) );
  MXI4X1 U2237 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n1571), .S1(n1551), .Y(
        n1156) );
  MXI4X1 U2238 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1571), .S1(n1551), .Y(
        n1160) );
  MXI4X1 U2239 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n1572), .S1(n1551), .Y(
        n1164) );
  MXI4X1 U2240 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1572), .S1(n1545), .Y(
        n1168) );
  MXI4X1 U2241 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n1572), .S1(n1554), .Y(
        n1172) );
  MXI4X1 U2242 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1572), .S1(n1544), .Y(
        n1176) );
  MXI4X1 U2243 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1573), .S1(n1545), .Y(
        n1180) );
  MXI4X1 U2244 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1573), .S1(n1544), .Y(
        n1184) );
  MXI4X1 U2245 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1573), .S1(n1555), .Y(
        n1188) );
  MXI4X1 U2246 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1573), .S1(n1547), .Y(
        n1192) );
  MXI4X1 U2247 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1574), .S1(n1553), .Y(
        n1196) );
  MXI4X1 U2248 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1574), .S1(n1546), 
        .Y(n1200) );
  MXI4X1 U2249 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1574), .S1(n1558), .Y(
        n1204) );
  MXI4X1 U2250 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1574), .S1(n1548), 
        .Y(n1208) );
  MXI4X1 U2251 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1575), .S1(n1547), .Y(
        n1212) );
  MXI4X1 U2252 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1575), .S1(n1551), 
        .Y(n1216) );
  MXI4X1 U2253 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1573), .S1(n1545), .Y(
        n1220) );
  MXI4X1 U2254 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1575), .S1(n1550), 
        .Y(n1224) );
  MXI4X1 U2255 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1575), .S1(n1548), .Y(
        n1228) );
  MXI4X1 U2256 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1576), .S1(n1557), 
        .Y(n1232) );
  MXI4X1 U2257 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1576), .S1(n1549), .Y(
        n1236) );
  MXI4X1 U2258 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1576), .S1(n1551), 
        .Y(n1240) );
  MXI4X1 U2259 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1573), .S1(n1545), .Y(
        n1244) );
  MXI4X1 U2260 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1562), .S1(n1546), .Y(
        n1252) );
  MXI4X1 U2261 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1248) );
  MXI4X1 U2262 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1562), .S1(n1546), .Y(
        n1260) );
  MXI4X1 U2263 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1256) );
  MXI4X1 U2264 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1563), .S1(n1546), .Y(
        n1268) );
  MXI4X1 U2265 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1563), .S1(n1546), 
        .Y(n1264) );
  MXI4X1 U2266 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1563), .S1(n1558), .Y(
        n1276) );
  MXI4X1 U2267 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1563), .S1(n1547), 
        .Y(n1272) );
  MXI4X1 U2268 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1564), .S1(n1554), .Y(
        n1284) );
  MXI4X1 U2269 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1564), .S1(n1548), 
        .Y(n1280) );
  MXI4X1 U2270 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1564), .S1(n1554), .Y(
        n1292) );
  MXI4X1 U2271 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1564), .S1(n1557), 
        .Y(n1288) );
  MXI4X1 U2272 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1565), .S1(n1547), .Y(
        n1300) );
  MXI4X1 U2273 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1564), .S1(n1547), 
        .Y(n1296) );
  MXI4X1 U2274 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1565), .S1(n1547), .Y(
        n1308) );
  MXI4X1 U2275 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1304) );
  MXI4X1 U2276 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1566), .S1(n1547), .Y(
        n1316) );
  MXI4X1 U2277 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1565), .S1(n1547), 
        .Y(n1312) );
  MXI4X1 U2278 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1566), .S1(n1548), .Y(
        n1324) );
  MXI4X1 U2279 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1566), .S1(n1548), 
        .Y(n1320) );
  MXI4X1 U2280 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1567), .S1(n1548), .Y(
        n1332) );
  MXI4X1 U2281 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1566), .S1(n1548), 
        .Y(n1328) );
  MXI4X1 U2282 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1567), .S1(n1548), .Y(
        n1340) );
  MXI4X1 U2283 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1336) );
  MXI4X1 U2284 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1568), .S1(n1549), .Y(
        n1348) );
  MXI4X1 U2285 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1567), .S1(n1548), 
        .Y(n1344) );
  MXI4X1 U2286 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1568), .S1(n1549), .Y(
        n1356) );
  MXI4X1 U2287 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1352) );
  MXI4X1 U2288 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1569), .S1(n1549), .Y(
        n1364) );
  MXI4X1 U2289 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1360) );
  MXI4X1 U2290 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1576), .S1(n1552), .Y(
        n1372) );
  MXI4X1 U2291 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1569), .S1(n1549), 
        .Y(n1368) );
  MXI4X1 U2292 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n2095), .S1(n2075), .Y(
        n1656) );
  MXI4X1 U2293 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n2095), .S1(n2075), .Y(
        n1664) );
  MXI4X1 U2294 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n2096), .S1(n2076), .Y(
        n1672) );
  MXI4X1 U2295 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n2096), .S1(n2076), .Y(
        n1680) );
  MXI4X1 U2296 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n2096), .S1(n2076), .Y(
        n1688) );
  MXI4X1 U2297 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n2097), .S1(n2077), .Y(
        n1696) );
  MXI4X1 U2298 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n2097), .S1(n2077), .Y(
        n1704) );
  MXI4X1 U2299 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n2098), .S1(n2077), .Y(
        n1712) );
  MXI4X1 U2300 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n2098), .S1(n2074), .Y(
        n1720) );
  MXI4X1 U2301 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n2099), .S1(n2072), 
        .Y(n1728) );
  MXI4X1 U2302 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n2099), .S1(n2074), 
        .Y(n1736) );
  MXI4X1 U2303 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n2100), .S1(n2078), 
        .Y(n1744) );
  MXI4X1 U2304 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1752) );
  MXI4X1 U2305 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n2101), .S1(n2078), 
        .Y(n1760) );
  MXI4X1 U2306 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n2101), .S1(n2078), 
        .Y(n1768) );
  MXI4X1 U2307 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1570), .S1(n1550), .Y(
        n1129) );
  MXI4X1 U2308 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1570), .S1(n1550), .Y(
        n1137) );
  MXI4X1 U2309 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1571), .S1(n1551), .Y(
        n1145) );
  MXI4X1 U2310 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1571), .S1(n1551), .Y(
        n1153) );
  MXI4X1 U2311 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1571), .S1(n1551), .Y(
        n1161) );
  MXI4X1 U2312 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1572), .S1(n1545), .Y(
        n1169) );
  MXI4X1 U2313 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1572), .S1(n1553), .Y(
        n1177) );
  MXI4X1 U2314 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1573), .S1(n1546), .Y(
        n1185) );
  MXI4X1 U2315 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1573), .S1(n1544), .Y(
        n1193) );
  MXI4X1 U2316 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1574), .S1(n1554), 
        .Y(n1201) );
  MXI4X1 U2317 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1574), .S1(n1545), 
        .Y(n1209) );
  MXI4X1 U2318 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1575), .S1(n1550), 
        .Y(n1217) );
  MXI4X1 U2319 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1575), .S1(n1548), 
        .Y(n1225) );
  MXI4X1 U2320 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1576), .S1(n1546), 
        .Y(n1233) );
  MXI4X1 U2321 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1576), .S1(n1550), 
        .Y(n1241) );
  MXI4X1 U2322 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n2094), .S1(n2075), .Y(
        n1649) );
  MXI4X1 U2323 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n2094), .S1(n2075), .Y(
        n1645) );
  MXI4X1 U2324 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n2094), .S1(n2075), .Y(
        n1653) );
  MXI4X1 U2325 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n2095), .S1(n2075), .Y(
        n1657) );
  MXI4X1 U2326 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n2095), .S1(n2075), .Y(
        n1661) );
  MXI4X1 U2327 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n2095), .S1(n2075), .Y(
        n1665) );
  MXI4X1 U2328 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n2095), .S1(n2076), .Y(
        n1669) );
  MXI4X1 U2329 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n2096), .S1(n2076), .Y(
        n1673) );
  MXI4X1 U2330 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n2096), .S1(n2076), .Y(
        n1677) );
  MXI4X1 U2331 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n2096), .S1(n2076), .Y(
        n1681) );
  MXI4X1 U2332 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n2096), .S1(n2076), .Y(
        n1685) );
  MXI4X1 U2333 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n2097), .S1(n2076), .Y(
        n1689) );
  MXI4X1 U2334 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n2097), .S1(n2076), .Y(
        n1693) );
  MXI4X1 U2335 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n2097), .S1(n2077), .Y(
        n1697) );
  MXI4X1 U2336 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n2097), .S1(n2077), .Y(
        n1701) );
  MXI4X1 U2337 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n2097), .S1(n2077), .Y(
        n1705) );
  MXI4X1 U2338 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n2101), .S1(n2079), .Y(
        n1709) );
  MXI4X1 U2339 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n2098), .S1(n2077), .Y(
        n1713) );
  MXI4X1 U2340 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n2098), .S1(n2077), .Y(
        n1717) );
  MXI4X1 U2341 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n2098), .S1(n2082), .Y(
        n1721) );
  MXI4X1 U2342 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n2099), .S1(n2071), 
        .Y(n1725) );
  MXI4X1 U2343 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n2099), .S1(n2078), 
        .Y(n1729) );
  MXI4X1 U2344 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n2099), .S1(n2070), 
        .Y(n1733) );
  MXI4X1 U2345 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n2099), .S1(n2075), 
        .Y(n1737) );
  MXI4X1 U2346 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n2100), .S1(n2077), 
        .Y(n1741) );
  MXI4X1 U2347 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n2100), .S1(n2078), 
        .Y(n1745) );
  MXI4X1 U2348 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1749) );
  MXI4X1 U2349 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1753) );
  MXI4X1 U2350 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n2100), .S1(n2078), 
        .Y(n1757) );
  MXI4X1 U2351 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n2101), .S1(n2078), 
        .Y(n1761) );
  MXI4X1 U2352 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n2101), .S1(n2078), 
        .Y(n1765) );
  MXI4X1 U2353 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n2101), .S1(n2079), 
        .Y(n1769) );
  MXI4X1 U2354 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1777) );
  MXI4X1 U2355 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1773) );
  MXI4X1 U2356 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1785) );
  MXI4X1 U2357 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1781) );
  MXI4X1 U2358 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n2088), .S1(n2070), 
        .Y(n1793) );
  MXI4X1 U2359 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n2087), .S1(n2070), 
        .Y(n1789) );
  MXI4X1 U2360 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n2088), .S1(n2071), 
        .Y(n1801) );
  MXI4X1 U2361 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n2088), .S1(n2070), 
        .Y(n1797) );
  MXI4X1 U2362 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n2089), .S1(n2071), 
        .Y(n1809) );
  MXI4X1 U2363 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n2088), .S1(n2071), 
        .Y(n1805) );
  MXI4X1 U2364 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1817) );
  MXI4X1 U2365 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1813) );
  MXI4X1 U2366 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n2090), .S1(n2072), 
        .Y(n1825) );
  MXI4X1 U2367 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n2089), .S1(n2071), 
        .Y(n1821) );
  MXI4X1 U2368 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1833) );
  MXI4X1 U2369 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1829) );
  MXI4X1 U2370 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n2091), .S1(n2072), 
        .Y(n1841) );
  MXI4X1 U2371 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n2090), .S1(n2072), 
        .Y(n1837) );
  MXI4X1 U2372 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n2091), .S1(n2073), 
        .Y(n1849) );
  MXI4X1 U2373 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n2091), .S1(n2072), 
        .Y(n1845) );
  MXI4X1 U2374 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n2092), .S1(n2073), 
        .Y(n1857) );
  MXI4X1 U2375 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n2091), .S1(n2073), 
        .Y(n1853) );
  MXI4X1 U2376 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1865) );
  MXI4X1 U2377 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1861) );
  MXI4X1 U2378 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n2092), .S1(n2074), 
        .Y(n1873) );
  MXI4X1 U2379 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n2092), .S1(n2073), 
        .Y(n1869) );
  MXI4X1 U2380 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1881) );
  MXI4X1 U2381 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1877) );
  MXI4X1 U2382 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1889) );
  MXI4X1 U2383 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1885) );
  MXI4X1 U2384 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n2094), .S1(n2075), 
        .Y(n1897) );
  MXI4X1 U2385 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n2094), .S1(n2074), 
        .Y(n1893) );
  MXI4X1 U2386 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1569), .S1(n1550), .Y(
        n1122) );
  MXI4X1 U2387 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1569), .S1(n1550), .Y(
        n1118) );
  MXI4X1 U2388 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1569), .S1(n1550), .Y(
        n1126) );
  MXI4X1 U2389 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1570), .S1(n1550), .Y(
        n1130) );
  MXI4X1 U2390 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1570), .S1(n1550), .Y(
        n1134) );
  MXI4X1 U2391 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1570), .S1(n1550), .Y(
        n1138) );
  MXI4X1 U2392 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1570), .S1(n1551), .Y(
        n1142) );
  MXI4X1 U2393 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1571), .S1(n1551), .Y(
        n1146) );
  MXI4X1 U2394 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1571), .S1(n1551), .Y(
        n1150) );
  MXI4X1 U2395 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1571), .S1(n1551), .Y(
        n1154) );
  MXI4X1 U2396 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1571), .S1(n1551), .Y(
        n1158) );
  MXI4X1 U2397 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1572), .S1(n1551), .Y(
        n1162) );
  MXI4X1 U2398 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1572), .S1(n1551), .Y(
        n1166) );
  MXI4X1 U2399 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1572), .S1(n1558), .Y(
        n1170) );
  MXI4X1 U2400 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1572), .S1(n1545), .Y(
        n1174) );
  MXI4X1 U2401 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1572), .S1(n1557), .Y(
        n1178) );
  MXI4X1 U2402 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1576), .S1(n1552), .Y(
        n1182) );
  MXI4X1 U2403 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1573), .S1(n1558), .Y(
        n1186) );
  MXI4X1 U2404 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1573), .S1(n1558), .Y(
        n1190) );
  MXI4X1 U2405 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1573), .S1(n1557), .Y(
        n1194) );
  MXI4X1 U2406 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1574), .S1(n1556), 
        .Y(n1198) );
  MXI4X1 U2407 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1574), .S1(n1545), 
        .Y(n1202) );
  MXI4X1 U2408 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1574), .S1(n1557), 
        .Y(n1206) );
  MXI4X1 U2409 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1574), .S1(n1553), 
        .Y(n1210) );
  MXI4X1 U2410 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1575), .S1(n1555), 
        .Y(n1214) );
  MXI4X1 U2411 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1575), .S1(n1557), 
        .Y(n1218) );
  MXI4X1 U2412 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1575), .S1(n1558), 
        .Y(n1222) );
  MXI4X1 U2413 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1575), .S1(n1556), 
        .Y(n1226) );
  MXI4X1 U2414 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1575), .S1(n1551), 
        .Y(n1230) );
  MXI4X1 U2415 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1576), .S1(n1551), 
        .Y(n1234) );
  MXI4X1 U2416 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1576), .S1(n1558), 
        .Y(n1238) );
  MXI4X1 U2417 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1576), .S1(n1552), 
        .Y(n1242) );
  MXI4X1 U2418 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1250) );
  MXI4X1 U2419 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1246) );
  MXI4X1 U2420 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1258) );
  MXI4X1 U2421 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1254) );
  MXI4X1 U2422 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1563), .S1(n1546), 
        .Y(n1266) );
  MXI4X1 U2423 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1562), .S1(n1546), 
        .Y(n1262) );
  MXI4X1 U2424 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1563), .S1(n1549), 
        .Y(n1274) );
  MXI4X1 U2425 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1563), .S1(n1546), 
        .Y(n1270) );
  MXI4X1 U2426 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1564), .S1(n1549), 
        .Y(n1282) );
  MXI4X1 U2427 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1563), .S1(n1544), 
        .Y(n1278) );
  MXI4X1 U2428 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1564), .S1(n1556), 
        .Y(n1290) );
  MXI4X1 U2429 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1564), .S1(n1545), 
        .Y(n1286) );
  MXI4X1 U2430 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1565), .S1(n1547), 
        .Y(n1298) );
  MXI4X1 U2431 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1564), .S1(n1545), 
        .Y(n1294) );
  MXI4X1 U2432 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1306) );
  MXI4X1 U2433 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1302) );
  MXI4X1 U2434 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1566), .S1(n1547), 
        .Y(n1314) );
  MXI4X1 U2435 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1565), .S1(n1547), 
        .Y(n1310) );
  MXI4X1 U2436 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1566), .S1(n1548), 
        .Y(n1322) );
  MXI4X1 U2437 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1566), .S1(n1547), 
        .Y(n1318) );
  MXI4X1 U2438 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1567), .S1(n1548), 
        .Y(n1330) );
  MXI4X1 U2439 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1566), .S1(n1548), 
        .Y(n1326) );
  MXI4X1 U2440 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1338) );
  MXI4X1 U2441 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1334) );
  MXI4X1 U2442 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1567), .S1(n1549), 
        .Y(n1346) );
  MXI4X1 U2443 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1567), .S1(n1548), 
        .Y(n1342) );
  MXI4X1 U2444 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1354) );
  MXI4X1 U2445 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1350) );
  MXI4X1 U2446 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1362) );
  MXI4X1 U2447 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1358) );
  MXI4X1 U2448 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1569), .S1(n1550), 
        .Y(n1370) );
  MXI4X1 U2449 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1569), .S1(n1549), 
        .Y(n1366) );
  MXI4X1 U2450 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n2094), .S1(n2075), .Y(
        n1650) );
  MXI4X1 U2451 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n2094), .S1(n2075), .Y(
        n1646) );
  MXI4X1 U2452 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n2094), .S1(n2075), .Y(
        n1654) );
  MXI4X1 U2453 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n2095), .S1(n2075), .Y(
        n1662) );
  MXI4X1 U2454 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n2095), .S1(n2076), .Y(
        n1670) );
  MXI4X1 U2455 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n2096), .S1(n2076), .Y(
        n1678) );
  MXI4X1 U2456 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n2096), .S1(n2076), .Y(
        n1686) );
  MXI4X1 U2457 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n2097), .S1(n2077), .Y(
        n1694) );
  MXI4X1 U2458 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n2097), .S1(n2077), .Y(
        n1702) );
  MXI4X1 U2459 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n2098), .S1(n2077), .Y(
        n1710) );
  MXI4X1 U2460 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n2098), .S1(n2075), .Y(
        n1718) );
  MXI4X1 U2461 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n2099), .S1(n2070), 
        .Y(n1726) );
  MXI4X1 U2462 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n2099), .S1(n2080), 
        .Y(n1734) );
  MXI4X1 U2463 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n2100), .S1(n2078), 
        .Y(n1742) );
  MXI4X1 U2464 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n2100), .S1(n2078), 
        .Y(n1750) );
  MXI4X1 U2465 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n2101), .S1(n2078), 
        .Y(n1758) );
  MXI4X1 U2466 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n2101), .S1(n2078), 
        .Y(n1766) );
  MXI4X1 U2467 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1778) );
  MXI4X1 U2468 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n2087), .S1(n2070), 
        .Y(n1774) );
  MXI4X1 U2469 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1786) );
  MXI4X1 U2470 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n2087), .S1(n2070), 
        .Y(n1782) );
  MXI4X1 U2471 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n2088), .S1(n2070), 
        .Y(n1794) );
  MXI4X1 U2472 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n2088), .S1(n2070), 
        .Y(n1790) );
  MXI4X1 U2473 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n2088), .S1(n2071), 
        .Y(n1802) );
  MXI4X1 U2474 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n2088), .S1(n2071), 
        .Y(n1798) );
  MXI4X1 U2475 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n2089), .S1(n2071), 
        .Y(n1810) );
  MXI4X1 U2476 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n2088), .S1(n2071), 
        .Y(n1806) );
  MXI4X1 U2477 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1818) );
  MXI4X1 U2478 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n2089), .S1(n2071), 
        .Y(n1814) );
  MXI4X1 U2479 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n2090), .S1(n2072), 
        .Y(n1826) );
  MXI4X1 U2480 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n2089), .S1(n2071), 
        .Y(n1822) );
  MXI4X1 U2481 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1834) );
  MXI4X1 U2482 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n2090), .S1(n2072), 
        .Y(n1830) );
  MXI4X1 U2483 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n2091), .S1(n2072), 
        .Y(n1842) );
  MXI4X1 U2484 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n2090), .S1(n2072), 
        .Y(n1838) );
  MXI4X1 U2485 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n2091), .S1(n2073), 
        .Y(n1850) );
  MXI4X1 U2486 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n2091), .S1(n2072), 
        .Y(n1846) );
  MXI4X1 U2487 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n2092), .S1(n2073), 
        .Y(n1858) );
  MXI4X1 U2488 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n2091), .S1(n2073), 
        .Y(n1854) );
  MXI4X1 U2489 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1866) );
  MXI4X1 U2490 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n2092), .S1(n2073), 
        .Y(n1862) );
  MXI4X1 U2491 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n2093), .S1(n2074), 
        .Y(n1874) );
  MXI4X1 U2492 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n2092), .S1(n2073), 
        .Y(n1870) );
  MXI4X1 U2493 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1882) );
  MXI4X1 U2494 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n2093), .S1(n2074), 
        .Y(n1878) );
  MXI4X1 U2495 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1890) );
  MXI4X1 U2496 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n2093), .S1(n2074), 
        .Y(n1886) );
  MXI4X1 U2497 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n2090), .S1(n2072), 
        .Y(n1898) );
  MXI4X1 U2498 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n2094), .S1(n2074), 
        .Y(n1894) );
  MXI4X1 U2499 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1569), .S1(n1550), .Y(
        n1123) );
  MXI4X1 U2500 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1569), .S1(n1550), .Y(
        n1119) );
  MXI4X1 U2501 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1569), .S1(n1550), .Y(
        n1127) );
  MXI4X1 U2502 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1570), .S1(n1550), .Y(
        n1135) );
  MXI4X1 U2503 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1570), .S1(n1551), .Y(
        n1143) );
  MXI4X1 U2504 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1571), .S1(n1551), .Y(
        n1151) );
  MXI4X1 U2505 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1571), .S1(n1551), .Y(
        n1159) );
  MXI4X1 U2506 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1572), .S1(n1554), .Y(
        n1167) );
  MXI4X1 U2507 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1572), .S1(n1556), .Y(
        n1175) );
  MXI4X1 U2508 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1573), .S1(n1554), .Y(
        n1183) );
  MXI4X1 U2509 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1573), .S1(n1544), .Y(
        n1191) );
  MXI4X1 U2510 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1574), .S1(n1554), 
        .Y(n1199) );
  MXI4X1 U2511 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1574), .S1(n1545), 
        .Y(n1207) );
  MXI4X1 U2512 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1575), .S1(n1557), 
        .Y(n1215) );
  MXI4X1 U2513 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1575), .S1(n1556), 
        .Y(n1223) );
  MXI4X1 U2514 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1576), .S1(n1549), 
        .Y(n1231) );
  MXI4X1 U2515 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1576), .S1(n1547), 
        .Y(n1239) );
  MXI4X1 U2516 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1251) );
  MXI4X1 U2517 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1562), .S1(n1546), 
        .Y(n1247) );
  MXI4X1 U2518 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1259) );
  MXI4X1 U2519 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1562), .S1(n1546), 
        .Y(n1255) );
  MXI4X1 U2520 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1563), .S1(n1546), 
        .Y(n1267) );
  MXI4X1 U2521 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1563), .S1(n1546), 
        .Y(n1263) );
  MXI4X1 U2522 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1563), .S1(n1555), 
        .Y(n1275) );
  MXI4X1 U2523 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1563), .S1(N13), .Y(
        n1271) );
  MXI4X1 U2524 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1564), .S1(n1545), 
        .Y(n1283) );
  MXI4X1 U2525 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1563), .S1(n1555), 
        .Y(n1279) );
  MXI4X1 U2526 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1564), .S1(n1544), 
        .Y(n1291) );
  MXI4X1 U2527 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1564), .S1(n1545), 
        .Y(n1287) );
  MXI4X1 U2528 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1565), .S1(n1547), 
        .Y(n1299) );
  MXI4X1 U2529 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1564), .S1(n1555), 
        .Y(n1295) );
  MXI4X1 U2530 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1307) );
  MXI4X1 U2531 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1565), .S1(n1547), 
        .Y(n1303) );
  MXI4X1 U2532 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1566), .S1(n1547), 
        .Y(n1315) );
  MXI4X1 U2533 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1565), .S1(n1547), 
        .Y(n1311) );
  MXI4X1 U2534 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1566), .S1(n1548), 
        .Y(n1323) );
  MXI4X1 U2535 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1566), .S1(n1547), 
        .Y(n1319) );
  MXI4X1 U2536 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1567), .S1(n1548), 
        .Y(n1331) );
  MXI4X1 U2537 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1566), .S1(n1548), 
        .Y(n1327) );
  MXI4X1 U2538 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1339) );
  MXI4X1 U2539 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1567), .S1(n1548), 
        .Y(n1335) );
  MXI4X1 U2540 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1568), .S1(n1549), 
        .Y(n1347) );
  MXI4X1 U2541 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1567), .S1(n1548), 
        .Y(n1343) );
  MXI4X1 U2542 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1355) );
  MXI4X1 U2543 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1568), .S1(n1549), 
        .Y(n1351) );
  MXI4X1 U2544 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1363) );
  MXI4X1 U2545 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1568), .S1(n1549), 
        .Y(n1359) );
  MXI4X1 U2546 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1565), .S1(n1547), 
        .Y(n1371) );
  MXI4X1 U2547 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1569), .S1(n1549), 
        .Y(n1367) );
  NOR3X1 U2548 ( .A(wsel[1]), .B(wsel[2]), .C(wsel[0]), .Y(n82) );
  XNOR2XL U2549 ( .A(N13), .B(wsel[1]), .Y(n57) );
  XNOR2XL U2550 ( .A(N18), .B(wsel[1]), .Y(n48) );
  NOR3X1 U2551 ( .A(wsel[1]), .B(wsel[2]), .C(n2454), .Y(n66) );
  XNOR2XL U2552 ( .A(N14), .B(wsel[2]), .Y(n59) );
  XNOR2XL U2553 ( .A(N19), .B(wsel[2]), .Y(n50) );
endmodule


module extender ( shamt_i, immed_i, ExtOp_i, ExtOut_o );
  input [4:0] shamt_i;
  input [15:0] immed_i;
  output [31:0] ExtOut_o;
  input ExtOp_i;
  wire   n2, n1, n19, n20;

  INVX3 U1 ( .A(ExtOp_i), .Y(n20) );
  INVX3 U2 ( .A(ExtOut_o[30]), .Y(n1) );
  AO22X1 U3 ( .A0(shamt_i[1]), .A1(ExtOp_i), .B0(immed_i[1]), .B1(n20), .Y(
        ExtOut_o[1]) );
  AO22X1 U4 ( .A0(shamt_i[2]), .A1(ExtOp_i), .B0(immed_i[2]), .B1(n20), .Y(
        ExtOut_o[2]) );
  AO22X1 U5 ( .A0(shamt_i[3]), .A1(ExtOp_i), .B0(immed_i[3]), .B1(n20), .Y(
        ExtOut_o[3]) );
  OAI2BB1X1 U6 ( .A0N(immed_i[4]), .A1N(n20), .B0(n19), .Y(ExtOut_o[4]) );
  OAI2BB1X1 U7 ( .A0N(immed_i[5]), .A1N(n20), .B0(n19), .Y(ExtOut_o[5]) );
  OAI2BB1X1 U8 ( .A0N(immed_i[6]), .A1N(n20), .B0(n19), .Y(ExtOut_o[6]) );
  OAI2BB1X1 U9 ( .A0N(immed_i[7]), .A1N(n20), .B0(n19), .Y(ExtOut_o[7]) );
  OAI2BB1X1 U10 ( .A0N(immed_i[8]), .A1N(n20), .B0(n19), .Y(ExtOut_o[8]) );
  OAI2BB1X1 U11 ( .A0N(immed_i[9]), .A1N(n20), .B0(n19), .Y(ExtOut_o[9]) );
  OAI2BB1X1 U12 ( .A0N(immed_i[10]), .A1N(n20), .B0(n19), .Y(ExtOut_o[10]) );
  OAI2BB1X1 U13 ( .A0N(immed_i[11]), .A1N(n20), .B0(n19), .Y(ExtOut_o[11]) );
  OAI2BB1X1 U14 ( .A0N(immed_i[12]), .A1N(n20), .B0(n19), .Y(ExtOut_o[12]) );
  OAI2BB1X1 U15 ( .A0N(immed_i[13]), .A1N(n20), .B0(n19), .Y(ExtOut_o[13]) );
  OAI2BB1X1 U16 ( .A0N(immed_i[14]), .A1N(n20), .B0(n19), .Y(ExtOut_o[14]) );
  CLKINVX1 U17 ( .A(n1), .Y(ExtOut_o[15]) );
  CLKINVX1 U18 ( .A(n1), .Y(ExtOut_o[16]) );
  CLKINVX1 U19 ( .A(n1), .Y(ExtOut_o[17]) );
  CLKINVX1 U20 ( .A(n1), .Y(ExtOut_o[18]) );
  CLKINVX1 U21 ( .A(n1), .Y(ExtOut_o[19]) );
  CLKINVX1 U22 ( .A(n1), .Y(ExtOut_o[20]) );
  CLKINVX1 U23 ( .A(n1), .Y(ExtOut_o[21]) );
  CLKINVX1 U24 ( .A(n1), .Y(ExtOut_o[22]) );
  CLKINVX1 U25 ( .A(n1), .Y(ExtOut_o[23]) );
  CLKINVX1 U26 ( .A(n1), .Y(ExtOut_o[24]) );
  CLKINVX1 U27 ( .A(n1), .Y(ExtOut_o[25]) );
  CLKINVX1 U28 ( .A(n1), .Y(ExtOut_o[26]) );
  CLKINVX1 U29 ( .A(n1), .Y(ExtOut_o[27]) );
  CLKINVX1 U30 ( .A(n1), .Y(ExtOut_o[28]) );
  CLKINVX1 U31 ( .A(n1), .Y(ExtOut_o[29]) );
  CLKINVX1 U32 ( .A(n1), .Y(ExtOut_o[31]) );
  AO22X1 U33 ( .A0(shamt_i[0]), .A1(ExtOp_i), .B0(immed_i[0]), .B1(n20), .Y(
        ExtOut_o[0]) );
  CLKBUFX3 U34 ( .A(n2), .Y(n19) );
  NAND2X1 U35 ( .A(shamt_i[4]), .B(ExtOp_i), .Y(n2) );
  OAI2BB1X1 U36 ( .A0N(immed_i[15]), .A1N(n20), .B0(n19), .Y(ExtOut_o[30]) );
endmodule


module MUX_5_3to1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [4:0] data0_i;
  input [4:0] data1_i;
  input [4:0] data2_i;
  input [1:0] select_i;
  output [4:0] data_o;
  wire   n6, n7, n8, n9, n10, n11, n12, n13;

  NOR2BX1 U2 ( .AN(select_i[1]), .B(select_i[0]), .Y(n8) );
  NOR2BX1 U3 ( .AN(select_i[0]), .B(select_i[1]), .Y(n9) );
  NOR2X1 U4 ( .A(select_i[0]), .B(select_i[1]), .Y(n7) );
  CLKINVX1 U5 ( .A(n12), .Y(data_o[1]) );
  AOI222XL U6 ( .A0(data0_i[1]), .A1(n7), .B0(data2_i[1]), .B1(n8), .C0(
        data1_i[1]), .C1(n9), .Y(n12) );
  CLKINVX1 U7 ( .A(n11), .Y(data_o[2]) );
  AOI222XL U8 ( .A0(data0_i[2]), .A1(n7), .B0(data2_i[2]), .B1(n8), .C0(
        data1_i[2]), .C1(n9), .Y(n11) );
  CLKINVX1 U9 ( .A(n10), .Y(data_o[3]) );
  AOI222XL U10 ( .A0(data0_i[3]), .A1(n7), .B0(data2_i[3]), .B1(n8), .C0(
        data1_i[3]), .C1(n9), .Y(n10) );
  CLKINVX1 U11 ( .A(n13), .Y(data_o[0]) );
  AOI222XL U12 ( .A0(data0_i[0]), .A1(n7), .B0(data2_i[0]), .B1(n8), .C0(
        data1_i[0]), .C1(n9), .Y(n13) );
  CLKINVX1 U13 ( .A(n6), .Y(data_o[4]) );
  AOI222XL U14 ( .A0(data0_i[4]), .A1(n7), .B0(data2_i[4]), .B1(n8), .C0(
        data1_i[4]), .C1(n9), .Y(n6) );
endmodule


module MUX_32_3to1_0 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AO21X2 U2 ( .A0(data0_i[1]), .A1(n9), .B0(n14), .Y(data_o[1]) );
  AO21X2 U3 ( .A0(data0_i[6]), .A1(n9), .B0(n19), .Y(data_o[6]) );
  AO21X2 U4 ( .A0(data0_i[2]), .A1(n9), .B0(n15), .Y(data_o[2]) );
  CLKBUFX8 U5 ( .A(n3), .Y(n9) );
  BUFX8 U6 ( .A(n4), .Y(n7) );
  CLKAND2X2 U7 ( .A(select_i[1]), .B(n11), .Y(n4) );
  AO21X2 U8 ( .A0(data0_i[13]), .A1(n9), .B0(n25), .Y(data_o[13]) );
  OR2X1 U9 ( .A(n1), .B(n34), .Y(data_o[22]) );
  AO22X1 U10 ( .A0(data2_i[6]), .A1(n7), .B0(data1_i[6]), .B1(n6), .Y(n19) );
  AOI22X1 U11 ( .A0(data2_i[10]), .A1(n7), .B0(data1_i[10]), .B1(n6), .Y(n2)
         );
  AO21X4 U12 ( .A0(data0_i[11]), .A1(n9), .B0(n23), .Y(data_o[11]) );
  AND2X8 U13 ( .A(select_i[0]), .B(n12), .Y(n5) );
  AND2X2 U14 ( .A(n12), .B(n11), .Y(n3) );
  BUFX4 U15 ( .A(n5), .Y(n6) );
  AO22XL U16 ( .A0(data2_i[21]), .A1(n7), .B0(data1_i[21]), .B1(n5), .Y(n33)
         );
  AO21X4 U17 ( .A0(data0_i[25]), .A1(n9), .B0(n37), .Y(data_o[25]) );
  AO22XL U18 ( .A0(data2_i[13]), .A1(n7), .B0(data1_i[13]), .B1(n5), .Y(n25)
         );
  AO21X4 U19 ( .A0(data0_i[18]), .A1(n9), .B0(n30), .Y(data_o[18]) );
  AO22XL U20 ( .A0(data2_i[18]), .A1(n7), .B0(data1_i[18]), .B1(n5), .Y(n30)
         );
  AO21X4 U21 ( .A0(data0_i[12]), .A1(n9), .B0(n24), .Y(data_o[12]) );
  AO22XL U22 ( .A0(data2_i[12]), .A1(n7), .B0(data1_i[12]), .B1(n5), .Y(n24)
         );
  AO21X4 U23 ( .A0(data0_i[21]), .A1(n9), .B0(n33), .Y(data_o[21]) );
  AO21X4 U24 ( .A0(data0_i[3]), .A1(n9), .B0(n16), .Y(data_o[3]) );
  AND2XL U25 ( .A(data0_i[22]), .B(n9), .Y(n1) );
  INVX2 U26 ( .A(select_i[0]), .Y(n11) );
  INVX2 U27 ( .A(select_i[1]), .Y(n12) );
  OAI2BB1X1 U28 ( .A0N(data0_i[10]), .A1N(n9), .B0(n2), .Y(data_o[10]) );
  CLKBUFX2 U29 ( .A(n3), .Y(n10) );
  CLKBUFX3 U30 ( .A(n4), .Y(n8) );
  AO21X1 U31 ( .A0(data0_i[0]), .A1(n9), .B0(n13), .Y(data_o[0]) );
  AO22X1 U32 ( .A0(data2_i[0]), .A1(n7), .B0(data1_i[0]), .B1(n6), .Y(n13) );
  AO22X1 U33 ( .A0(data2_i[1]), .A1(n7), .B0(data1_i[1]), .B1(n6), .Y(n14) );
  AO21X1 U34 ( .A0(data0_i[4]), .A1(n9), .B0(n17), .Y(data_o[4]) );
  AO22X1 U35 ( .A0(data2_i[4]), .A1(n7), .B0(data1_i[4]), .B1(n6), .Y(n17) );
  AO21X1 U36 ( .A0(data0_i[5]), .A1(n9), .B0(n18), .Y(data_o[5]) );
  AO22X1 U37 ( .A0(data2_i[5]), .A1(n7), .B0(data1_i[5]), .B1(n6), .Y(n18) );
  AO21X1 U38 ( .A0(data0_i[19]), .A1(n9), .B0(n31), .Y(data_o[19]) );
  AO22X1 U39 ( .A0(data2_i[19]), .A1(n7), .B0(data1_i[19]), .B1(n5), .Y(n31)
         );
  AO22X1 U40 ( .A0(data2_i[22]), .A1(n7), .B0(data1_i[22]), .B1(n5), .Y(n34)
         );
  AO21X1 U41 ( .A0(data0_i[23]), .A1(n9), .B0(n35), .Y(data_o[23]) );
  AO22X1 U42 ( .A0(data2_i[23]), .A1(n7), .B0(data1_i[23]), .B1(n5), .Y(n35)
         );
  AO21X1 U43 ( .A0(data0_i[24]), .A1(n9), .B0(n36), .Y(data_o[24]) );
  AO22X1 U44 ( .A0(data2_i[24]), .A1(n8), .B0(data1_i[24]), .B1(n5), .Y(n36)
         );
  AO21X1 U45 ( .A0(data0_i[27]), .A1(n10), .B0(n39), .Y(data_o[27]) );
  AO22X1 U46 ( .A0(data2_i[27]), .A1(n8), .B0(data1_i[27]), .B1(n6), .Y(n39)
         );
  AO22X1 U47 ( .A0(data2_i[3]), .A1(n7), .B0(data1_i[3]), .B1(n6), .Y(n16) );
  AO21X1 U48 ( .A0(data0_i[15]), .A1(n9), .B0(n27), .Y(data_o[15]) );
  AO22X1 U49 ( .A0(data2_i[15]), .A1(n7), .B0(data1_i[15]), .B1(n5), .Y(n27)
         );
  AO21X1 U50 ( .A0(data0_i[29]), .A1(n10), .B0(n41), .Y(data_o[29]) );
  AO22X1 U51 ( .A0(data2_i[29]), .A1(n8), .B0(data1_i[29]), .B1(n5), .Y(n41)
         );
  AO22X1 U52 ( .A0(data2_i[2]), .A1(n7), .B0(data1_i[2]), .B1(n6), .Y(n15) );
  AO21X1 U53 ( .A0(data0_i[31]), .A1(n10), .B0(n43), .Y(data_o[31]) );
  AO22X1 U54 ( .A0(data2_i[31]), .A1(n8), .B0(data1_i[31]), .B1(n5), .Y(n43)
         );
  AO21X1 U55 ( .A0(data0_i[30]), .A1(n10), .B0(n42), .Y(data_o[30]) );
  AO22X1 U56 ( .A0(data2_i[30]), .A1(n8), .B0(data1_i[30]), .B1(n5), .Y(n42)
         );
  AO21X1 U57 ( .A0(data0_i[7]), .A1(n9), .B0(n20), .Y(data_o[7]) );
  AO22X1 U58 ( .A0(data2_i[7]), .A1(n7), .B0(data1_i[7]), .B1(n6), .Y(n20) );
  AO21X1 U59 ( .A0(data0_i[14]), .A1(n9), .B0(n26), .Y(data_o[14]) );
  AO22X1 U60 ( .A0(data2_i[14]), .A1(n7), .B0(data1_i[14]), .B1(n5), .Y(n26)
         );
  AO21X1 U61 ( .A0(data0_i[17]), .A1(n9), .B0(n29), .Y(data_o[17]) );
  AO22X1 U62 ( .A0(data2_i[17]), .A1(n7), .B0(data1_i[17]), .B1(n5), .Y(n29)
         );
  AO21X1 U63 ( .A0(data0_i[26]), .A1(n10), .B0(n38), .Y(data_o[26]) );
  AO22X1 U64 ( .A0(data2_i[26]), .A1(n8), .B0(data1_i[26]), .B1(n5), .Y(n38)
         );
  AO22X1 U65 ( .A0(data2_i[11]), .A1(n7), .B0(data1_i[11]), .B1(n6), .Y(n23)
         );
  AO21X1 U66 ( .A0(data0_i[8]), .A1(n9), .B0(n21), .Y(data_o[8]) );
  AO22X1 U67 ( .A0(data2_i[8]), .A1(n7), .B0(data1_i[8]), .B1(n6), .Y(n21) );
  AO21X1 U68 ( .A0(data0_i[9]), .A1(n9), .B0(n22), .Y(data_o[9]) );
  AO22X1 U69 ( .A0(data2_i[9]), .A1(n7), .B0(data1_i[9]), .B1(n6), .Y(n22) );
  AO21X1 U70 ( .A0(data0_i[28]), .A1(n10), .B0(n40), .Y(data_o[28]) );
  AO22X1 U71 ( .A0(data2_i[28]), .A1(n8), .B0(data1_i[28]), .B1(n6), .Y(n40)
         );
  AO21X1 U72 ( .A0(data0_i[16]), .A1(n9), .B0(n28), .Y(data_o[16]) );
  AO22X1 U73 ( .A0(data2_i[16]), .A1(n7), .B0(data1_i[16]), .B1(n5), .Y(n28)
         );
  AO21X1 U74 ( .A0(data0_i[20]), .A1(n9), .B0(n32), .Y(data_o[20]) );
  AO22X1 U75 ( .A0(data2_i[20]), .A1(n7), .B0(data1_i[20]), .B1(n5), .Y(n32)
         );
  AO22XL U76 ( .A0(data2_i[25]), .A1(n8), .B0(data1_i[25]), .B1(n5), .Y(n37)
         );
endmodule


module MUX_32_3to1_2 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  BUFX12 U2 ( .A(n18), .Y(n1) );
  BUFX16 U3 ( .A(n18), .Y(n2) );
  CLKAND2X6 U4 ( .A(select_i[0]), .B(n21), .Y(n18) );
  OAI2BB1X2 U5 ( .A0N(data0_i[30]), .A1N(n16), .B0(n15), .Y(data_o[30]) );
  CLKINVX1 U6 ( .A(select_i[1]), .Y(n21) );
  BUFX16 U7 ( .A(n17), .Y(n9) );
  OR2X6 U8 ( .A(n8), .B(n36), .Y(data_o[16]) );
  AO22X1 U9 ( .A0(data2_i[16]), .A1(n10), .B0(data1_i[16]), .B1(n1), .Y(n36)
         );
  AO22X1 U10 ( .A0(data2_i[10]), .A1(n11), .B0(data1_i[10]), .B1(n1), .Y(n30)
         );
  AND2X8 U11 ( .A(n21), .B(n20), .Y(n16) );
  INVX4 U12 ( .A(select_i[0]), .Y(n20) );
  AO22X4 U13 ( .A0(data2_i[3]), .A1(n11), .B0(data1_i[3]), .B1(n1), .Y(n23) );
  AO22X2 U14 ( .A0(data2_i[11]), .A1(n11), .B0(data1_i[11]), .B1(n1), .Y(n31)
         );
  AO22X4 U15 ( .A0(data2_i[0]), .A1(n11), .B0(data1_i[0]), .B1(n2), .Y(n14) );
  AO22X4 U16 ( .A0(data2_i[7]), .A1(n11), .B0(data1_i[7]), .B1(n2), .Y(n27) );
  AO22X4 U17 ( .A0(data2_i[2]), .A1(n10), .B0(data1_i[2]), .B1(n1), .Y(n13) );
  AO22X1 U18 ( .A0(data2_i[5]), .A1(n10), .B0(data1_i[5]), .B1(n2), .Y(n25) );
  AO22X4 U19 ( .A0(data2_i[4]), .A1(n11), .B0(data1_i[4]), .B1(n2), .Y(n24) );
  CLKAND2X12 U20 ( .A(select_i[1]), .B(n20), .Y(n17) );
  AO22X4 U21 ( .A0(data2_i[20]), .A1(n10), .B0(data1_i[20]), .B1(n2), .Y(n40)
         );
  AO22X1 U22 ( .A0(n10), .A1(data2_i[25]), .B0(data1_i[25]), .B1(n2), .Y(n43)
         );
  AO22X4 U23 ( .A0(data2_i[14]), .A1(n10), .B0(data1_i[14]), .B1(n2), .Y(n34)
         );
  AO22X4 U24 ( .A0(data2_i[15]), .A1(n10), .B0(data1_i[15]), .B1(n2), .Y(n35)
         );
  BUFX20 U25 ( .A(n9), .Y(n10) );
  AND2X1 U26 ( .A(data0_i[25]), .B(n16), .Y(n3) );
  OR2X8 U27 ( .A(n3), .B(n43), .Y(data_o[25]) );
  AND2X2 U28 ( .A(data0_i[27]), .B(n16), .Y(n4) );
  OR2X8 U29 ( .A(n4), .B(n45), .Y(data_o[27]) );
  AO22X1 U30 ( .A0(data2_i[27]), .A1(n11), .B0(data1_i[27]), .B1(n1), .Y(n45)
         );
  AND2X1 U31 ( .A(data0_i[18]), .B(n16), .Y(n5) );
  OR2X8 U32 ( .A(n5), .B(n38), .Y(data_o[18]) );
  AO22X1 U33 ( .A0(data2_i[18]), .A1(n11), .B0(data1_i[18]), .B1(n1), .Y(n38)
         );
  AND2X1 U34 ( .A(data0_i[23]), .B(n16), .Y(n6) );
  OR2X8 U35 ( .A(n6), .B(n12), .Y(data_o[23]) );
  AO22XL U36 ( .A0(data2_i[23]), .A1(n11), .B0(data1_i[23]), .B1(n2), .Y(n12)
         );
  CLKAND2X2 U37 ( .A(data0_i[17]), .B(n16), .Y(n7) );
  OR2X8 U38 ( .A(n7), .B(n37), .Y(data_o[17]) );
  AND2X1 U39 ( .A(data0_i[16]), .B(n16), .Y(n8) );
  AO22X4 U40 ( .A0(data2_i[22]), .A1(n11), .B0(data1_i[22]), .B1(n2), .Y(n42)
         );
  BUFX20 U41 ( .A(n9), .Y(n11) );
  AO22X4 U42 ( .A0(data2_i[26]), .A1(n10), .B0(data1_i[26]), .B1(n2), .Y(n44)
         );
  AO21X4 U43 ( .A0(data0_i[2]), .A1(n16), .B0(n13), .Y(data_o[2]) );
  AO21X4 U44 ( .A0(data0_i[0]), .A1(n16), .B0(n14), .Y(data_o[0]) );
  AOI22XL U45 ( .A0(data2_i[30]), .A1(n11), .B0(data1_i[30]), .B1(n2), .Y(n15)
         );
  AO21X4 U46 ( .A0(data0_i[10]), .A1(n16), .B0(n30), .Y(data_o[10]) );
  OAI2BB1X4 U47 ( .A0N(data0_i[24]), .A1N(n16), .B0(n19), .Y(data_o[24]) );
  AOI22X1 U48 ( .A0(data2_i[24]), .A1(n10), .B0(data1_i[24]), .B1(n2), .Y(n19)
         );
  AO22X1 U49 ( .A0(data2_i[17]), .A1(n10), .B0(data1_i[17]), .B1(n2), .Y(n37)
         );
  AO21X1 U50 ( .A0(data0_i[13]), .A1(n16), .B0(n33), .Y(data_o[13]) );
  AO22X1 U51 ( .A0(data2_i[13]), .A1(n10), .B0(data1_i[13]), .B1(n1), .Y(n33)
         );
  AO21X2 U52 ( .A0(data0_i[22]), .A1(n16), .B0(n42), .Y(data_o[22]) );
  AO22X4 U53 ( .A0(data2_i[12]), .A1(n11), .B0(data1_i[12]), .B1(n2), .Y(n32)
         );
  AO22X1 U54 ( .A0(data2_i[8]), .A1(n10), .B0(data1_i[8]), .B1(n1), .Y(n28) );
  AO22X1 U55 ( .A0(data2_i[9]), .A1(n11), .B0(data1_i[9]), .B1(n2), .Y(n29) );
  AO22X1 U56 ( .A0(data2_i[28]), .A1(n10), .B0(data1_i[28]), .B1(n2), .Y(n46)
         );
  AO21X2 U57 ( .A0(data0_i[15]), .A1(n16), .B0(n35), .Y(data_o[15]) );
  AO22X2 U58 ( .A0(data2_i[21]), .A1(n11), .B0(data1_i[21]), .B1(n2), .Y(n41)
         );
  AO22X2 U59 ( .A0(data2_i[29]), .A1(n10), .B0(data1_i[29]), .B1(n2), .Y(n47)
         );
  AO22X4 U60 ( .A0(data2_i[1]), .A1(n11), .B0(data1_i[1]), .B1(n2), .Y(n22) );
  AO21X4 U61 ( .A0(data0_i[1]), .A1(n16), .B0(n22), .Y(data_o[1]) );
  AO21X4 U62 ( .A0(data0_i[3]), .A1(n16), .B0(n23), .Y(data_o[3]) );
  AO21X4 U63 ( .A0(data0_i[4]), .A1(n16), .B0(n24), .Y(data_o[4]) );
  AO21X4 U64 ( .A0(data0_i[5]), .A1(n16), .B0(n25), .Y(data_o[5]) );
  AO22X4 U65 ( .A0(data2_i[6]), .A1(n11), .B0(data1_i[6]), .B1(n1), .Y(n26) );
  AO21X4 U66 ( .A0(data0_i[6]), .A1(n16), .B0(n26), .Y(data_o[6]) );
  AO21X4 U67 ( .A0(data0_i[7]), .A1(n16), .B0(n27), .Y(data_o[7]) );
  AO21X4 U68 ( .A0(data0_i[8]), .A1(n16), .B0(n28), .Y(data_o[8]) );
  AO21X4 U69 ( .A0(data0_i[9]), .A1(n16), .B0(n29), .Y(data_o[9]) );
  AO21X4 U70 ( .A0(data0_i[11]), .A1(n16), .B0(n31), .Y(data_o[11]) );
  AO21X4 U71 ( .A0(data0_i[12]), .A1(n16), .B0(n32), .Y(data_o[12]) );
  AO21X4 U72 ( .A0(data0_i[14]), .A1(n16), .B0(n34), .Y(data_o[14]) );
  AO22X4 U73 ( .A0(data2_i[19]), .A1(n10), .B0(data1_i[19]), .B1(n2), .Y(n39)
         );
  AO21X4 U74 ( .A0(data0_i[19]), .A1(n16), .B0(n39), .Y(data_o[19]) );
  AO21X4 U75 ( .A0(data0_i[20]), .A1(n16), .B0(n40), .Y(data_o[20]) );
  AO21X4 U76 ( .A0(data0_i[21]), .A1(n16), .B0(n41), .Y(data_o[21]) );
  AO21X4 U77 ( .A0(data0_i[26]), .A1(n16), .B0(n44), .Y(data_o[26]) );
  AO21X4 U78 ( .A0(data0_i[28]), .A1(n16), .B0(n46), .Y(data_o[28]) );
  AO21X4 U79 ( .A0(data0_i[29]), .A1(n16), .B0(n47), .Y(data_o[29]) );
  AO22X4 U80 ( .A0(data2_i[31]), .A1(n10), .B0(data1_i[31]), .B1(n2), .Y(n48)
         );
  AO21X4 U81 ( .A0(data0_i[31]), .A1(n16), .B0(n48), .Y(data_o[31]) );
endmodule


module MUX_32_3to1_1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  AO21X2 U2 ( .A0(data0_i[21]), .A1(n8), .B0(n39), .Y(data_o[21]) );
  AND2X4 U3 ( .A(select_i[0]), .B(n26), .Y(n15) );
  INVX4 U4 ( .A(select_i[0]), .Y(n25) );
  BUFX12 U5 ( .A(n13), .Y(n8) );
  AND2X2 U6 ( .A(n26), .B(n25), .Y(n13) );
  AO21X2 U7 ( .A0(data0_i[31]), .A1(n8), .B0(n48), .Y(data_o[31]) );
  AO21X2 U8 ( .A0(data0_i[30]), .A1(n8), .B0(n47), .Y(data_o[30]) );
  AO21X1 U9 ( .A0(data0_i[29]), .A1(n8), .B0(n46), .Y(data_o[29]) );
  AO21X2 U10 ( .A0(data0_i[28]), .A1(n8), .B0(n45), .Y(data_o[28]) );
  AO21X2 U11 ( .A0(data0_i[25]), .A1(n8), .B0(n42), .Y(data_o[25]) );
  AO21X2 U12 ( .A0(data0_i[24]), .A1(n8), .B0(n41), .Y(data_o[24]) );
  NAND2X1 U13 ( .A(n4), .B(n1), .Y(data_o[23]) );
  AO21X1 U14 ( .A0(data0_i[22]), .A1(n8), .B0(n40), .Y(data_o[22]) );
  AO22X2 U15 ( .A0(data2_i[22]), .A1(n11), .B0(data1_i[22]), .B1(n5), .Y(n40)
         );
  AO21X1 U16 ( .A0(data0_i[20]), .A1(n8), .B0(n38), .Y(data_o[20]) );
  AOI22X1 U17 ( .A0(data2_i[18]), .A1(n12), .B0(data1_i[18]), .B1(n5), .Y(n17)
         );
  AO22X1 U18 ( .A0(data2_i[14]), .A1(n12), .B0(data1_i[14]), .B1(n5), .Y(n33)
         );
  AO21X2 U19 ( .A0(data0_i[12]), .A1(n8), .B0(n31), .Y(data_o[12]) );
  OAI2BB1X1 U20 ( .A0N(data0_i[11]), .A1N(n8), .B0(n16), .Y(data_o[11]) );
  AOI22X1 U21 ( .A0(data2_i[11]), .A1(n12), .B0(data1_i[11]), .B1(n5), .Y(n16)
         );
  AO21X2 U22 ( .A0(data0_i[10]), .A1(n8), .B0(n30), .Y(data_o[10]) );
  AO21X2 U23 ( .A0(data0_i[8]), .A1(n8), .B0(n29), .Y(data_o[8]) );
  OAI2BB1X2 U24 ( .A0N(data0_i[7]), .A1N(n8), .B0(n22), .Y(data_o[7]) );
  OAI2BB1X1 U25 ( .A0N(data0_i[6]), .A1N(n8), .B0(n21), .Y(data_o[6]) );
  AOI22X1 U26 ( .A0(data2_i[6]), .A1(n10), .B0(data1_i[6]), .B1(n6), .Y(n21)
         );
  AO21X2 U27 ( .A0(data0_i[4]), .A1(n8), .B0(n28), .Y(data_o[4]) );
  OAI2BB1X2 U28 ( .A0N(data0_i[3]), .A1N(n8), .B0(n18), .Y(data_o[3]) );
  CLKAND2X3 U29 ( .A(n2), .B(n3), .Y(n18) );
  NAND2X2 U30 ( .A(data2_i[3]), .B(n11), .Y(n2) );
  OAI2BB1X2 U31 ( .A0N(data0_i[2]), .A1N(n8), .B0(n20), .Y(data_o[2]) );
  AOI22X1 U32 ( .A0(data2_i[23]), .A1(n12), .B0(data1_i[23]), .B1(n6), .Y(n1)
         );
  CLKAND2X2 U33 ( .A(select_i[1]), .B(n25), .Y(n14) );
  AO22X4 U34 ( .A0(data2_i[10]), .A1(n10), .B0(data1_i[10]), .B1(n5), .Y(n30)
         );
  AO22X4 U35 ( .A0(data2_i[0]), .A1(n10), .B0(data1_i[0]), .B1(n6), .Y(n27) );
  AOI22X2 U36 ( .A0(data2_i[2]), .A1(n12), .B0(data1_i[2]), .B1(n6), .Y(n20)
         );
  AO22X2 U37 ( .A0(data2_i[29]), .A1(n12), .B0(data1_i[29]), .B1(n5), .Y(n46)
         );
  AO22X4 U38 ( .A0(data2_i[25]), .A1(n12), .B0(data1_i[25]), .B1(n5), .Y(n42)
         );
  INVX12 U39 ( .A(n9), .Y(n12) );
  AO21X4 U40 ( .A0(data0_i[0]), .A1(n8), .B0(n27), .Y(data_o[0]) );
  OAI2BB1X2 U41 ( .A0N(data0_i[1]), .A1N(n8), .B0(n23), .Y(data_o[1]) );
  AO22X1 U42 ( .A0(data2_i[8]), .A1(n12), .B0(data1_i[8]), .B1(n5), .Y(n29) );
  AOI22X2 U43 ( .A0(data2_i[5]), .A1(n12), .B0(data1_i[5]), .B1(n5), .Y(n24)
         );
  OAI2BB1X4 U44 ( .A0N(data0_i[5]), .A1N(n8), .B0(n24), .Y(data_o[5]) );
  INVX1 U45 ( .A(select_i[1]), .Y(n26) );
  AO22X4 U46 ( .A0(data2_i[13]), .A1(n11), .B0(data1_i[13]), .B1(n6), .Y(n32)
         );
  INVX20 U47 ( .A(n9), .Y(n11) );
  AO21X4 U48 ( .A0(data0_i[15]), .A1(n8), .B0(n34), .Y(data_o[15]) );
  NAND2X1 U49 ( .A(data1_i[3]), .B(n6), .Y(n3) );
  BUFX12 U50 ( .A(n15), .Y(n6) );
  NAND2X1 U51 ( .A(data0_i[23]), .B(n8), .Y(n4) );
  AO21X4 U52 ( .A0(data0_i[27]), .A1(n8), .B0(n44), .Y(data_o[27]) );
  OAI2BB1X2 U53 ( .A0N(data0_i[18]), .A1N(n8), .B0(n17), .Y(data_o[18]) );
  CLKBUFX12 U54 ( .A(n15), .Y(n5) );
  BUFX8 U55 ( .A(n14), .Y(n7) );
  AO21X2 U56 ( .A0(data0_i[19]), .A1(n8), .B0(n37), .Y(data_o[19]) );
  CLKINVX12 U57 ( .A(n7), .Y(n9) );
  INVX20 U58 ( .A(n9), .Y(n10) );
  AO21X4 U59 ( .A0(data0_i[13]), .A1(n8), .B0(n32), .Y(data_o[13]) );
  AO21X4 U60 ( .A0(data0_i[14]), .A1(n8), .B0(n33), .Y(data_o[14]) );
  AO21X4 U61 ( .A0(data0_i[17]), .A1(n8), .B0(n36), .Y(data_o[17]) );
  AO21X4 U62 ( .A0(data0_i[26]), .A1(n8), .B0(n43), .Y(data_o[26]) );
  AO21X4 U63 ( .A0(data0_i[16]), .A1(n8), .B0(n35), .Y(data_o[16]) );
  OAI2BB1X1 U64 ( .A0N(data0_i[9]), .A1N(n8), .B0(n19), .Y(data_o[9]) );
  AOI22X1 U65 ( .A0(data2_i[9]), .A1(n11), .B0(data1_i[9]), .B1(n5), .Y(n19)
         );
  AOI22X1 U66 ( .A0(data2_i[7]), .A1(n11), .B0(data1_i[7]), .B1(n6), .Y(n22)
         );
  AO22X1 U67 ( .A0(data2_i[27]), .A1(n10), .B0(data1_i[27]), .B1(n6), .Y(n44)
         );
  AO22X1 U68 ( .A0(data2_i[24]), .A1(n10), .B0(data1_i[24]), .B1(n6), .Y(n41)
         );
  AOI22X1 U69 ( .A0(data2_i[1]), .A1(n10), .B0(data1_i[1]), .B1(n6), .Y(n23)
         );
  AO22X1 U70 ( .A0(data2_i[4]), .A1(n11), .B0(data1_i[4]), .B1(n5), .Y(n28) );
  AO22XL U71 ( .A0(data2_i[15]), .A1(n10), .B0(data1_i[15]), .B1(n5), .Y(n34)
         );
  AO22X1 U72 ( .A0(data2_i[19]), .A1(n10), .B0(data1_i[19]), .B1(n6), .Y(n37)
         );
  AO22X1 U73 ( .A0(data2_i[12]), .A1(n11), .B0(data1_i[12]), .B1(n5), .Y(n31)
         );
  AO22XL U74 ( .A0(data2_i[28]), .A1(n11), .B0(data1_i[28]), .B1(n6), .Y(n45)
         );
  AO22X1 U75 ( .A0(data2_i[16]), .A1(n11), .B0(data1_i[16]), .B1(n6), .Y(n35)
         );
  AO22X1 U76 ( .A0(data2_i[20]), .A1(n10), .B0(data1_i[20]), .B1(n5), .Y(n38)
         );
  AO22XL U77 ( .A0(data2_i[31]), .A1(n12), .B0(data1_i[31]), .B1(n5), .Y(n48)
         );
  AO22XL U78 ( .A0(data2_i[21]), .A1(n10), .B0(data1_i[21]), .B1(n6), .Y(n39)
         );
  AO22XL U79 ( .A0(data2_i[30]), .A1(n11), .B0(data1_i[30]), .B1(n6), .Y(n47)
         );
  AO22XL U80 ( .A0(data2_i[17]), .A1(n10), .B0(data1_i[17]), .B1(n5), .Y(n36)
         );
  AO22XL U81 ( .A0(data2_i[26]), .A1(n11), .B0(data1_i[26]), .B1(n6), .Y(n43)
         );
endmodule


module forwarding ( Rs_regD, Rt_regD, RegWrite_regE, wsel_regE, RegWrite_regM, 
        wsel_regM, FU_Asel, FU_Bsel );
  input [4:0] Rs_regD;
  input [4:0] Rt_regD;
  input [4:0] wsel_regE;
  input [4:0] wsel_regM;
  output [1:0] FU_Asel;
  output [1:0] FU_Bsel;
  input RegWrite_regE, RegWrite_regM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  CLKXOR2X4 U2 ( .A(n26), .B(Rs_regD[4]), .Y(n37) );
  CLKXOR2X4 U3 ( .A(n27), .B(Rs_regD[3]), .Y(n36) );
  INVX4 U4 ( .A(wsel_regE[3]), .Y(n27) );
  INVX4 U5 ( .A(wsel_regE[4]), .Y(n26) );
  NOR4X6 U6 ( .A(n42), .B(n41), .C(n40), .D(n39), .Y(FU_Asel[0]) );
  INVX3 U7 ( .A(wsel_regM[0]), .Y(n20) );
  INVX3 U8 ( .A(wsel_regM[3]), .Y(n19) );
  INVX3 U9 ( .A(wsel_regM[1]), .Y(n18) );
  XOR2X1 U10 ( .A(n28), .B(Rs_regD[0]), .Y(n33) );
  XOR2X1 U11 ( .A(n20), .B(Rt_regD[0]), .Y(n3) );
  XOR2X1 U12 ( .A(n18), .B(Rt_regD[1]), .Y(n5) );
  CLKXOR2X2 U13 ( .A(n19), .B(Rs_regD[3]), .Y(n24) );
  XOR2X1 U14 ( .A(n20), .B(Rs_regD[0]), .Y(n23) );
  AND4X4 U15 ( .A(n14), .B(n13), .C(n35), .D(n12), .Y(FU_Bsel[1]) );
  XOR2X1 U16 ( .A(n26), .B(Rt_regD[4]), .Y(n14) );
  XOR2X1 U17 ( .A(n27), .B(Rt_regD[3]), .Y(n13) );
  XOR2X1 U18 ( .A(n19), .B(Rt_regD[3]), .Y(n4) );
  XOR2X1 U19 ( .A(n30), .B(Rs_regD[1]), .Y(n31) );
  CLKINVX4 U20 ( .A(wsel_regE[1]), .Y(n30) );
  NOR4X8 U21 ( .A(n17), .B(n16), .C(FU_Bsel[1]), .D(n15), .Y(FU_Bsel[0]) );
  XOR2X1 U22 ( .A(n29), .B(Rt_regD[2]), .Y(n10) );
  NAND3BX4 U23 ( .AN(wsel_regE[1]), .B(n28), .C(n29), .Y(n7) );
  XOR2X2 U24 ( .A(n28), .B(Rt_regD[0]), .Y(n11) );
  XOR2X1 U25 ( .A(n30), .B(Rt_regD[1]), .Y(n9) );
  NAND2X2 U26 ( .A(RegWrite_regM), .B(n38), .Y(n16) );
  NAND3BX2 U27 ( .AN(wsel_regM[4]), .B(n19), .C(n6), .Y(n38) );
  INVX6 U28 ( .A(n43), .Y(FU_Asel[1]) );
  NAND4X8 U29 ( .A(n37), .B(n36), .C(n35), .D(n34), .Y(n43) );
  OAI31X2 U30 ( .A0(n7), .A1(wsel_regE[4]), .A2(wsel_regE[3]), .B0(
        RegWrite_regE), .Y(n8) );
  AND3X6 U31 ( .A(n33), .B(n32), .C(n31), .Y(n34) );
  XOR2X1 U32 ( .A(n21), .B(Rt_regD[2]), .Y(n2) );
  NAND4X2 U33 ( .A(n5), .B(n4), .C(n3), .D(n2), .Y(n17) );
  INVX2 U34 ( .A(n38), .Y(n40) );
  INVX4 U35 ( .A(n8), .Y(n35) );
  CLKINVX8 U36 ( .A(wsel_regE[2]), .Y(n29) );
  CLKINVX8 U37 ( .A(wsel_regE[0]), .Y(n28) );
  XOR2X1 U38 ( .A(n21), .B(Rs_regD[2]), .Y(n22) );
  XOR2X1 U39 ( .A(n18), .B(Rs_regD[1]), .Y(n25) );
  NAND2X6 U40 ( .A(RegWrite_regM), .B(n43), .Y(n41) );
  XOR2X1 U41 ( .A(n29), .B(Rs_regD[2]), .Y(n32) );
  INVX3 U42 ( .A(wsel_regM[2]), .Y(n21) );
  AND3X4 U43 ( .A(n20), .B(n18), .C(n21), .Y(n6) );
  AND3X4 U44 ( .A(n11), .B(n10), .C(n9), .Y(n12) );
  XOR2X2 U45 ( .A(Rt_regD[4]), .B(wsel_regM[4]), .Y(n15) );
  NAND4X2 U46 ( .A(n25), .B(n24), .C(n23), .D(n22), .Y(n42) );
  XOR2X2 U47 ( .A(Rs_regD[4]), .B(wsel_regM[4]), .Y(n39) );
endmodule


module hazard_detection ( Branch_EX, equal, branchpred_his, JumpReg_regD, 
        MemRead_regD, Rt_regD, Rs, Rt, ICACHE_stall, DCACHE_stall, 
        stall_lw_use, stallcache, flush, pred_cond );
  input [4:0] Rt_regD;
  input [4:0] Rs;
  input [4:0] Rt;
  input Branch_EX, equal, branchpred_his, JumpReg_regD, MemRead_regD,
         ICACHE_stall, DCACHE_stall;
  output stall_lw_use, stallcache, flush, pred_cond;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;

  NOR2X2 U2 ( .A(n20), .B(JumpReg_regD), .Y(stall_lw_use) );
  OR2X8 U3 ( .A(DCACHE_stall), .B(ICACHE_stall), .Y(stallcache) );
  XOR2XL U4 ( .A(Rt[4]), .B(Rt_regD[4]), .Y(n13) );
  XOR2XL U5 ( .A(Rt[1]), .B(Rt_regD[1]), .Y(n14) );
  XOR2XL U6 ( .A(Rs[1]), .B(Rt_regD[1]), .Y(n17) );
  XOR2XL U7 ( .A(Rs[4]), .B(Rt_regD[4]), .Y(n16) );
  INVXL U8 ( .A(Rt_regD[3]), .Y(n9) );
  INVXL U9 ( .A(Rt_regD[2]), .Y(n8) );
  CLKINVX1 U10 ( .A(Branch_EX), .Y(n2) );
  NAND2X1 U11 ( .A(MemRead_regD), .B(n19), .Y(n20) );
  OAI33X1 U12 ( .A0(n18), .A1(n17), .A2(n16), .B0(n15), .B1(n14), .B2(n13), 
        .Y(n19) );
  NAND3BX1 U13 ( .AN(n12), .B(n11), .C(n10), .Y(n15) );
  XOR2X1 U14 ( .A(n8), .B(Rt[2]), .Y(n11) );
  XOR2X1 U15 ( .A(Rt[0]), .B(Rt_regD[0]), .Y(n12) );
  XOR2X1 U16 ( .A(n9), .B(Rt[3]), .Y(n10) );
  NAND3BX1 U17 ( .AN(n7), .B(n6), .C(n5), .Y(n18) );
  XOR2X1 U18 ( .A(n8), .B(Rs[2]), .Y(n6) );
  XOR2X1 U19 ( .A(Rs[0]), .B(Rt_regD[0]), .Y(n7) );
  XOR2X1 U20 ( .A(n9), .B(Rs[3]), .Y(n5) );
  NOR2X8 U21 ( .A(n3), .B(n2), .Y(pred_cond) );
  XNOR2X4 U22 ( .A(branchpred_his), .B(equal), .Y(n3) );
  INVXL U23 ( .A(pred_cond), .Y(n4) );
  NAND3BXL U24 ( .AN(JumpReg_regD), .B(n20), .C(n4), .Y(flush) );
endmodule


module branch_prediction ( clk, rst_n, branch, equal, predict, branchpred_his
 );
  input clk, rst_n, branch, equal;
  output predict, branchpred_his;
  wire   n9, n10, n1, n2, n3, n4, n5;
  wire   [1:0] state;

  DFFRX1 branchpred_reg_reg ( .D(predict), .CK(clk), .RN(rst_n), .Q(
        branchpred_his) );
  DFFRX1 \state_reg[1]  ( .D(n9), .CK(clk), .RN(rst_n), .Q(state[1]), .QN(
        predict) );
  DFFSX1 \state_reg[0]  ( .D(n10), .CK(clk), .SN(rst_n), .Q(state[0]), .QN(n5)
         );
  OAI2BB2XL U3 ( .B0(state[0]), .B1(equal), .A0N(state[1]), .A1N(n5), .Y(n1)
         );
  INVXL U4 ( .A(branch), .Y(n4) );
  OAI2BB2XL U5 ( .B0(n2), .B1(n5), .A0N(branch), .A1N(n1), .Y(n10) );
  OAI32XL U6 ( .A0(equal), .A1(n5), .A2(n4), .B0(n3), .B1(predict), .Y(n9) );
  AND3X2 U7 ( .A(equal), .B(branch), .C(n5), .Y(n3) );
  AOI2BB1XL U8 ( .A0N(equal), .A1N(predict), .B0(n4), .Y(n2) );
endmodule


module precontrolDec ( instruction_next, Jump_IF, Branch_IF );
  input [31:0] instruction_next;
  output Jump_IF, Branch_IF;
  wire   n1, n2, n3, n4;

  OR3X6 U1 ( .A(instruction_next[30]), .B(instruction_next[29]), .C(
        instruction_next[31]), .Y(n2) );
  CLKINVX4 U2 ( .A(n2), .Y(n4) );
  OR2X2 U3 ( .A(instruction_next[26]), .B(instruction_next[27]), .Y(n1) );
  NOR3X6 U4 ( .A(n3), .B(n1), .C(n2), .Y(Branch_IF) );
  AND3X8 U5 ( .A(n4), .B(instruction_next[27]), .C(n3), .Y(Jump_IF) );
  INVX3 U6 ( .A(instruction_next[28]), .Y(n3) );
endmodule


module nextPCcalculator_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n21, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n40, n41, n44, n45, n47, n48, n49, n51, n52, n53, n55,
         n56, n57, n58, n59, n62, n63, n67, n68, n70, n71, n73, n74, n75, n78,
         n79, n81, n85, n86, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n104, n105, n106, n107, n108, n109, n111, n114, n115,
         n116, n118, n120, n121, n122, n123, n124, n125, n126, n127, n130,
         n131, n132, n133, n134, n135, n136, n138, n139, n140, n141, n142,
         n143, n144, n145, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n169, n171,
         n172, n174, n177, n178, n179, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n198,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n315, n316, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354;
  assign n21 = A[30];
  assign n27 = A[29];
  assign n37 = A[27];
  assign n41 = A[26];
  assign n49 = A[25];
  assign n53 = A[24];
  assign n59 = A[23];
  assign n63 = A[22];
  assign n71 = A[21];
  assign n75 = A[20];
  assign n81 = A[19];
  assign n85 = A[18];

  OAI21X4 U179 ( .A0(n185), .A1(n157), .B0(n158), .Y(n156) );
  AOI21X4 U220 ( .A0(n194), .A1(n186), .B0(n187), .Y(n185) );
  NAND2X2 U248 ( .A(n319), .B(A[31]), .Y(n322) );
  OAI21X2 U249 ( .A0(n193), .A1(n191), .B0(n192), .Y(n190) );
  NOR2X6 U250 ( .A(n121), .B(n114), .Y(n108) );
  INVX1 U251 ( .A(n121), .Y(n202) );
  OAI21X2 U252 ( .A0(n155), .A1(n153), .B0(n154), .Y(n152) );
  NAND2X2 U253 ( .A(n45), .B(n41), .Y(n40) );
  CLKINVX8 U254 ( .A(n44), .Y(n45) );
  INVX6 U255 ( .A(n156), .Y(n155) );
  BUFX8 U256 ( .A(B[17]), .Y(n339) );
  NAND2X2 U257 ( .A(B[13]), .B(A[13]), .Y(n133) );
  NAND2XL U258 ( .A(n208), .B(n169), .Y(n11) );
  NAND2X1 U259 ( .A(n324), .B(n169), .Y(n165) );
  OAI21X4 U260 ( .A0(n188), .A1(n192), .B0(n189), .Y(n187) );
  INVXL U261 ( .A(n166), .Y(n208) );
  OR2X1 U262 ( .A(n174), .B(n166), .Y(n324) );
  NOR2BX1 U263 ( .AN(n315), .B(n166), .Y(n164) );
  NOR2X6 U264 ( .A(n166), .B(n161), .Y(n159) );
  NOR2X4 U265 ( .A(n191), .B(n188), .Y(n186) );
  INVXL U266 ( .A(n188), .Y(n211) );
  NOR2X6 U267 ( .A(B[5]), .B(A[5]), .Y(n188) );
  INVX3 U268 ( .A(n125), .Y(n127) );
  NAND2X6 U269 ( .A(n345), .B(n118), .Y(n116) );
  NAND2X6 U270 ( .A(n344), .B(n318), .Y(n345) );
  CLKAND2X12 U271 ( .A(n127), .B(n202), .Y(n323) );
  OR2X8 U272 ( .A(n325), .B(n127), .Y(n123) );
  AOI21X4 U273 ( .A0(n127), .A1(n99), .B0(n100), .Y(n98) );
  NOR2X2 U274 ( .A(n1), .B(n24), .Y(n23) );
  INVX1 U275 ( .A(n25), .Y(n24) );
  NOR2X4 U276 ( .A(n1), .B(n30), .Y(n29) );
  CLKINVX12 U277 ( .A(n346), .Y(n1) );
  AND2X8 U278 ( .A(n109), .B(n92), .Y(n326) );
  NAND2X6 U279 ( .A(B[16]), .B(A[16]), .Y(n104) );
  INVXL U280 ( .A(n101), .Y(n200) );
  NOR2BX2 U281 ( .AN(n108), .B(n101), .Y(n99) );
  NOR2X6 U282 ( .A(B[16]), .B(A[16]), .Y(n101) );
  NOR2X8 U283 ( .A(B[15]), .B(A[15]), .Y(n114) );
  INVXL U284 ( .A(n114), .Y(n201) );
  NAND2X6 U285 ( .A(n315), .B(n159), .Y(n157) );
  AOI21X4 U286 ( .A0(n172), .A1(n159), .B0(n160), .Y(n158) );
  NAND2XL U287 ( .A(n200), .B(n104), .Y(n3) );
  INVX4 U288 ( .A(n104), .Y(n342) );
  INVX4 U289 ( .A(n172), .Y(n174) );
  AO21X4 U290 ( .A0(n184), .A1(n315), .B0(n172), .Y(n348) );
  OAI21X4 U291 ( .A0(n177), .A1(n183), .B0(n178), .Y(n172) );
  BUFX6 U292 ( .A(n171), .Y(n315) );
  NOR2X6 U293 ( .A(B[7]), .B(A[7]), .Y(n177) );
  NAND2X4 U294 ( .A(B[9]), .B(A[9]), .Y(n162) );
  NAND2X4 U295 ( .A(n108), .B(n92), .Y(n90) );
  NOR2X4 U296 ( .A(n101), .B(n94), .Y(n92) );
  OAI21X2 U297 ( .A0(n161), .A1(n169), .B0(n162), .Y(n160) );
  NOR2X4 U298 ( .A(B[9]), .B(A[9]), .Y(n161) );
  NOR2X4 U299 ( .A(B[3]), .B(A[3]), .Y(n195) );
  NAND2X4 U300 ( .A(n41), .B(n37), .Y(n36) );
  NOR2X4 U301 ( .A(B[11]), .B(A[11]), .Y(n150) );
  NAND2X4 U302 ( .A(n331), .B(n332), .Y(SUM[27]) );
  NAND2X2 U303 ( .A(n329), .B(n330), .Y(n332) );
  NAND2X4 U304 ( .A(n321), .B(n322), .Y(SUM[31]) );
  INVX3 U305 ( .A(n191), .Y(n212) );
  NOR2X4 U306 ( .A(n139), .B(n132), .Y(n130) );
  NOR2X4 U307 ( .A(n153), .B(n150), .Y(n144) );
  NAND2X2 U308 ( .A(B[7]), .B(A[7]), .Y(n178) );
  NOR2X4 U309 ( .A(B[8]), .B(A[8]), .Y(n166) );
  NOR2X2 U310 ( .A(n182), .B(n177), .Y(n171) );
  NAND2X2 U311 ( .A(B[8]), .B(A[8]), .Y(n169) );
  CLKINVX1 U312 ( .A(n349), .Y(n329) );
  INVX3 U313 ( .A(n29), .Y(n334) );
  NOR2X4 U314 ( .A(n323), .B(n120), .Y(n118) );
  INVX3 U315 ( .A(n155), .Y(n344) );
  NAND2X2 U316 ( .A(B[15]), .B(A[15]), .Y(n115) );
  NOR2X2 U317 ( .A(n58), .B(n48), .Y(n47) );
  NAND2X2 U318 ( .A(n53), .B(n49), .Y(n48) );
  NAND2X1 U319 ( .A(n99), .B(n126), .Y(n97) );
  NAND2X2 U320 ( .A(B[12]), .B(A[12]), .Y(n140) );
  OR2X6 U321 ( .A(n327), .B(n328), .Y(n145) );
  CLKBUFX3 U322 ( .A(n133), .Y(n340) );
  XNOR2X1 U323 ( .A(n190), .B(n14), .Y(SUM[5]) );
  NAND2X1 U324 ( .A(n211), .B(n189), .Y(n14) );
  NAND2X1 U325 ( .A(n213), .B(n196), .Y(n16) );
  CLKINVX1 U326 ( .A(n195), .Y(n213) );
  BUFX6 U327 ( .A(n123), .Y(n338) );
  NAND2X1 U328 ( .A(n206), .B(n154), .Y(n9) );
  XNOR2X2 U329 ( .A(n152), .B(n8), .Y(SUM[11]) );
  XNOR2X1 U330 ( .A(n184), .B(n13), .Y(SUM[6]) );
  INVX3 U331 ( .A(n94), .Y(n341) );
  OR2X1 U332 ( .A(B[2]), .B(A[2]), .Y(n316) );
  AND2X2 U333 ( .A(n316), .B(n198), .Y(SUM[2]) );
  AND2X2 U334 ( .A(n126), .B(n202), .Y(n318) );
  NOR2X6 U335 ( .A(n1), .B(n20), .Y(n19) );
  NAND2X6 U336 ( .A(n333), .B(n107), .Y(n105) );
  AOI21X2 U337 ( .A0(n127), .A1(n108), .B0(n109), .Y(n107) );
  OR2X6 U338 ( .A(n1), .B(n78), .Y(n353) );
  XOR2X1 U339 ( .A(n155), .B(n9), .Y(SUM[10]) );
  NOR2X4 U340 ( .A(n155), .B(n124), .Y(n325) );
  NOR2X4 U341 ( .A(n1), .B(n74), .Y(n73) );
  XOR2X4 U342 ( .A(n73), .B(n71), .Y(SUM[21]) );
  OR2X4 U343 ( .A(n155), .B(n106), .Y(n333) );
  NAND2X1 U344 ( .A(n126), .B(n108), .Y(n106) );
  OR2X6 U345 ( .A(n1), .B(n86), .Y(n354) );
  OAI21X2 U346 ( .A0(n155), .A1(n135), .B0(n136), .Y(n134) );
  OAI21X2 U347 ( .A0(n155), .A1(n142), .B0(n143), .Y(n141) );
  XOR2X4 U348 ( .A(n51), .B(n49), .Y(SUM[25]) );
  NOR2X4 U349 ( .A(n1), .B(n52), .Y(n51) );
  NAND2X1 U350 ( .A(n144), .B(n204), .Y(n135) );
  XNOR2X4 U351 ( .A(n338), .B(n5), .Y(SUM[14]) );
  OAI21X1 U352 ( .A0(n111), .A1(n101), .B0(n104), .Y(n100) );
  NOR2X6 U353 ( .A(n44), .B(n26), .Y(n25) );
  NAND2X4 U354 ( .A(n31), .B(n27), .Y(n26) );
  XOR2X4 U355 ( .A(n23), .B(n21), .Y(SUM[30]) );
  OAI2BB1X4 U356 ( .A0N(n156), .A1N(n88), .B0(n347), .Y(n346) );
  NOR2X2 U357 ( .A(n1), .B(n34), .Y(n33) );
  OR2X6 U358 ( .A(n1), .B(n68), .Y(n352) );
  XNOR2X4 U359 ( .A(n353), .B(n75), .Y(SUM[20]) );
  OR2X6 U360 ( .A(n1), .B(n62), .Y(n350) );
  XNOR2X4 U361 ( .A(n351), .B(n41), .Y(SUM[26]) );
  OR2X4 U362 ( .A(n1), .B(n44), .Y(n351) );
  NOR2X2 U363 ( .A(n326), .B(n93), .Y(n91) );
  NAND2X2 U364 ( .A(n343), .B(n95), .Y(n93) );
  NAND2X2 U365 ( .A(n341), .B(n342), .Y(n343) );
  NOR2X4 U366 ( .A(n1), .B(n56), .Y(n55) );
  INVX6 U367 ( .A(n124), .Y(n126) );
  NAND2X4 U368 ( .A(B[3]), .B(A[3]), .Y(n196) );
  NAND2X4 U369 ( .A(n25), .B(n21), .Y(n20) );
  NOR2X8 U370 ( .A(B[4]), .B(A[4]), .Y(n191) );
  OR2X8 U371 ( .A(n1), .B(n40), .Y(n349) );
  NOR2X2 U372 ( .A(n124), .B(n90), .Y(n88) );
  NOR2X6 U373 ( .A(n339), .B(A[17]), .Y(n94) );
  NAND2X1 U374 ( .A(n45), .B(n31), .Y(n30) );
  NAND2X2 U375 ( .A(n19), .B(n320), .Y(n321) );
  INVX3 U376 ( .A(n19), .Y(n319) );
  CLKINVX1 U377 ( .A(A[31]), .Y(n320) );
  XOR2X2 U378 ( .A(n1), .B(n86), .Y(SUM[18]) );
  XNOR2X4 U379 ( .A(n350), .B(n59), .Y(SUM[23]) );
  AOI21X2 U380 ( .A0(n184), .A1(n164), .B0(n165), .Y(n163) );
  XNOR2X2 U381 ( .A(n33), .B(n32), .Y(SUM[28]) );
  OA21X4 U382 ( .A0(n125), .A1(n90), .B0(n91), .Y(n347) );
  NOR2X6 U383 ( .A(n150), .B(n154), .Y(n327) );
  CLKINVX2 U384 ( .A(n151), .Y(n328) );
  NAND2X8 U385 ( .A(B[10]), .B(A[10]), .Y(n154) );
  NAND2X4 U386 ( .A(B[11]), .B(A[11]), .Y(n151) );
  AOI21X1 U387 ( .A0(n145), .A1(n204), .B0(n138), .Y(n136) );
  INVX3 U388 ( .A(n145), .Y(n143) );
  NAND2X2 U389 ( .A(n349), .B(n37), .Y(n331) );
  INVX1 U390 ( .A(n37), .Y(n330) );
  XNOR2X4 U391 ( .A(n105), .B(n3), .Y(SUM[16]) );
  NAND2X2 U392 ( .A(n29), .B(n335), .Y(n336) );
  NAND2X4 U393 ( .A(n334), .B(n27), .Y(n337) );
  NAND2X4 U394 ( .A(n336), .B(n337), .Y(SUM[29]) );
  INVXL U395 ( .A(n27), .Y(n335) );
  OAI21X4 U396 ( .A0(n132), .A1(n140), .B0(n340), .Y(n131) );
  INVX3 U397 ( .A(n132), .Y(n203) );
  NOR2X4 U398 ( .A(B[13]), .B(A[13]), .Y(n132) );
  INVX4 U399 ( .A(n109), .Y(n111) );
  OAI21X4 U400 ( .A0(n114), .A1(n122), .B0(n115), .Y(n109) );
  NAND2X2 U401 ( .A(B[5]), .B(A[5]), .Y(n189) );
  XNOR2X4 U402 ( .A(n348), .B(n11), .Y(SUM[8]) );
  XNOR2X2 U403 ( .A(n141), .B(n7), .Y(SUM[12]) );
  XNOR2X2 U404 ( .A(n134), .B(n6), .Y(SUM[13]) );
  INVX2 U405 ( .A(n185), .Y(n184) );
  XNOR2X4 U406 ( .A(n96), .B(n2), .Y(SUM[17]) );
  XNOR2X4 U407 ( .A(n354), .B(n81), .Y(SUM[19]) );
  INVXL U408 ( .A(n194), .Y(n193) );
  XNOR2X4 U409 ( .A(n352), .B(n63), .Y(SUM[22]) );
  XOR2X2 U410 ( .A(n55), .B(n53), .Y(SUM[24]) );
  AOI21X4 U411 ( .A0(n145), .A1(n130), .B0(n131), .Y(n125) );
  NAND2X4 U412 ( .A(n144), .B(n130), .Y(n124) );
  XNOR2X4 U413 ( .A(n116), .B(n4), .Y(SUM[15]) );
  NOR2X2 U414 ( .A(B[12]), .B(A[12]), .Y(n139) );
  INVXL U415 ( .A(n144), .Y(n142) );
  NOR2X4 U416 ( .A(B[10]), .B(A[10]), .Y(n153) );
  OAI21X2 U417 ( .A0(n155), .A1(n97), .B0(n98), .Y(n96) );
  NAND2X4 U418 ( .A(n67), .B(n47), .Y(n44) );
  INVXL U419 ( .A(n122), .Y(n120) );
  NAND2X2 U420 ( .A(n63), .B(n59), .Y(n58) );
  INVX1 U421 ( .A(n57), .Y(n56) );
  NAND2X1 U422 ( .A(n45), .B(n35), .Y(n34) );
  INVXL U423 ( .A(n36), .Y(n35) );
  NAND2XL U424 ( .A(n79), .B(n75), .Y(n74) );
  NAND2X4 U425 ( .A(B[6]), .B(A[6]), .Y(n183) );
  OAI21X4 U426 ( .A0(n195), .A1(n198), .B0(n196), .Y(n194) );
  NAND2XL U427 ( .A(n341), .B(n95), .Y(n2) );
  NAND2XL U428 ( .A(n203), .B(n340), .Y(n6) );
  NAND2XL U429 ( .A(n204), .B(n140), .Y(n7) );
  INVXL U430 ( .A(n140), .Y(n138) );
  INVXL U431 ( .A(n161), .Y(n207) );
  NAND2XL U432 ( .A(n212), .B(n192), .Y(n15) );
  NAND2XL U433 ( .A(n202), .B(n122), .Y(n5) );
  INVXL U434 ( .A(n182), .Y(n210) );
  INVX3 U435 ( .A(n67), .Y(n68) );
  INVXL U436 ( .A(n78), .Y(n79) );
  NAND2X4 U437 ( .A(B[2]), .B(A[2]), .Y(n198) );
  NOR2X4 U438 ( .A(n32), .B(n36), .Y(n31) );
  INVXL U439 ( .A(n85), .Y(n86) );
  BUFX2 U440 ( .A(A[1]), .Y(SUM[1]) );
  BUFX2 U441 ( .A(A[0]), .Y(SUM[0]) );
  NAND2X1 U442 ( .A(n201), .B(n115), .Y(n4) );
  NAND2X1 U443 ( .A(n205), .B(n151), .Y(n8) );
  CLKINVX1 U444 ( .A(n150), .Y(n205) );
  NAND2X1 U445 ( .A(n210), .B(n183), .Y(n13) );
  XOR2X1 U446 ( .A(n179), .B(n12), .Y(SUM[7]) );
  NAND2X1 U447 ( .A(n209), .B(n178), .Y(n12) );
  AOI21X1 U448 ( .A0(n184), .A1(n210), .B0(n181), .Y(n179) );
  CLKINVX1 U449 ( .A(n177), .Y(n209) );
  NOR2X1 U450 ( .A(n68), .B(n58), .Y(n57) );
  CLKINVX1 U451 ( .A(n153), .Y(n206) );
  CLKINVX1 U452 ( .A(n139), .Y(n204) );
  XOR2X1 U453 ( .A(n16), .B(n198), .Y(SUM[3]) );
  CLKINVX1 U454 ( .A(n183), .Y(n181) );
  XOR2X1 U455 ( .A(n163), .B(n10), .Y(SUM[9]) );
  NAND2X1 U456 ( .A(n207), .B(n162), .Y(n10) );
  XOR2X1 U457 ( .A(n193), .B(n15), .Y(SUM[4]) );
  NOR2X4 U458 ( .A(n78), .B(n70), .Y(n67) );
  NAND2X1 U459 ( .A(n75), .B(n71), .Y(n70) );
  NAND2X1 U460 ( .A(n57), .B(n53), .Y(n52) );
  NAND2X1 U461 ( .A(n67), .B(n63), .Y(n62) );
  NAND2X4 U462 ( .A(B[4]), .B(A[4]), .Y(n192) );
  NOR2X2 U463 ( .A(B[14]), .B(A[14]), .Y(n121) );
  NAND2X4 U464 ( .A(n85), .B(n81), .Y(n78) );
  NAND2X4 U465 ( .A(B[14]), .B(A[14]), .Y(n122) );
  NOR2X2 U466 ( .A(B[6]), .B(A[6]), .Y(n182) );
  NAND2X1 U467 ( .A(n339), .B(A[17]), .Y(n95) );
  INVX3 U468 ( .A(A[28]), .Y(n32) );
endmodule


module nextPCcalculator ( PCcur, PCplus4, PCplus4_regD, targetAddr, 
        branchOffset_I, branchOffset_regD, JumpRegAddr, PCsrc, PCnext );
  input [31:0] PCcur;
  input [31:0] PCplus4;
  input [31:0] PCplus4_regD;
  input [25:0] targetAddr;
  input [15:0] branchOffset_I;
  input [15:0] branchOffset_regD;
  input [31:0] JumpRegAddr;
  input [2:0] PCsrc;
  output [31:0] PCnext;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198;
  wire   [31:0] PCplus4_actual;
  wire   [17:2] branchOffset_actual;
  wire   [31:0] ADDresult;

  nextPCcalculator_DW01_add_1 add_1346 ( .A({PCplus4_actual[31:11], n42, 
        PCplus4_actual[9:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, branchOffset_actual, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(ADDresult) );
  CLKMX2X4 U4 ( .A(PCplus4[27]), .B(PCplus4_regD[27]), .S0(n41), .Y(
        PCplus4_actual[27]) );
  OAI211X2 U5 ( .A0(n52), .A1(n161), .B0(n160), .C0(n159), .Y(PCnext[23]) );
  CLKAND2X3 U6 ( .A(ADDresult[24]), .B(n55), .Y(n17) );
  CLKAND2X8 U7 ( .A(ADDresult[14]), .B(n55), .Y(n6) );
  OAI211X2 U8 ( .A0(n53), .A1(n97), .B0(n96), .C0(n95), .Y(PCnext[7]) );
  OAI211X2 U9 ( .A0(n52), .A1(n173), .B0(n172), .C0(n171), .Y(PCnext[26]) );
  OAI211X2 U10 ( .A0(n53), .A1(n117), .B0(n116), .C0(n115), .Y(PCnext[12]) );
  CLKAND2X3 U11 ( .A(ADDresult[28]), .B(n55), .Y(n20) );
  INVX4 U12 ( .A(n66), .Y(n191) );
  NAND2X1 U13 ( .A(JumpRegAddr[31]), .B(n56), .Y(n25) );
  AOI222X4 U14 ( .A0(JumpRegAddr[6]), .A1(n57), .B0(targetAddr[4]), .B1(n51), 
        .C0(ADDresult[6]), .C1(n55), .Y(n91) );
  OA21X2 U15 ( .A0(n52), .A1(n178), .B0(n177), .Y(n21) );
  AOI222X2 U16 ( .A0(JumpRegAddr[11]), .A1(n56), .B0(targetAddr[9]), .B1(n51), 
        .C0(ADDresult[11]), .C1(n55), .Y(n111) );
  INVX1 U17 ( .A(n64), .Y(n39) );
  CLKMX2X2 U18 ( .A(branchOffset_regD[15]), .B(branchOffset_I[15]), .S0(n64), 
        .Y(branchOffset_actual[17]) );
  MX2X6 U19 ( .A(PCplus4_regD[29]), .B(PCplus4[29]), .S0(n50), .Y(
        PCplus4_actual[29]) );
  MX2X2 U20 ( .A(PCplus4[25]), .B(PCplus4_regD[25]), .S0(n39), .Y(
        PCplus4_actual[25]) );
  NOR3X4 U21 ( .A(n32), .B(n33), .C(n34), .Y(n167) );
  CLKAND2X12 U22 ( .A(ADDresult[25]), .B(n55), .Y(n34) );
  INVX3 U23 ( .A(n180), .Y(n175) );
  BUFX8 U24 ( .A(n175), .Y(n51) );
  BUFX4 U25 ( .A(n194), .Y(n62) );
  OAI211X2 U26 ( .A0(n52), .A1(n133), .B0(n131), .C0(n132), .Y(PCnext[16]) );
  CLKMX2X3 U27 ( .A(branchOffset_regD[5]), .B(branchOffset_I[5]), .S0(n64), 
        .Y(branchOffset_actual[7]) );
  AOI222X2 U28 ( .A0(JumpRegAddr[22]), .A1(n191), .B0(targetAddr[20]), .B1(n51), .C0(ADDresult[22]), .C1(n55), .Y(n155) );
  NAND2X2 U29 ( .A(n28), .B(n167), .Y(PCnext[25]) );
  AOI222X2 U30 ( .A0(JumpRegAddr[20]), .A1(n191), .B0(targetAddr[18]), .B1(
        n175), .C0(ADDresult[20]), .C1(n55), .Y(n147) );
  CLKMX2X3 U31 ( .A(PCplus4_regD[7]), .B(PCplus4[7]), .S0(n64), .Y(
        PCplus4_actual[7]) );
  MX2X2 U32 ( .A(PCplus4_regD[16]), .B(PCplus4[16]), .S0(n64), .Y(
        PCplus4_actual[16]) );
  CLKMX2X3 U33 ( .A(branchOffset_regD[14]), .B(branchOffset_I[14]), .S0(n64), 
        .Y(branchOffset_actual[16]) );
  MX2X2 U34 ( .A(branchOffset_regD[13]), .B(branchOffset_I[13]), .S0(n64), .Y(
        branchOffset_actual[15]) );
  CLKMX2X12 U35 ( .A(PCplus4_regD[15]), .B(PCplus4[15]), .S0(n64), .Y(
        PCplus4_actual[15]) );
  AND2X6 U36 ( .A(PCsrc[2]), .B(n74), .Y(n49) );
  NOR3X8 U37 ( .A(n12), .B(n13), .C(n14), .Y(n159) );
  CLKAND2X12 U38 ( .A(ADDresult[23]), .B(n55), .Y(n14) );
  NAND2X4 U39 ( .A(n21), .B(n176), .Y(PCnext[27]) );
  NOR3X6 U40 ( .A(n29), .B(n30), .C(n31), .Y(n176) );
  OAI211X2 U41 ( .A0(n52), .A1(n149), .B0(n148), .C0(n147), .Y(PCnext[20]) );
  OAI211X2 U42 ( .A0(n53), .A1(n157), .B0(n155), .C0(n156), .Y(PCnext[22]) );
  CLKMX2X8 U43 ( .A(PCplus4_regD[9]), .B(PCplus4[9]), .S0(n64), .Y(
        PCplus4_actual[9]) );
  CLKMX2X8 U44 ( .A(branchOffset_regD[7]), .B(branchOffset_I[7]), .S0(n64), 
        .Y(branchOffset_actual[9]) );
  CLKMX2X3 U45 ( .A(branchOffset_regD[6]), .B(branchOffset_I[6]), .S0(n64), 
        .Y(branchOffset_actual[8]) );
  CLKMX2X2 U46 ( .A(branchOffset_regD[3]), .B(branchOffset_I[3]), .S0(n64), 
        .Y(branchOffset_actual[5]) );
  CLKMX2X2 U47 ( .A(PCplus4_regD[5]), .B(PCplus4[5]), .S0(n64), .Y(
        PCplus4_actual[5]) );
  MX2X2 U48 ( .A(branchOffset_regD[12]), .B(branchOffset_I[12]), .S0(n64), .Y(
        branchOffset_actual[14]) );
  CLKAND2X8 U49 ( .A(ADDresult[29]), .B(n55), .Y(n45) );
  CLKMX2X2 U50 ( .A(PCplus4_regD[8]), .B(PCplus4[8]), .S0(n64), .Y(
        PCplus4_actual[8]) );
  CLKMX2X2 U51 ( .A(PCplus4_regD[18]), .B(PCplus4[18]), .S0(n64), .Y(
        PCplus4_actual[18]) );
  CLKMX2X2 U52 ( .A(PCplus4_regD[17]), .B(PCplus4[17]), .S0(n64), .Y(
        PCplus4_actual[17]) );
  CLKMX2X2 U53 ( .A(PCplus4_regD[12]), .B(PCplus4[12]), .S0(n64), .Y(
        PCplus4_actual[12]) );
  CLKMX2X2 U54 ( .A(branchOffset_regD[10]), .B(branchOffset_I[10]), .S0(n64), 
        .Y(branchOffset_actual[12]) );
  CLKMX2X2 U55 ( .A(branchOffset_regD[11]), .B(branchOffset_I[11]), .S0(n64), 
        .Y(branchOffset_actual[13]) );
  CLKMX2X2 U56 ( .A(PCplus4_regD[13]), .B(PCplus4[13]), .S0(n64), .Y(
        PCplus4_actual[13]) );
  CLKMX2X2 U57 ( .A(PCplus4_regD[30]), .B(PCplus4[30]), .S0(n50), .Y(
        PCplus4_actual[30]) );
  CLKMX2X2 U58 ( .A(PCplus4[26]), .B(PCplus4_regD[26]), .S0(n40), .Y(
        PCplus4_actual[26]) );
  CLKMX2X2 U59 ( .A(PCplus4_regD[31]), .B(PCplus4[31]), .S0(n50), .Y(
        PCplus4_actual[31]) );
  NAND2X1 U60 ( .A(n11), .B(n143), .Y(PCnext[19]) );
  OA21XL U61 ( .A0(n52), .A1(n145), .B0(n144), .Y(n11) );
  NOR3X2 U62 ( .A(n36), .B(n37), .C(n38), .Y(n143) );
  OA21XL U63 ( .A0(n52), .A1(n169), .B0(n168), .Y(n28) );
  NAND2X1 U64 ( .A(n35), .B(n151), .Y(PCnext[21]) );
  NAND2X2 U65 ( .A(n189), .B(n188), .Y(PCnext[30]) );
  AOI222X1 U66 ( .A0(JumpRegAddr[8]), .A1(n56), .B0(targetAddr[6]), .B1(n51), 
        .C0(ADDresult[8]), .C1(n55), .Y(n99) );
  NAND2X2 U67 ( .A(n183), .B(n182), .Y(PCnext[28]) );
  NOR3X2 U68 ( .A(n18), .B(n19), .C(n20), .Y(n183) );
  NAND2X2 U69 ( .A(n186), .B(n185), .Y(PCnext[29]) );
  NOR3X4 U70 ( .A(n8), .B(n9), .C(n10), .Y(n139) );
  NOR3X4 U71 ( .A(n22), .B(n23), .C(n24), .Y(n171) );
  OAI211X1 U72 ( .A0(n52), .A1(n137), .B0(n136), .C0(n135), .Y(PCnext[17]) );
  OAI211X1 U73 ( .A0(n53), .A1(n121), .B0(n120), .C0(n119), .Y(PCnext[13]) );
  NAND2X2 U74 ( .A(n196), .B(n195), .Y(PCnext[31]) );
  AND3X6 U75 ( .A(n25), .B(n26), .C(n27), .Y(n196) );
  AOI222X1 U76 ( .A0(JumpRegAddr[4]), .A1(n57), .B0(targetAddr[2]), .B1(n51), 
        .C0(ADDresult[4]), .C1(n55), .Y(n83) );
  NAND2X1 U77 ( .A(n180), .B(n54), .Y(n190) );
  AOI222X1 U78 ( .A0(JumpRegAddr[9]), .A1(n56), .B0(targetAddr[7]), .B1(n51), 
        .C0(ADDresult[9]), .C1(n55), .Y(n103) );
  AOI222X1 U79 ( .A0(JumpRegAddr[21]), .A1(n191), .B0(targetAddr[19]), .B1(
        n175), .C0(ADDresult[21]), .C1(n55), .Y(n151) );
  CLKINVX3 U80 ( .A(n60), .Y(n58) );
  INVX3 U81 ( .A(n67), .Y(n194) );
  CLKINVX1 U82 ( .A(n193), .Y(n60) );
  OR2X1 U83 ( .A(n47), .B(n46), .Y(n1) );
  CLKBUFX3 U84 ( .A(n179), .Y(n54) );
  AND2XL U85 ( .A(JumpRegAddr[14]), .B(n56), .Y(n2) );
  AND2X2 U86 ( .A(targetAddr[12]), .B(n51), .Y(n5) );
  NOR3X4 U87 ( .A(n2), .B(n5), .C(n6), .Y(n123) );
  CLKBUFX6 U88 ( .A(n49), .Y(n55) );
  CLKBUFX3 U89 ( .A(n191), .Y(n56) );
  MX2X4 U90 ( .A(PCplus4_regD[11]), .B(PCplus4[11]), .S0(n64), .Y(
        PCplus4_actual[11]) );
  INVX3 U91 ( .A(n7), .Y(n73) );
  OAI211XL U92 ( .A0(n53), .A1(n101), .B0(n100), .C0(n99), .Y(PCnext[8]) );
  CLKAND2X12 U93 ( .A(ADDresult[26]), .B(n55), .Y(n24) );
  OAI211X2 U94 ( .A0(n52), .A1(n125), .B0(n124), .C0(n123), .Y(PCnext[14]) );
  MX2X2 U95 ( .A(branchOffset_regD[9]), .B(branchOffset_I[9]), .S0(n64), .Y(
        branchOffset_actual[11]) );
  CLKMX2X2 U96 ( .A(PCplus4_regD[10]), .B(PCplus4[10]), .S0(n64), .Y(
        PCplus4_actual[10]) );
  CLKBUFX2 U97 ( .A(PCsrc[2]), .Y(n7) );
  CLKMX2X3 U98 ( .A(PCplus4_regD[4]), .B(PCplus4[4]), .S0(n64), .Y(
        PCplus4_actual[4]) );
  AOI222X2 U99 ( .A0(JumpRegAddr[17]), .A1(n56), .B0(targetAddr[15]), .B1(n175), .C0(ADDresult[17]), .C1(n55), .Y(n135) );
  CLKMX2X8 U100 ( .A(branchOffset_regD[1]), .B(branchOffset_I[1]), .S0(n64), 
        .Y(branchOffset_actual[3]) );
  INVX8 U101 ( .A(PCsrc[1]), .Y(n74) );
  BUFX16 U102 ( .A(n64), .Y(n50) );
  OAI211X2 U103 ( .A0(n52), .A1(n129), .B0(n128), .C0(n127), .Y(PCnext[15]) );
  CLKMX2X2 U104 ( .A(PCplus4_regD[3]), .B(PCplus4[3]), .S0(n64), .Y(
        PCplus4_actual[3]) );
  AOI222X2 U105 ( .A0(JumpRegAddr[12]), .A1(n56), .B0(targetAddr[10]), .B1(n51), .C0(ADDresult[12]), .C1(n55), .Y(n115) );
  AOI222X2 U106 ( .A0(JumpRegAddr[13]), .A1(n56), .B0(targetAddr[11]), .B1(n51), .C0(ADDresult[13]), .C1(n55), .Y(n119) );
  AND2X8 U107 ( .A(ADDresult[27]), .B(n55), .Y(n31) );
  AND2X2 U108 ( .A(JumpRegAddr[27]), .B(n191), .Y(n29) );
  CLKAND2X2 U109 ( .A(JumpRegAddr[18]), .B(n56), .Y(n8) );
  AND2X1 U110 ( .A(targetAddr[16]), .B(n51), .Y(n9) );
  CLKAND2X12 U111 ( .A(ADDresult[18]), .B(n55), .Y(n10) );
  OAI211X2 U112 ( .A0(n52), .A1(n141), .B0(n140), .C0(n139), .Y(PCnext[18]) );
  AND2X1 U113 ( .A(JumpRegAddr[23]), .B(n191), .Y(n12) );
  AND2X1 U114 ( .A(targetAddr[21]), .B(n51), .Y(n13) );
  AND2X1 U115 ( .A(JumpRegAddr[24]), .B(n57), .Y(n15) );
  AND2X1 U116 ( .A(targetAddr[22]), .B(n51), .Y(n16) );
  NOR3X4 U117 ( .A(n15), .B(n16), .C(n17), .Y(n163) );
  OAI211X2 U118 ( .A0(n52), .A1(n165), .B0(n164), .C0(n163), .Y(PCnext[24]) );
  AND2X1 U119 ( .A(JumpRegAddr[28]), .B(n191), .Y(n18) );
  AND2X1 U120 ( .A(PCplus4[28]), .B(n190), .Y(n19) );
  NOR2X4 U121 ( .A(n48), .B(n1), .Y(n189) );
  CLKAND2X3 U122 ( .A(ADDresult[30]), .B(n55), .Y(n48) );
  AND2X1 U123 ( .A(JumpRegAddr[26]), .B(n56), .Y(n22) );
  AND2X2 U124 ( .A(targetAddr[24]), .B(n51), .Y(n23) );
  NAND2XL U125 ( .A(PCplus4[31]), .B(n190), .Y(n26) );
  NAND2X6 U126 ( .A(ADDresult[31]), .B(n55), .Y(n27) );
  BUFX4 U127 ( .A(n54), .Y(n52) );
  AND2X2 U128 ( .A(targetAddr[25]), .B(n51), .Y(n30) );
  AND2XL U129 ( .A(JumpRegAddr[25]), .B(n56), .Y(n32) );
  AND2XL U130 ( .A(targetAddr[23]), .B(n51), .Y(n33) );
  OA21XL U131 ( .A0(n52), .A1(n153), .B0(n152), .Y(n35) );
  AND2X1 U132 ( .A(JumpRegAddr[19]), .B(n56), .Y(n36) );
  CLKAND2X2 U133 ( .A(targetAddr[17]), .B(n175), .Y(n37) );
  CLKAND2X12 U134 ( .A(ADDresult[19]), .B(n55), .Y(n38) );
  CLKINVX1 U135 ( .A(n50), .Y(n40) );
  CLKINVX1 U136 ( .A(n50), .Y(n41) );
  NAND2X8 U137 ( .A(n49), .B(n65), .Y(n63) );
  AOI222X1 U138 ( .A0(JumpRegAddr[5]), .A1(n57), .B0(targetAddr[3]), .B1(n51), 
        .C0(ADDresult[5]), .C1(n55), .Y(n87) );
  AOI222X1 U139 ( .A0(JumpRegAddr[7]), .A1(n57), .B0(targetAddr[5]), .B1(n51), 
        .C0(ADDresult[7]), .C1(n55), .Y(n95) );
  AOI222X2 U140 ( .A0(JumpRegAddr[16]), .A1(n56), .B0(targetAddr[14]), .B1(n51), .C0(ADDresult[16]), .C1(n55), .Y(n131) );
  AOI222X2 U141 ( .A0(JumpRegAddr[15]), .A1(n56), .B0(targetAddr[13]), .B1(n51), .C0(ADDresult[15]), .C1(n55), .Y(n127) );
  CLKINVX3 U142 ( .A(n60), .Y(n59) );
  BUFX6 U143 ( .A(PCplus4_actual[10]), .Y(n42) );
  AND2XL U144 ( .A(PCplus4[30]), .B(n190), .Y(n47) );
  AND2XL U145 ( .A(JumpRegAddr[29]), .B(n56), .Y(n43) );
  AND2XL U146 ( .A(PCplus4[29]), .B(n190), .Y(n44) );
  NOR3X2 U147 ( .A(n43), .B(n44), .C(n45), .Y(n186) );
  MX2X1 U148 ( .A(PCplus4_regD[23]), .B(PCplus4[23]), .S0(n64), .Y(
        PCplus4_actual[23]) );
  CLKBUFX2 U149 ( .A(n191), .Y(n57) );
  CLKINVX20 U150 ( .A(n63), .Y(n64) );
  INVXL U151 ( .A(PCplus4[20]), .Y(n149) );
  AOI2BB2XL U152 ( .B0(PCcur[20]), .B1(n62), .A0N(n59), .A1N(n146), .Y(n148)
         );
  INVXL U153 ( .A(PCplus4[19]), .Y(n145) );
  AOI2BB2XL U154 ( .B0(PCcur[19]), .B1(n62), .A0N(n59), .A1N(n142), .Y(n144)
         );
  CLKMX2X3 U155 ( .A(PCplus4_regD[21]), .B(PCplus4[21]), .S0(n64), .Y(
        PCplus4_actual[21]) );
  AND2XL U156 ( .A(JumpRegAddr[30]), .B(n191), .Y(n46) );
  INVXL U157 ( .A(PCplus4[27]), .Y(n178) );
  AOI2BB2XL U158 ( .B0(PCcur[27]), .B1(n194), .A0N(n58), .A1N(n174), .Y(n177)
         );
  INVXL U159 ( .A(PCplus4[25]), .Y(n169) );
  AOI2BB2XL U160 ( .B0(PCcur[25]), .B1(n62), .A0N(n59), .A1N(n166), .Y(n168)
         );
  AOI2BB2XL U161 ( .B0(PCcur[21]), .B1(n62), .A0N(n59), .A1N(n150), .Y(n152)
         );
  INVXL U162 ( .A(PCplus4[18]), .Y(n141) );
  AOI2BB2XL U163 ( .B0(PCcur[18]), .B1(n62), .A0N(n59), .A1N(n138), .Y(n140)
         );
  INVXL U164 ( .A(PCplus4[16]), .Y(n133) );
  AOI2BB2XL U165 ( .B0(PCcur[16]), .B1(n62), .A0N(n59), .A1N(n130), .Y(n132)
         );
  INVXL U166 ( .A(PCplus4[15]), .Y(n129) );
  AOI2BB2XL U167 ( .B0(PCcur[15]), .B1(n62), .A0N(n59), .A1N(n126), .Y(n128)
         );
  AOI2BB2XL U168 ( .B0(PCcur[17]), .B1(n62), .A0N(n59), .A1N(n134), .Y(n136)
         );
  AOI2BB2XL U169 ( .B0(PCcur[31]), .B1(n61), .A0N(n59), .A1N(n192), .Y(n195)
         );
  AOI2BB2XL U170 ( .B0(PCcur[30]), .B1(n62), .A0N(n58), .A1N(n187), .Y(n188)
         );
  AOI2BB2XL U171 ( .B0(PCcur[29]), .B1(n194), .A0N(n58), .A1N(n184), .Y(n185)
         );
  AOI2BB2XL U172 ( .B0(PCcur[28]), .B1(n61), .A0N(n58), .A1N(n181), .Y(n182)
         );
  AOI2BB2XL U173 ( .B0(PCcur[6]), .B1(n61), .A0N(n58), .A1N(n90), .Y(n92) );
  INVXL U174 ( .A(PCplus4[14]), .Y(n125) );
  AOI2BB2XL U175 ( .B0(PCcur[14]), .B1(n62), .A0N(n59), .A1N(n122), .Y(n124)
         );
  INVXL U176 ( .A(PCplus4[13]), .Y(n121) );
  AOI2BB2XL U177 ( .B0(PCcur[13]), .B1(n62), .A0N(n58), .A1N(n118), .Y(n120)
         );
  INVXL U178 ( .A(PCplus4[12]), .Y(n117) );
  AOI2BB2XL U179 ( .B0(PCcur[12]), .B1(n61), .A0N(n58), .A1N(n114), .Y(n116)
         );
  INVXL U180 ( .A(PCplus4[11]), .Y(n113) );
  AOI2BB2XL U181 ( .B0(PCcur[11]), .B1(n61), .A0N(n58), .A1N(n110), .Y(n112)
         );
  AOI2BB2XL U182 ( .B0(PCcur[8]), .B1(n61), .A0N(n58), .A1N(n98), .Y(n100) );
  AOI2BB2XL U183 ( .B0(PCcur[7]), .B1(n61), .A0N(n58), .A1N(n94), .Y(n96) );
  AOI2BB2XL U184 ( .B0(PCcur[9]), .B1(n61), .A0N(n58), .A1N(n102), .Y(n104) );
  INVXL U185 ( .A(PCplus4[10]), .Y(n109) );
  AOI2BB2XL U186 ( .B0(PCcur[10]), .B1(n61), .A0N(n58), .A1N(n106), .Y(n108)
         );
  AOI222X1 U187 ( .A0(JumpRegAddr[10]), .A1(n56), .B0(targetAddr[8]), .B1(n51), 
        .C0(ADDresult[10]), .C1(n55), .Y(n107) );
  AOI2BB2XL U188 ( .B0(PCcur[3]), .B1(n61), .A0N(n58), .A1N(n78), .Y(n80) );
  OAI211XL U189 ( .A0(n53), .A1(n81), .B0(n80), .C0(n79), .Y(PCnext[3]) );
  CLKMX2X4 U190 ( .A(PCplus4_regD[28]), .B(PCplus4[28]), .S0(n50), .Y(
        PCplus4_actual[28]) );
  AOI2BB2XL U191 ( .B0(PCcur[2]), .B1(n61), .A0N(n58), .A1N(n72), .Y(n76) );
  MX2XL U192 ( .A(PCplus4_regD[1]), .B(PCplus4[1]), .S0(n50), .Y(
        PCplus4_actual[1]) );
  MX2XL U193 ( .A(PCplus4_regD[0]), .B(PCplus4[0]), .S0(n50), .Y(
        PCplus4_actual[0]) );
  CLKBUFX3 U194 ( .A(n179), .Y(n53) );
  CLKBUFX3 U195 ( .A(n194), .Y(n61) );
  CLKINVX1 U196 ( .A(PCplus4[5]), .Y(n89) );
  CLKINVX1 U197 ( .A(PCplus4[17]), .Y(n137) );
  OAI211X1 U198 ( .A0(n53), .A1(n113), .B0(n112), .C0(n111), .Y(PCnext[11]) );
  OAI211X1 U199 ( .A0(n53), .A1(n109), .B0(n108), .C0(n107), .Y(PCnext[10]) );
  CLKINVX1 U200 ( .A(PCplus4[26]), .Y(n173) );
  AOI2BB2X1 U201 ( .B0(PCcur[26]), .B1(n194), .A0N(n58), .A1N(n170), .Y(n172)
         );
  CLKINVX1 U202 ( .A(PCplus4[24]), .Y(n165) );
  AOI2BB2X1 U203 ( .B0(PCcur[24]), .B1(n62), .A0N(n59), .A1N(n162), .Y(n164)
         );
  CLKINVX1 U204 ( .A(PCplus4[23]), .Y(n161) );
  AOI2BB2X1 U205 ( .B0(PCcur[23]), .B1(n62), .A0N(n59), .A1N(n158), .Y(n160)
         );
  CLKINVX1 U206 ( .A(PCplus4[22]), .Y(n157) );
  AOI2BB2X1 U207 ( .B0(PCcur[22]), .B1(n62), .A0N(n59), .A1N(n154), .Y(n156)
         );
  CLKINVX1 U208 ( .A(PCplus4[21]), .Y(n153) );
  OAI211X1 U209 ( .A0(n53), .A1(n105), .B0(n104), .C0(n103), .Y(PCnext[9]) );
  CLKINVX1 U210 ( .A(PCplus4[9]), .Y(n105) );
  CLKINVX1 U211 ( .A(PCplus4[8]), .Y(n101) );
  CLKINVX1 U212 ( .A(PCplus4[7]), .Y(n97) );
  OAI211X1 U213 ( .A0(n53), .A1(n93), .B0(n92), .C0(n91), .Y(PCnext[6]) );
  CLKINVX1 U214 ( .A(PCplus4[6]), .Y(n93) );
  OAI211X1 U215 ( .A0(n53), .A1(n85), .B0(n84), .C0(n83), .Y(PCnext[4]) );
  CLKINVX1 U216 ( .A(PCplus4[4]), .Y(n85) );
  CLKINVX1 U217 ( .A(PCplus4[3]), .Y(n81) );
  OAI211X1 U218 ( .A0(n53), .A1(n77), .B0(n76), .C0(n75), .Y(PCnext[2]) );
  CLKINVX1 U219 ( .A(PCplus4[2]), .Y(n77) );
  CLKMX2X2 U220 ( .A(PCplus4_regD[19]), .B(PCplus4[19]), .S0(n64), .Y(
        PCplus4_actual[19]) );
  NAND2X1 U221 ( .A(n71), .B(n70), .Y(PCnext[1]) );
  AOI2BB2X1 U222 ( .B0(PCcur[1]), .B1(n61), .A0N(n197), .A1N(n54), .Y(n70) );
  AOI222XL U223 ( .A0(PCplus4_regD[1]), .A1(n60), .B0(ADDresult[1]), .B1(n55), 
        .C0(JumpRegAddr[1]), .C1(n57), .Y(n71) );
  CLKINVX1 U224 ( .A(PCplus4[1]), .Y(n197) );
  NAND2X1 U225 ( .A(n69), .B(n68), .Y(PCnext[0]) );
  AOI2BB2X1 U226 ( .B0(PCcur[0]), .B1(n61), .A0N(n198), .A1N(n54), .Y(n68) );
  AOI222XL U227 ( .A0(PCplus4_regD[0]), .A1(n60), .B0(ADDresult[0]), .B1(n55), 
        .C0(JumpRegAddr[0]), .C1(n57), .Y(n69) );
  CLKINVX1 U228 ( .A(PCplus4[0]), .Y(n198) );
  CLKINVX1 U229 ( .A(PCplus4_regD[29]), .Y(n184) );
  CLKINVX1 U230 ( .A(PCplus4_regD[31]), .Y(n192) );
  CLKINVX1 U231 ( .A(PCplus4_regD[30]), .Y(n187) );
  CLKINVX1 U232 ( .A(PCplus4_regD[28]), .Y(n181) );
  CLKINVX1 U233 ( .A(PCplus4_regD[10]), .Y(n106) );
  CLKINVX1 U234 ( .A(PCplus4_regD[3]), .Y(n78) );
  CLKINVX1 U235 ( .A(PCplus4_regD[13]), .Y(n118) );
  CLKINVX1 U236 ( .A(PCplus4_regD[11]), .Y(n110) );
  CLKINVX1 U237 ( .A(PCplus4_regD[27]), .Y(n174) );
  CLKINVX1 U238 ( .A(PCplus4_regD[26]), .Y(n170) );
  CLKINVX1 U239 ( .A(PCplus4_regD[25]), .Y(n166) );
  CLKINVX1 U240 ( .A(PCplus4_regD[24]), .Y(n162) );
  CLKINVX1 U241 ( .A(PCplus4_regD[23]), .Y(n158) );
  CLKINVX1 U242 ( .A(PCplus4_regD[22]), .Y(n154) );
  CLKINVX1 U243 ( .A(PCplus4_regD[21]), .Y(n150) );
  CLKINVX1 U244 ( .A(PCplus4_regD[20]), .Y(n146) );
  CLKINVX1 U245 ( .A(PCplus4_regD[19]), .Y(n142) );
  CLKINVX1 U246 ( .A(PCplus4_regD[18]), .Y(n138) );
  CLKINVX1 U247 ( .A(PCplus4_regD[17]), .Y(n134) );
  CLKINVX1 U248 ( .A(PCplus4_regD[16]), .Y(n130) );
  CLKINVX1 U249 ( .A(PCplus4_regD[15]), .Y(n126) );
  CLKINVX1 U250 ( .A(PCplus4_regD[14]), .Y(n122) );
  CLKINVX1 U251 ( .A(PCplus4_regD[12]), .Y(n114) );
  CLKINVX1 U252 ( .A(PCplus4_regD[9]), .Y(n102) );
  CLKINVX1 U253 ( .A(PCplus4_regD[8]), .Y(n98) );
  CLKINVX1 U254 ( .A(PCplus4_regD[7]), .Y(n94) );
  CLKINVX1 U255 ( .A(PCplus4_regD[6]), .Y(n90) );
  CLKINVX1 U256 ( .A(PCplus4_regD[2]), .Y(n72) );
  CLKINVX1 U257 ( .A(PCplus4_regD[4]), .Y(n82) );
  CLKINVX1 U258 ( .A(PCplus4_regD[5]), .Y(n86) );
  AOI2BB2XL U259 ( .B0(PCcur[5]), .B1(n61), .A0N(n58), .A1N(n86), .Y(n88) );
  OAI211X1 U260 ( .A0(n53), .A1(n89), .B0(n88), .C0(n87), .Y(PCnext[5]) );
  AOI222XL U261 ( .A0(JumpRegAddr[2]), .A1(n57), .B0(targetAddr[0]), .B1(n51), 
        .C0(ADDresult[2]), .C1(n55), .Y(n75) );
  AOI2BB2XL U262 ( .B0(PCcur[4]), .B1(n61), .A0N(n58), .A1N(n82), .Y(n84) );
  AOI222XL U263 ( .A0(JumpRegAddr[3]), .A1(n57), .B0(targetAddr[1]), .B1(n51), 
        .C0(ADDresult[3]), .C1(n55), .Y(n79) );
  NAND3BXL U264 ( .AN(PCsrc[1]), .B(PCsrc[0]), .C(n73), .Y(n67) );
  NAND3BXL U265 ( .AN(PCsrc[0]), .B(PCsrc[1]), .C(n73), .Y(n193) );
  NAND3BXL U266 ( .AN(n74), .B(n7), .C(n65), .Y(n66) );
  NAND3BXL U267 ( .AN(PCsrc[0]), .B(n74), .C(n73), .Y(n179) );
  NAND3BXL U268 ( .AN(n74), .B(PCsrc[0]), .C(n73), .Y(n180) );
  CLKINVX3 U269 ( .A(PCsrc[0]), .Y(n65) );
  CLKMX2X4 U270 ( .A(PCplus4_regD[24]), .B(PCplus4[24]), .S0(n50), .Y(
        PCplus4_actual[24]) );
  CLKMX2X4 U271 ( .A(PCplus4_regD[22]), .B(PCplus4[22]), .S0(n64), .Y(
        PCplus4_actual[22]) );
  CLKMX2X4 U272 ( .A(PCplus4_regD[20]), .B(PCplus4[20]), .S0(n64), .Y(
        PCplus4_actual[20]) );
  CLKMX2X4 U273 ( .A(PCplus4_regD[14]), .B(PCplus4[14]), .S0(n64), .Y(
        PCplus4_actual[14]) );
  CLKMX2X4 U274 ( .A(PCplus4_regD[6]), .B(PCplus4[6]), .S0(n64), .Y(
        PCplus4_actual[6]) );
  CLKMX2X4 U275 ( .A(PCplus4_regD[2]), .B(PCplus4[2]), .S0(n64), .Y(
        PCplus4_actual[2]) );
  CLKMX2X4 U276 ( .A(branchOffset_regD[8]), .B(branchOffset_I[8]), .S0(n64), 
        .Y(branchOffset_actual[10]) );
  CLKMX2X4 U277 ( .A(branchOffset_regD[4]), .B(branchOffset_I[4]), .S0(n64), 
        .Y(branchOffset_actual[6]) );
  CLKMX2X4 U278 ( .A(branchOffset_regD[2]), .B(branchOffset_I[2]), .S0(n64), 
        .Y(branchOffset_actual[4]) );
  CLKMX2X4 U279 ( .A(branchOffset_regD[0]), .B(branchOffset_I[0]), .S0(n64), 
        .Y(branchOffset_actual[2]) );
endmodule


module PCsrcLogic ( pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, 
        predict, stallcache, stall_lw_use, PCsrc );
  output [2:0] PCsrc;
  input pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, predict,
         stallcache, stall_lw_use;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  INVX1 U3 ( .A(n3), .Y(n2) );
  CLKINVX12 U4 ( .A(stallcache), .Y(n3) );
  CLKMX2X4 U5 ( .A(Jump), .B(n7), .S0(n1), .Y(n6) );
  MX2X2 U6 ( .A(Jump), .B(equal), .S0(n1), .Y(n4) );
  AOI211X2 U7 ( .A0(n10), .A1(n9), .B0(n2), .C0(stall_lw_use), .Y(PCsrc[2]) );
  CLKMX2X6 U8 ( .A(n8), .B(n7), .S0(n1), .Y(n10) );
  AOI2BB1X4 U9 ( .A0N(JumpReg), .A1N(n6), .B0(n5), .Y(PCsrc[1]) );
  NAND2BX4 U10 ( .AN(stall_lw_use), .B(n3), .Y(n5) );
  AND2X8 U11 ( .A(Branch_EX), .B(pred_cond), .Y(n1) );
  INVXL U12 ( .A(JumpReg), .Y(n9) );
  CLKINVX1 U13 ( .A(equal), .Y(n7) );
  NAND3BX4 U14 ( .AN(Jump), .B(Branch_IF), .C(predict), .Y(n8) );
  AO21X4 U15 ( .A0(n4), .A1(n9), .B0(n5), .Y(PCsrc[0]) );
endmodule


module ALU_DW_leftsh_0 ( A, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  wire   n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497;

  NOR4X1 U255 ( .A(n353), .B(n351), .C(n385), .D(n327), .Y(B[14]) );
  MXI2X1 U256 ( .A(n414), .B(n415), .S0(n345), .Y(n368) );
  NOR4X1 U257 ( .A(n354), .B(n351), .C(n329), .D(n374), .Y(B[3]) );
  INVX4 U258 ( .A(n338), .Y(n336) );
  BUFX6 U259 ( .A(n344), .Y(n343) );
  CLKINVX8 U260 ( .A(n334), .Y(n331) );
  MX2XL U261 ( .A(A[24]), .B(A[25]), .S0(n330), .Y(n405) );
  MXI2X1 U262 ( .A(n448), .B(n449), .S0(n345), .Y(n402) );
  CLKMX2X2 U263 ( .A(A[17]), .B(A[18]), .S0(n330), .Y(n445) );
  CLKMX2X2 U264 ( .A(A[16]), .B(A[17]), .S0(n330), .Y(n451) );
  CLKMX2X2 U265 ( .A(A[18]), .B(A[19]), .S0(n330), .Y(n440) );
  CLKMX2X2 U266 ( .A(A[22]), .B(A[23]), .S0(n330), .Y(n418) );
  MXI2X1 U267 ( .A(n451), .B(n461), .S0(n336), .Y(n439) );
  MXI2X1 U268 ( .A(n321), .B(n458), .S0(n341), .Y(n437) );
  CLKMX2X2 U269 ( .A(A[23]), .B(A[24]), .S0(n330), .Y(n411) );
  CLKMX2X2 U270 ( .A(A[25]), .B(A[26]), .S0(n330), .Y(n398) );
  MXI2X1 U271 ( .A(n472), .B(n473), .S0(n341), .Y(n432) );
  MXI2X1 U272 ( .A(n459), .B(n321), .S0(n342), .Y(n414) );
  NAND2X1 U273 ( .A(n427), .B(n347), .Y(n370) );
  MXI2X1 U274 ( .A(n464), .B(n465), .S0(n341), .Y(n421) );
  MXI2X1 U275 ( .A(n460), .B(n459), .S0(n341), .Y(n438) );
  CLKMX2X2 U276 ( .A(A[27]), .B(A[28]), .S0(n330), .Y(n388) );
  NOR4X1 U277 ( .A(n354), .B(n351), .C(n329), .D(n370), .Y(B[7]) );
  CLKINVX1 U278 ( .A(n402), .Y(n363) );
  CLKINVX1 U279 ( .A(SH[2]), .Y(n344) );
  INVX6 U280 ( .A(n339), .Y(n335) );
  CLKBUFX2 U281 ( .A(n340), .Y(n339) );
  BUFX4 U282 ( .A(n328), .Y(n327) );
  INVXL U283 ( .A(SH[3]), .Y(n348) );
  CLKBUFX3 U284 ( .A(n349), .Y(n351) );
  CLKBUFX3 U285 ( .A(n326), .Y(n329) );
  AND2X2 U286 ( .A(n322), .B(n323), .Y(n321) );
  NOR4X1 U287 ( .A(n497), .B(SH[16]), .C(SH[18]), .D(SH[17]), .Y(n491) );
  MX2X1 U288 ( .A(A[4]), .B(A[5]), .S0(n331), .Y(n477) );
  MX2X1 U289 ( .A(A[0]), .B(A[1]), .S0(n331), .Y(n476) );
  MX2XL U290 ( .A(A[11]), .B(A[12]), .S0(n331), .Y(n475) );
  MX2XL U291 ( .A(A[6]), .B(A[7]), .S0(n331), .Y(n480) );
  MX2XL U292 ( .A(A[3]), .B(A[4]), .S0(n331), .Y(n483) );
  NOR4X1 U293 ( .A(n353), .B(n351), .C(n402), .D(n329), .Y(B[11]) );
  CLKMX2X2 U294 ( .A(A[26]), .B(A[27]), .S0(n330), .Y(n393) );
  NAND2XL U295 ( .A(n477), .B(n339), .Y(n322) );
  NAND2X1 U296 ( .A(n478), .B(n335), .Y(n323) );
  NAND2XL U297 ( .A(n437), .B(n347), .Y(n372) );
  CLKMX2X2 U298 ( .A(n411), .B(n398), .S0(n339), .Y(n387) );
  MX2X1 U299 ( .A(n439), .B(n416), .S0(n343), .Y(n391) );
  NAND2XL U300 ( .A(n476), .B(n339), .Y(n458) );
  NAND2X1 U301 ( .A(n442), .B(n347), .Y(n373) );
  NAND2X1 U302 ( .A(n453), .B(n347), .Y(n389) );
  NOR2X1 U303 ( .A(n458), .B(n342), .Y(n415) );
  CLKINVX1 U304 ( .A(n394), .Y(n355) );
  CLKINVX1 U305 ( .A(n399), .Y(n356) );
  NOR2X1 U306 ( .A(n482), .B(n342), .Y(n422) );
  MXI2X1 U307 ( .A(n425), .B(n435), .S0(n336), .Y(n410) );
  MXI2X1 U308 ( .A(n456), .B(n467), .S0(n336), .Y(n444) );
  MXI2X1 U309 ( .A(n418), .B(n430), .S0(n336), .Y(n404) );
  NAND4X1 U310 ( .A(n489), .B(n490), .C(n491), .D(n492), .Y(n326) );
  NOR3XL U311 ( .A(SH[10]), .B(SH[12]), .C(SH[11]), .Y(n489) );
  INVXL U312 ( .A(n438), .Y(n361) );
  INVXL U313 ( .A(n433), .Y(n360) );
  INVXL U314 ( .A(n428), .Y(n359) );
  NOR4XL U315 ( .A(n353), .B(n351), .C(n392), .D(n327), .Y(B[13]) );
  NOR4XL U316 ( .A(n353), .B(n351), .C(n397), .D(n327), .Y(B[12]) );
  NAND2XL U317 ( .A(n432), .B(n347), .Y(n371) );
  MXI2XL U318 ( .A(n387), .B(n358), .S0(n342), .Y(n407) );
  INVX1 U319 ( .A(n414), .Y(n365) );
  NOR4XL U320 ( .A(n353), .B(n351), .C(n378), .D(n329), .Y(B[15]) );
  NOR4XL U321 ( .A(n353), .B(n351), .C(n409), .D(n329), .Y(B[10]) );
  NOR4XL U322 ( .A(n354), .B(n351), .C(n329), .D(n372), .Y(B[5]) );
  INVXL U323 ( .A(n443), .Y(n362) );
  INVX1 U324 ( .A(n421), .Y(n366) );
  INVXL U325 ( .A(n454), .Y(n364) );
  CLKBUFX2 U326 ( .A(n348), .Y(n347) );
  MX2XL U327 ( .A(n466), .B(n444), .S0(n343), .Y(n424) );
  MX2XL U328 ( .A(n460), .B(n439), .S0(n343), .Y(n417) );
  MX2XL U329 ( .A(n455), .B(n434), .S0(n343), .Y(n408) );
  MX2XL U330 ( .A(n429), .B(n404), .S0(n343), .Y(n377) );
  CLKBUFX2 U331 ( .A(n340), .Y(n338) );
  MXI3X1 U332 ( .A(n381), .B(n393), .C(n355), .S0(n337), .S1(n342), .Y(n324)
         );
  MXI3X1 U333 ( .A(n388), .B(n398), .C(n356), .S0(n337), .S1(n342), .Y(n325)
         );
  MXI2XL U334 ( .A(n430), .B(n440), .S0(n336), .Y(n416) );
  NAND2XL U335 ( .A(n488), .B(n339), .Y(n482) );
  MX2XL U336 ( .A(n405), .B(n393), .S0(n339), .Y(n380) );
  CLKBUFX2 U337 ( .A(SH[0]), .Y(n334) );
  NOR4XL U338 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n496) );
  NOR3XL U339 ( .A(SH[26]), .B(SH[28]), .C(SH[27]), .Y(n494) );
  NOR3XL U340 ( .A(SH[23]), .B(SH[25]), .C(SH[24]), .Y(n493) );
  OR4XL U341 ( .A(SH[20]), .B(SH[19]), .C(SH[22]), .D(SH[21]), .Y(n497) );
  CLKBUFX2 U342 ( .A(SH[0]), .Y(n333) );
  INVX3 U343 ( .A(n343), .Y(n341) );
  INVX3 U344 ( .A(n343), .Y(n342) );
  INVX3 U345 ( .A(n348), .Y(n345) );
  INVX3 U346 ( .A(n347), .Y(n346) );
  CLKINVX1 U347 ( .A(n338), .Y(n337) );
  CLKINVX1 U348 ( .A(n410), .Y(n358) );
  CLKINVX1 U349 ( .A(n374), .Y(n367) );
  CLKINVX1 U350 ( .A(n404), .Y(n357) );
  CLKBUFX3 U351 ( .A(n349), .Y(n350) );
  CLKBUFX3 U352 ( .A(n352), .Y(n354) );
  CLKBUFX3 U353 ( .A(n352), .Y(n353) );
  INVX3 U354 ( .A(SH[0]), .Y(n330) );
  CLKBUFX3 U355 ( .A(n326), .Y(n328) );
  CLKINVX1 U356 ( .A(SH[1]), .Y(n340) );
  CLKINVX1 U357 ( .A(n333), .Y(n332) );
  CLKBUFX3 U358 ( .A(SH[4]), .Y(n349) );
  CLKBUFX3 U359 ( .A(SH[5]), .Y(n352) );
  MX2XL U360 ( .A(A[12]), .B(A[13]), .S0(n331), .Y(n471) );
  MX2XL U361 ( .A(A[10]), .B(A[11]), .S0(n331), .Y(n481) );
  MX2XL U362 ( .A(A[8]), .B(A[9]), .S0(n331), .Y(n479) );
  MX2XL U363 ( .A(A[7]), .B(A[8]), .S0(n332), .Y(n485) );
  MX2XL U364 ( .A(A[9]), .B(A[10]), .S0(n332), .Y(n487) );
  MX2X1 U365 ( .A(A[28]), .B(A[29]), .S0(n330), .Y(n381) );
  MX2XL U366 ( .A(A[15]), .B(A[16]), .S0(n331), .Y(n456) );
  MX2XL U367 ( .A(A[19]), .B(A[20]), .S0(n330), .Y(n435) );
  MX2XL U368 ( .A(A[20]), .B(A[21]), .S0(n330), .Y(n430) );
  MX2XL U369 ( .A(A[13]), .B(A[14]), .S0(n331), .Y(n467) );
  MX2XL U370 ( .A(A[21]), .B(A[22]), .S0(n330), .Y(n425) );
  MX2XL U371 ( .A(A[14]), .B(A[15]), .S0(n331), .Y(n461) );
  MX2X1 U372 ( .A(A[1]), .B(A[2]), .S0(n331), .Y(n484) );
  MX2XL U373 ( .A(A[2]), .B(A[3]), .S0(n331), .Y(n478) );
  NOR4X1 U374 ( .A(n353), .B(n351), .C(n368), .D(n329), .Y(B[9]) );
  NOR4X1 U375 ( .A(n353), .B(n351), .C(n369), .D(n329), .Y(B[8]) );
  NOR4X1 U376 ( .A(n354), .B(n351), .C(n329), .D(n371), .Y(B[6]) );
  NOR4X1 U377 ( .A(n353), .B(n351), .C(n329), .D(n373), .Y(B[4]) );
  NOR3X1 U378 ( .A(n375), .B(SH[5]), .C(n327), .Y(B[31]) );
  MX3XL U379 ( .A(n376), .B(n377), .C(n378), .S0(n346), .S1(n350), .Y(n375) );
  MXI2X1 U380 ( .A(n379), .B(n380), .S0(n341), .Y(n376) );
  MX3XL U381 ( .A(A[31]), .B(A[30]), .C(n381), .S0(n333), .S1(n336), .Y(n379)
         );
  NOR3X1 U382 ( .A(n382), .B(n354), .C(n327), .Y(B[30]) );
  MX3XL U383 ( .A(n383), .B(n384), .C(n385), .S0(n345), .S1(n350), .Y(n382) );
  MXI2X1 U384 ( .A(n386), .B(n387), .S0(n341), .Y(n383) );
  MX3XL U385 ( .A(A[30]), .B(A[29]), .C(n388), .S0(n334), .S1(n336), .Y(n386)
         );
  NOR4X1 U386 ( .A(n353), .B(n351), .C(n329), .D(n389), .Y(B[2]) );
  NOR3X1 U387 ( .A(n390), .B(n354), .C(n327), .Y(B[29]) );
  MX3XL U388 ( .A(n324), .B(n391), .C(n392), .S0(n346), .S1(n350), .Y(n390) );
  NOR3X1 U389 ( .A(n395), .B(SH[5]), .C(n327), .Y(B[28]) );
  MX3XL U390 ( .A(n325), .B(n396), .C(n397), .S0(n346), .S1(n350), .Y(n395) );
  NOR3X1 U391 ( .A(n400), .B(n354), .C(n327), .Y(B[27]) );
  MXI2X1 U392 ( .A(n401), .B(n363), .S0(n350), .Y(n400) );
  MX3XL U393 ( .A(n380), .B(n357), .C(n403), .S0(n342), .S1(n345), .Y(n401) );
  NOR3X1 U394 ( .A(n406), .B(n354), .C(n327), .Y(B[26]) );
  MX3XL U395 ( .A(n407), .B(n408), .C(n409), .S0(n346), .S1(n350), .Y(n406) );
  NOR3X1 U396 ( .A(n412), .B(n354), .C(n327), .Y(B[25]) );
  CLKMX2X2 U397 ( .A(n413), .B(n368), .S0(n350), .Y(n412) );
  MX3XL U398 ( .A(n394), .B(n416), .C(n417), .S0(n342), .S1(n345), .Y(n413) );
  MXI2X1 U399 ( .A(n405), .B(n418), .S0(n336), .Y(n394) );
  NOR3X1 U400 ( .A(n419), .B(n354), .C(n327), .Y(B[24]) );
  CLKMX2X2 U401 ( .A(n420), .B(n369), .S0(n350), .Y(n419) );
  MXI2X1 U402 ( .A(n421), .B(n422), .S0(n345), .Y(n369) );
  MX3XL U403 ( .A(n399), .B(n423), .C(n424), .S0(n342), .S1(n345), .Y(n420) );
  MXI2X1 U404 ( .A(n411), .B(n425), .S0(n336), .Y(n399) );
  NOR3X1 U405 ( .A(n426), .B(n354), .C(n327), .Y(B[23]) );
  MX3XL U406 ( .A(n377), .B(n359), .C(n370), .S0(n346), .S1(n350), .Y(n426) );
  NOR3X1 U407 ( .A(n431), .B(n354), .C(n327), .Y(B[22]) );
  MX3XL U408 ( .A(n384), .B(n360), .C(n371), .S0(n346), .S1(n350), .Y(n431) );
  CLKMX2X2 U409 ( .A(n434), .B(n410), .S0(n344), .Y(n384) );
  NOR3X1 U410 ( .A(n436), .B(n354), .C(n327), .Y(B[21]) );
  MX3XL U411 ( .A(n391), .B(n361), .C(n372), .S0(n346), .S1(n350), .Y(n436) );
  NOR3X1 U412 ( .A(n441), .B(n354), .C(n327), .Y(B[20]) );
  MX3XL U413 ( .A(n396), .B(n362), .C(n373), .S0(n346), .S1(n351), .Y(n441) );
  CLKMX2X2 U414 ( .A(n444), .B(n423), .S0(n343), .Y(n396) );
  MXI2X1 U415 ( .A(n435), .B(n445), .S0(n336), .Y(n423) );
  NOR4X1 U416 ( .A(n353), .B(n351), .C(n329), .D(n446), .Y(B[1]) );
  NOR3BXL U417 ( .AN(n447), .B(n354), .C(n327), .Y(B[19]) );
  MX3XL U418 ( .A(n403), .B(n448), .C(n367), .S0(n346), .S1(n351), .Y(n447) );
  NAND2X1 U419 ( .A(n449), .B(n347), .Y(n374) );
  MXI2X1 U420 ( .A(n429), .B(n450), .S0(n342), .Y(n403) );
  MXI2X1 U421 ( .A(n440), .B(n451), .S0(n336), .Y(n429) );
  NOR3X1 U422 ( .A(n452), .B(n354), .C(n327), .Y(B[18]) );
  MX3XL U423 ( .A(n408), .B(n364), .C(n389), .S0(n346), .S1(n350), .Y(n452) );
  MXI2X1 U424 ( .A(n445), .B(n456), .S0(n336), .Y(n434) );
  NOR3X1 U425 ( .A(n457), .B(n354), .C(n327), .Y(B[17]) );
  MX3XL U426 ( .A(n417), .B(n365), .C(n446), .S0(n346), .S1(n351), .Y(n457) );
  NAND2X1 U427 ( .A(n415), .B(n347), .Y(n446) );
  NOR3X1 U428 ( .A(n462), .B(SH[5]), .C(n328), .Y(B[16]) );
  MX3XL U429 ( .A(n424), .B(n366), .C(n463), .S0(n345), .S1(n350), .Y(n462) );
  MXI2X1 U430 ( .A(n428), .B(n427), .S0(n345), .Y(n378) );
  MXI2X1 U431 ( .A(n468), .B(n469), .S0(n341), .Y(n427) );
  MXI2X1 U432 ( .A(n450), .B(n470), .S0(n341), .Y(n428) );
  MXI2X1 U433 ( .A(n461), .B(n471), .S0(n335), .Y(n450) );
  MXI2X1 U434 ( .A(n433), .B(n432), .S0(n345), .Y(n385) );
  MXI2X1 U435 ( .A(n455), .B(n474), .S0(n341), .Y(n433) );
  MXI2X1 U436 ( .A(n467), .B(n475), .S0(n335), .Y(n455) );
  MXI2X1 U437 ( .A(n438), .B(n437), .S0(n345), .Y(n392) );
  MXI2X1 U438 ( .A(n479), .B(n480), .S0(n335), .Y(n459) );
  MXI2X1 U439 ( .A(n471), .B(n481), .S0(n335), .Y(n460) );
  MXI2X1 U440 ( .A(n443), .B(n442), .S0(n345), .Y(n397) );
  MXI2X1 U441 ( .A(n465), .B(n482), .S0(n341), .Y(n442) );
  MXI2X1 U442 ( .A(n483), .B(n484), .S0(n335), .Y(n465) );
  MXI2X1 U443 ( .A(n466), .B(n464), .S0(n341), .Y(n443) );
  MXI2X1 U444 ( .A(n485), .B(n486), .S0(n335), .Y(n464) );
  MXI2X1 U445 ( .A(n475), .B(n487), .S0(n335), .Y(n466) );
  NOR2X1 U446 ( .A(n469), .B(n342), .Y(n449) );
  MXI2X1 U447 ( .A(n478), .B(n476), .S0(n335), .Y(n469) );
  MXI2X1 U448 ( .A(n470), .B(n468), .S0(n341), .Y(n448) );
  MXI2X1 U449 ( .A(n480), .B(n477), .S0(n335), .Y(n468) );
  MXI2X1 U450 ( .A(n481), .B(n479), .S0(n335), .Y(n470) );
  MXI2X1 U451 ( .A(n454), .B(n453), .S0(n345), .Y(n409) );
  NOR2X1 U452 ( .A(n473), .B(n342), .Y(n453) );
  MXI2X1 U453 ( .A(n484), .B(n488), .S0(n335), .Y(n473) );
  MXI2X1 U454 ( .A(n474), .B(n472), .S0(n341), .Y(n454) );
  MXI2X1 U455 ( .A(n486), .B(n483), .S0(n335), .Y(n472) );
  CLKMX2X2 U456 ( .A(A[5]), .B(A[6]), .S0(n332), .Y(n486) );
  MXI2X1 U457 ( .A(n487), .B(n485), .S0(n336), .Y(n474) );
  NOR4X1 U458 ( .A(n353), .B(n351), .C(n329), .D(n463), .Y(B[0]) );
  NAND2X1 U459 ( .A(n422), .B(n347), .Y(n463) );
  NOR2BX1 U460 ( .AN(A[0]), .B(SH[0]), .Y(n488) );
  AND4X1 U461 ( .A(n493), .B(n494), .C(n495), .D(n496), .Y(n492) );
  NOR3X1 U462 ( .A(SH[29]), .B(SH[31]), .C(SH[30]), .Y(n495) );
  NOR3X1 U463 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n490) );
endmodule


module ALU_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;

  OAI21X1 U655 ( .A0(n1333), .A1(n1334), .B0(n1335), .Y(n1318) );
  OAI31X2 U656 ( .A0(n1314), .A1(n1315), .A2(n1316), .B0(n1317), .Y(
        GE_LT_GT_LE) );
  OAI2BB1X2 U657 ( .A0N(n1332), .A1N(n1278), .B0(n1321), .Y(n1319) );
  AOI211X4 U658 ( .A0(n1294), .A1(A[20]), .B0(n1325), .C0(n1290), .Y(n1332) );
  AND2X2 U659 ( .A(A[3]), .B(n1280), .Y(n1364) );
  OR2X1 U660 ( .A(B[11]), .B(n1304), .Y(n1374) );
  OAI32X1 U661 ( .A0(n1287), .A1(A[26]), .A2(n1345), .B0(A[27]), .B1(n1286), 
        .Y(n1341) );
  OAI32X1 U662 ( .A0(n1289), .A1(A[24]), .A2(n1344), .B0(A[25]), .B1(n1288), 
        .Y(n1342) );
  OAI211X1 U663 ( .A0(B[12]), .A1(n1303), .B0(n1370), .C0(n1368), .Y(n1350) );
  OA22X2 U664 ( .A0(n1327), .A1(n1328), .B0(n1329), .B1(n1327), .Y(n1278) );
  OAI32X1 U665 ( .A0(n1292), .A1(A[22]), .A2(n1326), .B0(A[23]), .B1(n1291), 
        .Y(n1322) );
  AOI211X1 U666 ( .A0(n1289), .A1(A[24]), .B0(n1344), .C0(n1375), .Y(n1320) );
  AOI21X1 U667 ( .A0(n1282), .A1(A[30]), .B0(n1340), .Y(n1337) );
  OAI32X1 U668 ( .A0(n1300), .A1(A[14]), .A2(n1371), .B0(A[15]), .B1(n1299), 
        .Y(n1367) );
  NAND2BXL U669 ( .AN(n1333), .B(n1343), .Y(n1375) );
  NOR2BX1 U670 ( .AN(A[25]), .B(B[25]), .Y(n1344) );
  NOR2BX2 U671 ( .AN(A[27]), .B(B[27]), .Y(n1345) );
  OAI32X4 U672 ( .A0(n1296), .A1(A[18]), .A2(n1331), .B0(A[19]), .B1(n1295), 
        .Y(n1327) );
  AOI21X1 U673 ( .A0(n1296), .A1(A[18]), .B0(n1331), .Y(n1329) );
  NOR2BX4 U674 ( .AN(A[23]), .B(B[23]), .Y(n1326) );
  AO21X1 U675 ( .A0(n1298), .A1(A[16]), .B0(n1330), .Y(n1315) );
  OAI32X1 U676 ( .A0(n1279), .A1(A[2]), .A2(n1364), .B0(A[3]), .B1(n1280), .Y(
        n1362) );
  OAI21X2 U677 ( .A0(n1350), .A1(n1365), .B0(n1366), .Y(n1346) );
  OAI22X1 U678 ( .A0(n1367), .A1(n1301), .B0(n1368), .B1(n1367), .Y(n1366) );
  INVX1 U679 ( .A(n1369), .Y(n1301) );
  INVX1 U680 ( .A(n1338), .Y(n1283) );
  INVXL U681 ( .A(A[13]), .Y(n1302) );
  INVXL U682 ( .A(B[23]), .Y(n1291) );
  INVXL U683 ( .A(B[27]), .Y(n1286) );
  INVXL U684 ( .A(B[31]), .Y(n1281) );
  OAI22X1 U685 ( .A0(n1318), .A1(n1319), .B0(n1320), .B1(n1318), .Y(n1317) );
  INVXL U686 ( .A(B[19]), .Y(n1295) );
  INVX1 U687 ( .A(n1359), .Y(n1308) );
  INVXL U688 ( .A(B[25]), .Y(n1288) );
  INVXL U689 ( .A(B[21]), .Y(n1293) );
  INVXL U690 ( .A(B[15]), .Y(n1299) );
  AOI32XL U691 ( .A0(B[12]), .A1(n1303), .A2(n1370), .B0(n1302), .B1(B[13]), 
        .Y(n1369) );
  OR2XL U692 ( .A(B[13]), .B(n1302), .Y(n1370) );
  OR2XL U693 ( .A(B[9]), .B(n1306), .Y(n1352) );
  INVX1 U694 ( .A(B[30]), .Y(n1282) );
  INVXL U695 ( .A(B[26]), .Y(n1287) );
  INVXL U696 ( .A(B[6]), .Y(n1310) );
  INVXL U697 ( .A(B[14]), .Y(n1300) );
  INVXL U698 ( .A(B[17]), .Y(n1297) );
  INVXL U699 ( .A(A[11]), .Y(n1304) );
  INVXL U700 ( .A(B[7]), .Y(n1309) );
  AOI32XL U701 ( .A0(B[10]), .A1(n1305), .A2(n1374), .B0(n1304), .B1(B[11]), 
        .Y(n1372) );
  AOI32XL U702 ( .A0(B[8]), .A1(n1307), .A2(n1352), .B0(n1306), .B1(B[9]), .Y(
        n1373) );
  INVXL U703 ( .A(B[20]), .Y(n1294) );
  INVXL U704 ( .A(B[18]), .Y(n1296) );
  INVXL U705 ( .A(B[22]), .Y(n1292) );
  INVXL U706 ( .A(B[16]), .Y(n1298) );
  INVXL U707 ( .A(A[12]), .Y(n1303) );
  INVXL U708 ( .A(A[28]), .Y(n1285) );
  INVXL U709 ( .A(A[5]), .Y(n1311) );
  INVXL U710 ( .A(A[4]), .Y(n1312) );
  INVXL U711 ( .A(A[8]), .Y(n1307) );
  INVXL U712 ( .A(A[29]), .Y(n1284) );
  INVXL U713 ( .A(B[24]), .Y(n1289) );
  CLKINVX1 U714 ( .A(B[3]), .Y(n1280) );
  CLKINVX1 U715 ( .A(B[2]), .Y(n1279) );
  CLKINVX1 U716 ( .A(A[1]), .Y(n1313) );
  CLKINVX1 U717 ( .A(n1324), .Y(n1290) );
  NOR2BX1 U718 ( .AN(A[15]), .B(B[15]), .Y(n1371) );
  INVXL U719 ( .A(A[10]), .Y(n1305) );
  INVXL U720 ( .A(A[9]), .Y(n1306) );
  OAI32XL U721 ( .A0(n1294), .A1(A[20]), .A2(n1325), .B0(A[21]), .B1(n1293), 
        .Y(n1323) );
  NOR2BXL U722 ( .AN(A[21]), .B(B[21]), .Y(n1325) );
  OAI32XL U723 ( .A0(n1282), .A1(A[30]), .A2(n1340), .B0(A[31]), .B1(n1281), 
        .Y(n1336) );
  OAI32XL U724 ( .A0(n1298), .A1(A[16]), .A2(n1330), .B0(A[17]), .B1(n1297), 
        .Y(n1328) );
  AND2XL U725 ( .A(A[17]), .B(n1297), .Y(n1330) );
  AOI21XL U726 ( .A0(n1287), .A1(A[26]), .B0(n1345), .Y(n1343) );
  AOI21XL U727 ( .A0(n1300), .A1(A[14]), .B0(n1371), .Y(n1368) );
  AOI21XL U728 ( .A0(A[2]), .A1(n1279), .B0(n1364), .Y(n1363) );
  OAI32XL U729 ( .A0(n1310), .A1(A[6]), .A2(n1360), .B0(A[7]), .B1(n1309), .Y(
        n1359) );
  NOR2BXL U730 ( .AN(A[7]), .B(B[7]), .Y(n1360) );
  AOI21XL U731 ( .A0(n1292), .A1(A[22]), .B0(n1326), .Y(n1324) );
  NOR2BXL U732 ( .AN(A[19]), .B(B[19]), .Y(n1331) );
  OAI22XL U733 ( .A0(n1322), .A1(n1323), .B0(n1324), .B1(n1322), .Y(n1321) );
  OAI22XL U734 ( .A0(n1336), .A1(n1283), .B0(n1337), .B1(n1336), .Y(n1335) );
  AOI32X1 U735 ( .A0(B[28]), .A1(n1285), .A2(n1339), .B0(n1284), .B1(B[29]), 
        .Y(n1338) );
  OAI22XL U736 ( .A0(n1341), .A1(n1342), .B0(n1343), .B1(n1341), .Y(n1334) );
  OAI22XL U737 ( .A0(n1346), .A1(n1347), .B0(n1348), .B1(n1346), .Y(n1316) );
  NOR3X1 U738 ( .A(n1349), .B(n1350), .C(n1351), .Y(n1348) );
  OAI21XL U739 ( .A0(B[8]), .A1(n1307), .B0(n1352), .Y(n1349) );
  OAI31XL U740 ( .A0(n1353), .A1(n1354), .A2(n1355), .B0(n1356), .Y(n1347) );
  AO22X1 U741 ( .A0(n1308), .A1(n1357), .B0(n1355), .B1(n1308), .Y(n1356) );
  AOI32X1 U742 ( .A0(B[4]), .A1(n1312), .A2(n1358), .B0(n1311), .B1(B[5]), .Y(
        n1357) );
  AO21X1 U743 ( .A0(n1310), .A1(A[6]), .B0(n1360), .Y(n1355) );
  AOI221XL U744 ( .A0(B[1]), .A1(n1313), .B0(n1361), .B1(B[0]), .C0(n1362), 
        .Y(n1354) );
  AOI2BB1X1 U745 ( .A0N(n1313), .A1N(B[1]), .B0(A[0]), .Y(n1361) );
  OAI221XL U746 ( .A0(B[4]), .A1(n1312), .B0(n1363), .B1(n1362), .C0(n1358), 
        .Y(n1353) );
  OR2X1 U747 ( .A(B[5]), .B(n1311), .Y(n1358) );
  AO22X1 U748 ( .A0(n1372), .A1(n1373), .B0(n1351), .B1(n1372), .Y(n1365) );
  OAI21XL U749 ( .A0(B[10]), .A1(n1305), .B0(n1374), .Y(n1351) );
  NAND3X1 U750 ( .A(n1320), .B(n1332), .C(n1329), .Y(n1314) );
  OAI211X1 U751 ( .A0(B[28]), .A1(n1285), .B0(n1339), .C0(n1337), .Y(n1333) );
  NOR2BX1 U752 ( .AN(A[31]), .B(B[31]), .Y(n1340) );
  OR2X1 U753 ( .A(B[29]), .B(n1284), .Y(n1339) );
endmodule


module ALU_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493;

  MX3X1 U256 ( .A(n352), .B(n383), .C(n411), .S0(n338), .S1(n343), .Y(n452) );
  NOR3BX1 U257 ( .AN(n463), .B(n345), .C(n326), .Y(B[12]) );
  NOR3X2 U258 ( .A(n394), .B(n345), .C(n326), .Y(B[3]) );
  BUFX4 U259 ( .A(n324), .Y(n326) );
  CLKMX2X2 U260 ( .A(A[29]), .B(A[30]), .S0(n327), .Y(n454) );
  CLKMX2X2 U261 ( .A(A[23]), .B(A[24]), .S0(n327), .Y(n459) );
  CLKMX2X2 U262 ( .A(A[25]), .B(A[26]), .S0(n328), .Y(n462) );
  CLKMX2X2 U263 ( .A(A[27]), .B(A[28]), .S0(n327), .Y(n461) );
  CLKMX2X2 U264 ( .A(A[17]), .B(A[18]), .S0(n327), .Y(n456) );
  INVX8 U265 ( .A(n329), .Y(n328) );
  CLKMX2X2 U266 ( .A(A[22]), .B(A[23]), .S0(n328), .Y(n481) );
  CLKMX2X2 U267 ( .A(A[18]), .B(A[19]), .S0(n328), .Y(n479) );
  CLKMX2X2 U268 ( .A(A[16]), .B(A[17]), .S0(n328), .Y(n474) );
  CLKMX2X2 U269 ( .A(A[26]), .B(A[27]), .S0(n328), .Y(n472) );
  CLKMX2X2 U270 ( .A(A[24]), .B(A[25]), .S0(n328), .Y(n480) );
  CLKMX2X2 U271 ( .A(A[30]), .B(A[31]), .S0(n328), .Y(n473) );
  CLKMX2X2 U272 ( .A(A[15]), .B(A[16]), .S0(n327), .Y(n457) );
  MXI2X1 U273 ( .A(n453), .B(n454), .S0(n332), .Y(n437) );
  MXI2X1 U274 ( .A(n454), .B(n461), .S0(n332), .Y(n444) );
  INVX4 U275 ( .A(n330), .Y(n327) );
  MXI2X1 U276 ( .A(n447), .B(n450), .S0(n334), .Y(n433) );
  NOR2X1 U277 ( .A(n464), .B(n336), .Y(n423) );
  MXI2X1 U278 ( .A(n441), .B(n444), .S0(n334), .Y(n431) );
  MXI2X1 U279 ( .A(n473), .B(n471), .S0(n332), .Y(n464) );
  MXI2X1 U280 ( .A(n435), .B(n436), .S0(n335), .Y(n365) );
  MXI2X1 U281 ( .A(n467), .B(n468), .S0(n334), .Y(n424) );
  MXI2X1 U282 ( .A(n423), .B(n424), .S0(n338), .Y(n390) );
  CLKBUFX3 U283 ( .A(n333), .Y(n337) );
  CLKBUFX3 U284 ( .A(n342), .Y(n343) );
  MXI2X1 U285 ( .A(n430), .B(n399), .S0(n332), .Y(n387) );
  INVX4 U286 ( .A(n341), .Y(n338) );
  CLKINVX6 U287 ( .A(SH[1]), .Y(n332) );
  CLKBUFX2 U288 ( .A(SH[5]), .Y(n345) );
  CLKBUFX2 U289 ( .A(SH[3]), .Y(n341) );
  MXI3X1 U290 ( .A(n397), .B(n398), .C(n359), .S0(n332), .S1(n336), .Y(n323)
         );
  MXI2X1 U291 ( .A(n464), .B(n467), .S0(n334), .Y(n416) );
  MX2X1 U292 ( .A(A[19]), .B(A[20]), .S0(n327), .Y(n455) );
  NAND2X1 U293 ( .A(n473), .B(n332), .Y(n447) );
  INVX1 U294 ( .A(SH[0]), .Y(n331) );
  MXI2XL U295 ( .A(n476), .B(n477), .S0(n332), .Y(n379) );
  CLKBUFX4 U296 ( .A(n342), .Y(n344) );
  NAND2X1 U297 ( .A(n421), .B(n338), .Y(n411) );
  MXI2X1 U298 ( .A(n456), .B(n457), .S0(n332), .Y(n442) );
  MXI2X1 U299 ( .A(n474), .B(n475), .S0(n332), .Y(n448) );
  INVX1 U300 ( .A(n365), .Y(n355) );
  NAND2X1 U301 ( .A(n453), .B(n332), .Y(n441) );
  NAND4X1 U302 ( .A(n483), .B(n484), .C(n485), .D(n486), .Y(n324) );
  NOR3XL U303 ( .A(SH[10]), .B(SH[12]), .C(SH[11]), .Y(n483) );
  NAND2XL U304 ( .A(n433), .B(n339), .Y(n414) );
  CLKINVX3 U305 ( .A(n336), .Y(n335) );
  MX2XL U306 ( .A(n442), .B(n443), .S0(n336), .Y(n375) );
  MX2XL U307 ( .A(n448), .B(n449), .S0(n336), .Y(n381) );
  MX2XL U308 ( .A(n379), .B(n448), .S0(n336), .Y(n404) );
  MX2XL U309 ( .A(n393), .B(n466), .S0(n336), .Y(n367) );
  MX2XL U310 ( .A(n429), .B(n436), .S0(n336), .Y(n383) );
  INVXL U311 ( .A(n432), .Y(n353) );
  INVXL U312 ( .A(n422), .Y(n352) );
  INVXL U313 ( .A(n434), .Y(n354) );
  INVX1 U314 ( .A(n369), .Y(n356) );
  INVX1 U315 ( .A(n420), .Y(n351) );
  INVX1 U316 ( .A(n418), .Y(n350) );
  MXI2XL U317 ( .A(n410), .B(n407), .S0(n332), .Y(n391) );
  INVX1 U318 ( .A(n410), .Y(n360) );
  MX2XL U319 ( .A(n397), .B(n400), .S0(SH[1]), .Y(n386) );
  NOR4XL U320 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n490) );
  NOR3XL U321 ( .A(SH[26]), .B(SH[28]), .C(SH[27]), .Y(n488) );
  NOR3XL U322 ( .A(SH[23]), .B(SH[25]), .C(SH[24]), .Y(n487) );
  NOR4XL U323 ( .A(n491), .B(SH[16]), .C(SH[18]), .D(SH[17]), .Y(n485) );
  OR4XL U324 ( .A(SH[20]), .B(SH[19]), .C(SH[22]), .D(SH[21]), .Y(n491) );
  INVX1 U325 ( .A(n408), .Y(n361) );
  CLKINVX1 U326 ( .A(n390), .Y(n349) );
  INVX3 U327 ( .A(n337), .Y(n334) );
  CLKINVX1 U328 ( .A(n387), .Y(n357) );
  CLKINVX1 U329 ( .A(n393), .Y(n358) );
  CLKBUFX3 U330 ( .A(n333), .Y(n336) );
  CLKBUFX3 U331 ( .A(SH[5]), .Y(n347) );
  CLKBUFX3 U332 ( .A(SH[5]), .Y(n346) );
  CLKINVX1 U333 ( .A(n341), .Y(n339) );
  CLKINVX1 U334 ( .A(n374), .Y(n359) );
  CLKBUFX3 U335 ( .A(n331), .Y(n329) );
  CLKINVX1 U336 ( .A(n412), .Y(n348) );
  CLKBUFX3 U337 ( .A(n324), .Y(n325) );
  CLKBUFX3 U338 ( .A(n331), .Y(n330) );
  CLKBUFX3 U339 ( .A(SH[2]), .Y(n333) );
  CLKBUFX3 U340 ( .A(SH[3]), .Y(n340) );
  CLKBUFX3 U341 ( .A(SH[4]), .Y(n342) );
  MX2XL U342 ( .A(A[20]), .B(A[21]), .S0(n328), .Y(n478) );
  MX2XL U343 ( .A(A[12]), .B(A[13]), .S0(n328), .Y(n476) );
  MX2XL U344 ( .A(A[11]), .B(A[12]), .S0(n327), .Y(n430) );
  MX2XL U345 ( .A(A[8]), .B(A[9]), .S0(n328), .Y(n409) );
  MX2XL U346 ( .A(A[7]), .B(A[8]), .S0(n327), .Y(n400) );
  MX2XL U347 ( .A(A[9]), .B(A[10]), .S0(n327), .Y(n399) );
  MX2X1 U348 ( .A(A[28]), .B(A[29]), .S0(n328), .Y(n471) );
  MX2XL U349 ( .A(A[13]), .B(A[14]), .S0(n327), .Y(n458) );
  MX2XL U350 ( .A(A[14]), .B(A[15]), .S0(n328), .Y(n475) );
  MX2XL U351 ( .A(A[10]), .B(A[11]), .S0(n328), .Y(n477) );
  MXI2XL U352 ( .A(A[7]), .B(A[6]), .S0(n330), .Y(n410) );
  MX2X1 U353 ( .A(A[21]), .B(A[22]), .S0(n327), .Y(n460) );
  MX2X1 U354 ( .A(A[3]), .B(A[4]), .S0(n327), .Y(n398) );
  MXI2XL U355 ( .A(A[3]), .B(A[2]), .S0(n329), .Y(n408) );
  NOR3X1 U356 ( .A(n362), .B(n347), .C(n326), .Y(B[9]) );
  MX3XL U357 ( .A(n355), .B(n363), .C(n364), .S0(n338), .S1(n343), .Y(n362) );
  NOR3X1 U358 ( .A(n366), .B(n345), .C(n326), .Y(B[8]) );
  MX3XL U359 ( .A(n356), .B(n367), .C(n368), .S0(n338), .S1(n343), .Y(n366) );
  NOR3X1 U360 ( .A(n370), .B(n345), .C(n326), .Y(B[7]) );
  CLKMX2X2 U361 ( .A(n371), .B(n372), .S0(n343), .Y(n370) );
  MX3XL U362 ( .A(n373), .B(n374), .C(n375), .S0(n335), .S1(n341), .Y(n371) );
  NOR3X1 U363 ( .A(n376), .B(n345), .C(n326), .Y(B[6]) );
  CLKMX2X2 U364 ( .A(n377), .B(n378), .S0(n343), .Y(n376) );
  MX3XL U365 ( .A(n379), .B(n380), .C(n381), .S0(n335), .S1(n340), .Y(n377) );
  NOR3X1 U366 ( .A(n382), .B(n345), .C(n326), .Y(B[5]) );
  MX3XL U367 ( .A(n383), .B(n384), .C(n385), .S0(n338), .S1(n344), .Y(n382) );
  MXI2X1 U368 ( .A(n357), .B(n386), .S0(n335), .Y(n384) );
  NOR3X1 U369 ( .A(n388), .B(n345), .C(n326), .Y(B[4]) );
  MXI2X1 U370 ( .A(n389), .B(n349), .S0(n343), .Y(n388) );
  MX3XL U371 ( .A(n358), .B(n391), .C(n392), .S0(n335), .S1(n341), .Y(n389) );
  MX3XL U372 ( .A(n395), .B(n323), .C(n396), .S0(n338), .S1(n344), .Y(n394) );
  MXI2X1 U373 ( .A(n399), .B(n400), .S0(n332), .Y(n374) );
  NOR4X1 U374 ( .A(n346), .B(n344), .C(n325), .D(n401), .Y(B[31]) );
  NOR4X1 U375 ( .A(n346), .B(n344), .C(n325), .D(n402), .Y(B[30]) );
  NOR3X1 U376 ( .A(n403), .B(n347), .C(n326), .Y(B[2]) );
  MX3XL U377 ( .A(n404), .B(n405), .C(n406), .S0(n338), .S1(n344), .Y(n403) );
  MX3XL U378 ( .A(n407), .B(n408), .C(n380), .S0(n332), .S1(n336), .Y(n405) );
  MXI2X1 U379 ( .A(n409), .B(n360), .S0(n332), .Y(n380) );
  NOR4X1 U380 ( .A(n346), .B(n344), .C(n325), .D(n411), .Y(B[29]) );
  NOR4X1 U381 ( .A(n346), .B(n344), .C(n325), .D(n412), .Y(B[28]) );
  NOR4X1 U382 ( .A(n346), .B(n344), .C(n325), .D(n413), .Y(B[27]) );
  NOR4X1 U383 ( .A(n346), .B(n344), .C(n325), .D(n414), .Y(B[26]) );
  NOR4X1 U384 ( .A(n346), .B(n344), .C(n325), .D(n364), .Y(B[25]) );
  NAND2X1 U385 ( .A(n415), .B(n339), .Y(n364) );
  NOR4X1 U386 ( .A(n346), .B(n344), .C(n325), .D(n368), .Y(B[24]) );
  NAND2X1 U387 ( .A(n416), .B(n338), .Y(n368) );
  NOR4X1 U388 ( .A(n347), .B(n344), .C(n372), .D(n326), .Y(B[23]) );
  MXI2X1 U389 ( .A(n417), .B(n418), .S0(n338), .Y(n372) );
  NOR4X1 U390 ( .A(n346), .B(n344), .C(n378), .D(n326), .Y(B[22]) );
  MXI2X1 U391 ( .A(n419), .B(n420), .S0(n338), .Y(n378) );
  NOR4X1 U392 ( .A(n347), .B(n344), .C(n385), .D(n326), .Y(B[21]) );
  MXI2X1 U393 ( .A(n421), .B(n422), .S0(n338), .Y(n385) );
  NOR4X1 U394 ( .A(n347), .B(n344), .C(n390), .D(n325), .Y(B[20]) );
  NOR3X1 U395 ( .A(n425), .B(n347), .C(n326), .Y(B[1]) );
  MX3XL U396 ( .A(n363), .B(n426), .C(n427), .S0(n338), .S1(n343), .Y(n425) );
  MXI2X1 U397 ( .A(n386), .B(n428), .S0(n335), .Y(n426) );
  MX3XL U398 ( .A(A[2]), .B(A[1]), .C(n398), .S0(n330), .S1(SH[1]), .Y(n428)
         );
  CLKMX2X2 U399 ( .A(A[5]), .B(A[6]), .S0(n327), .Y(n397) );
  CLKMX2X2 U400 ( .A(n387), .B(n429), .S0(n336), .Y(n363) );
  NOR4X1 U401 ( .A(n346), .B(n344), .C(n396), .D(n325), .Y(B[19]) );
  MXI2X1 U402 ( .A(n431), .B(n432), .S0(n338), .Y(n396) );
  NOR4X1 U403 ( .A(n347), .B(n344), .C(n406), .D(n325), .Y(B[18]) );
  MXI2X1 U404 ( .A(n433), .B(n434), .S0(n338), .Y(n406) );
  NOR4X1 U405 ( .A(n346), .B(n344), .C(n427), .D(n325), .Y(B[17]) );
  MXI2X1 U406 ( .A(n415), .B(n365), .S0(n338), .Y(n427) );
  MXI2X1 U407 ( .A(n437), .B(n438), .S0(n334), .Y(n415) );
  NOR4X1 U408 ( .A(n346), .B(n344), .C(n439), .D(n325), .Y(B[16]) );
  NOR3X1 U409 ( .A(n440), .B(n347), .C(n326), .Y(B[15]) );
  MX3XL U410 ( .A(n350), .B(n375), .C(n401), .S0(n338), .S1(n343), .Y(n440) );
  NAND2X1 U411 ( .A(n417), .B(n339), .Y(n401) );
  NOR2X1 U412 ( .A(n441), .B(n336), .Y(n417) );
  MXI2X1 U413 ( .A(n444), .B(n445), .S0(n334), .Y(n418) );
  NOR3X1 U414 ( .A(n446), .B(n347), .C(n326), .Y(B[14]) );
  MX3XL U415 ( .A(n351), .B(n381), .C(n402), .S0(n338), .S1(n343), .Y(n446) );
  NAND2X1 U416 ( .A(n419), .B(n339), .Y(n402) );
  NOR2X1 U417 ( .A(n447), .B(n336), .Y(n419) );
  MXI2X1 U418 ( .A(n450), .B(n451), .S0(n334), .Y(n420) );
  NOR3X1 U419 ( .A(n452), .B(n347), .C(n326), .Y(B[13]) );
  NOR2X1 U420 ( .A(n437), .B(n336), .Y(n421) );
  MXI2X1 U421 ( .A(n455), .B(n456), .S0(n332), .Y(n436) );
  MXI2X1 U422 ( .A(n457), .B(n458), .S0(n332), .Y(n429) );
  MXI2X1 U423 ( .A(n438), .B(n435), .S0(n334), .Y(n422) );
  MXI2X1 U424 ( .A(n459), .B(n460), .S0(n332), .Y(n435) );
  MXI2X1 U425 ( .A(n461), .B(n462), .S0(n332), .Y(n438) );
  MX3XL U426 ( .A(n424), .B(n392), .C(n348), .S0(n339), .S1(n343), .Y(n463) );
  NAND2X1 U427 ( .A(n423), .B(n338), .Y(n412) );
  MXI2X1 U428 ( .A(n465), .B(n466), .S0(n334), .Y(n392) );
  NOR3X1 U429 ( .A(n469), .B(n347), .C(n326), .Y(B[11]) );
  MX3XL U430 ( .A(n353), .B(n395), .C(n413), .S0(n338), .S1(n343), .Y(n469) );
  NAND2X1 U431 ( .A(n431), .B(n339), .Y(n413) );
  AND2X1 U432 ( .A(A[31]), .B(n330), .Y(n453) );
  CLKMX2X2 U433 ( .A(n373), .B(n442), .S0(n337), .Y(n395) );
  MXI2X1 U434 ( .A(n458), .B(n430), .S0(n332), .Y(n373) );
  MXI2X1 U435 ( .A(n445), .B(n443), .S0(n334), .Y(n432) );
  MXI2X1 U436 ( .A(n460), .B(n455), .S0(n332), .Y(n443) );
  MXI2X1 U437 ( .A(n462), .B(n459), .S0(n332), .Y(n445) );
  NOR3X1 U438 ( .A(n470), .B(n347), .C(n326), .Y(B[10]) );
  MX3XL U439 ( .A(n354), .B(n404), .C(n414), .S0(n338), .S1(n343), .Y(n470) );
  MXI2X1 U440 ( .A(n471), .B(n472), .S0(n332), .Y(n450) );
  MXI2X1 U441 ( .A(n451), .B(n449), .S0(n334), .Y(n434) );
  MXI2X1 U442 ( .A(n478), .B(n479), .S0(n332), .Y(n449) );
  MXI2X1 U443 ( .A(n480), .B(n481), .S0(n332), .Y(n451) );
  NOR3X1 U444 ( .A(n482), .B(n347), .C(n326), .Y(B[0]) );
  AND4X1 U445 ( .A(n487), .B(n488), .C(n489), .D(n490), .Y(n486) );
  NOR3X1 U446 ( .A(SH[29]), .B(SH[31]), .C(SH[30]), .Y(n489) );
  NOR3X1 U447 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n484) );
  MX3XL U448 ( .A(n367), .B(n492), .C(n439), .S0(n338), .S1(n343), .Y(n482) );
  MXI2X1 U449 ( .A(n416), .B(n369), .S0(n338), .Y(n439) );
  MXI2X1 U450 ( .A(n468), .B(n465), .S0(n334), .Y(n369) );
  MXI2X1 U451 ( .A(n479), .B(n474), .S0(n332), .Y(n465) );
  MXI2X1 U452 ( .A(n481), .B(n478), .S0(n332), .Y(n468) );
  MXI2X1 U453 ( .A(n472), .B(n480), .S0(n332), .Y(n467) );
  MXI2X1 U454 ( .A(n391), .B(n493), .S0(n334), .Y(n492) );
  MX3XL U455 ( .A(A[1]), .B(A[0]), .C(n361), .S0(n330), .S1(SH[1]), .Y(n493)
         );
  MXI2X1 U456 ( .A(A[5]), .B(A[4]), .S0(n329), .Y(n407) );
  MXI2X1 U457 ( .A(n475), .B(n476), .S0(n332), .Y(n466) );
  MXI2X1 U458 ( .A(n477), .B(n409), .S0(n332), .Y(n393) );
endmodule


module ALU_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n36, n38, n39, n40, n41, n42, n44, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n60, n62, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n133,
         n134, n135, n136, n138, n139, n140, n141, n142, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n208, n210, n212, n213, n214, n216, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394;

  AOI21X1 U304 ( .A0(n140), .A1(n127), .B0(n128), .Y(n126) );
  OAI21X2 U305 ( .A0(n99), .A1(n87), .B0(n88), .Y(n86) );
  INVX1 U306 ( .A(n99), .Y(n98) );
  NOR2X2 U307 ( .A(n251), .B(A[17]), .Y(n114) );
  OAI21X2 U308 ( .A0(n122), .A1(n48), .B0(n49), .Y(n47) );
  AOI21X2 U309 ( .A0(n121), .A1(n73), .B0(n74), .Y(n72) );
  CLKINVX8 U310 ( .A(n122), .Y(n121) );
  NOR2X1 U311 ( .A(n169), .B(n166), .Y(n164) );
  NOR2X2 U312 ( .A(n259), .B(A[9]), .Y(n166) );
  NOR2X1 U313 ( .A(n246), .B(A[22]), .Y(n84) );
  NOR2X2 U314 ( .A(n255), .B(A[13]), .Y(n141) );
  INVXL U315 ( .A(n185), .Y(n232) );
  OAI21X2 U316 ( .A0(n185), .A1(n191), .B0(n186), .Y(n184) );
  OAI21X1 U317 ( .A0(n171), .A1(n162), .B0(n163), .Y(n161) );
  INVX2 U318 ( .A(n172), .Y(n171) );
  NOR2X2 U319 ( .A(n243), .B(A[25]), .Y(n66) );
  INVX1 U320 ( .A(B[25]), .Y(n243) );
  INVX3 U321 ( .A(n199), .Y(n371) );
  CLKINVX4 U322 ( .A(n371), .Y(n372) );
  BUFX3 U323 ( .A(n197), .Y(n373) );
  CLKBUFX3 U324 ( .A(n177), .Y(n374) );
  NOR2X2 U325 ( .A(n129), .B(n134), .Y(n127) );
  NOR2X1 U326 ( .A(n254), .B(A[14]), .Y(n134) );
  NOR2X2 U327 ( .A(n146), .B(n141), .Y(n139) );
  NOR2X1 U328 ( .A(n256), .B(A[12]), .Y(n146) );
  INVX4 U329 ( .A(B[17]), .Y(n251) );
  BUFX6 U330 ( .A(n149), .Y(n375) );
  NOR2X4 U331 ( .A(n392), .B(A[3]), .Y(n196) );
  INVX2 U332 ( .A(B[3]), .Y(n392) );
  INVX8 U333 ( .A(B[5]), .Y(n394) );
  CLKINVX1 U334 ( .A(B[24]), .Y(n244) );
  AOI21X2 U335 ( .A0(n90), .A1(n77), .B0(n78), .Y(n76) );
  OAI21X1 U336 ( .A0(n91), .A1(n97), .B0(n92), .Y(n90) );
  INVX6 U337 ( .A(B[9]), .Y(n259) );
  INVX8 U338 ( .A(B[7]), .Y(n261) );
  NOR2X1 U339 ( .A(n390), .B(A[1]), .Y(n203) );
  INVX6 U340 ( .A(B[1]), .Y(n390) );
  NAND2X4 U341 ( .A(n262), .B(A[6]), .Y(n181) );
  INVX4 U342 ( .A(B[6]), .Y(n262) );
  NOR2X4 U343 ( .A(n159), .B(n154), .Y(n152) );
  NOR2X2 U344 ( .A(n257), .B(A[11]), .Y(n154) );
  NAND2X1 U345 ( .A(n391), .B(A[2]), .Y(n200) );
  INVX8 U346 ( .A(B[2]), .Y(n391) );
  INVXL U347 ( .A(n140), .Y(n138) );
  OAI21X1 U348 ( .A0(n141), .A1(n147), .B0(n142), .Y(n140) );
  NAND2X2 U349 ( .A(n104), .B(n112), .Y(n102) );
  NOR2X2 U350 ( .A(n102), .B(n75), .Y(n73) );
  NAND2X4 U351 ( .A(n376), .B(n138), .Y(n136) );
  NAND2XL U352 ( .A(n375), .B(n139), .Y(n376) );
  OAI21XL U353 ( .A0(n111), .A1(n109), .B0(n110), .Y(n108) );
  CLKINVX1 U354 ( .A(B[23]), .Y(n245) );
  CLKINVX1 U355 ( .A(B[22]), .Y(n246) );
  OAI21X1 U356 ( .A0(n66), .A1(n70), .B0(n67), .Y(n65) );
  AOI21X2 U357 ( .A0(n202), .A1(n194), .B0(n195), .Y(n193) );
  NAND2X1 U358 ( .A(n377), .B(n373), .Y(n195) );
  NOR2X1 U359 ( .A(n393), .B(A[4]), .Y(n190) );
  CLKINVX1 U360 ( .A(B[8]), .Y(n260) );
  CLKINVX1 U361 ( .A(B[11]), .Y(n257) );
  CLKINVX1 U362 ( .A(B[12]), .Y(n256) );
  CLKINVX1 U363 ( .A(B[13]), .Y(n255) );
  CLKINVX1 U364 ( .A(B[16]), .Y(n252) );
  AOI21X1 U365 ( .A0(n121), .A1(n100), .B0(n101), .Y(n99) );
  CLKINVX1 U366 ( .A(B[21]), .Y(n247) );
  CLKINVX1 U367 ( .A(B[19]), .Y(n249) );
  CLKINVX1 U368 ( .A(B[18]), .Y(n250) );
  AO21X1 U369 ( .A0(n136), .A1(n223), .B0(n133), .Y(n383) );
  CLKINVX1 U370 ( .A(n193), .Y(n192) );
  NOR2X1 U371 ( .A(n391), .B(A[2]), .Y(n199) );
  AOI21X1 U372 ( .A0(n192), .A1(n183), .B0(n184), .Y(n182) );
  CLKINVX1 U373 ( .A(n72), .Y(n71) );
  XNOR2X1 U374 ( .A(n136), .B(n18), .Y(DIFF[14]) );
  AOI21X1 U375 ( .A0(n39), .A1(n385), .B0(n36), .Y(n34) );
  OAI21X1 U376 ( .A0(n166), .A1(n170), .B0(n167), .Y(n165) );
  NOR2X1 U377 ( .A(n247), .B(A[21]), .Y(n91) );
  AOI21X1 U378 ( .A0(n121), .A1(n112), .B0(n113), .Y(n111) );
  CLKINVX1 U379 ( .A(n375), .Y(n148) );
  NAND2X4 U380 ( .A(n378), .B(n41), .Y(n39) );
  NAND2X1 U381 ( .A(n239), .B(A[29]), .Y(n41) );
  NOR2X1 U382 ( .A(n241), .B(A[27]), .Y(n52) );
  CLKINVX1 U383 ( .A(B[27]), .Y(n241) );
  AOI21X4 U384 ( .A0(n165), .A1(n152), .B0(n153), .Y(n151) );
  OAI21X2 U385 ( .A0(n151), .A1(n125), .B0(n126), .Y(n124) );
  NAND2X1 U386 ( .A(n393), .B(A[4]), .Y(n191) );
  OAI21X4 U387 ( .A0(n193), .A1(n173), .B0(n174), .Y(n172) );
  NAND2X2 U388 ( .A(n89), .B(n77), .Y(n75) );
  INVX1 U389 ( .A(B[20]), .Y(n248) );
  NAND2X1 U390 ( .A(n256), .B(A[12]), .Y(n147) );
  XNOR2X4 U391 ( .A(n108), .B(n13), .Y(DIFF[19]) );
  XNOR2X2 U392 ( .A(n71), .B(n8), .Y(DIFF[24]) );
  NAND2X2 U393 ( .A(n260), .B(A[8]), .Y(n170) );
  NAND2X1 U394 ( .A(n250), .B(A[18]), .Y(n110) );
  XOR2X1 U395 ( .A(n42), .B(n3), .Y(DIFF[29]) );
  NAND2X1 U396 ( .A(n164), .B(n152), .Y(n150) );
  NOR2X1 U397 ( .A(n258), .B(A[10]), .Y(n159) );
  NOR2X1 U398 ( .A(n245), .B(A[23]), .Y(n79) );
  OR2X2 U399 ( .A(n196), .B(n200), .Y(n377) );
  OR2X8 U400 ( .A(n42), .B(n40), .Y(n378) );
  AOI21X2 U401 ( .A0(n47), .A1(n387), .B0(n44), .Y(n42) );
  XNOR2X4 U402 ( .A(n39), .B(n2), .Y(DIFF[30]) );
  NOR2X1 U403 ( .A(n261), .B(A[7]), .Y(n177) );
  NAND2XL U404 ( .A(n245), .B(A[23]), .Y(n80) );
  NOR2X1 U405 ( .A(n249), .B(A[19]), .Y(n106) );
  OAI21X2 U406 ( .A0(n114), .A1(n120), .B0(n115), .Y(n113) );
  NAND2X1 U407 ( .A(n252), .B(A[16]), .Y(n120) );
  AOI21X2 U408 ( .A0(n172), .A1(n123), .B0(n124), .Y(n122) );
  OAI21X2 U409 ( .A0(n154), .A1(n160), .B0(n155), .Y(n153) );
  NAND2XL U410 ( .A(n231), .B(n181), .Y(n26) );
  OAI21X1 U411 ( .A0(n374), .A1(n181), .B0(n178), .Y(n176) );
  NOR2X2 U412 ( .A(n66), .B(n69), .Y(n64) );
  OAI21XL U413 ( .A0(n79), .A1(n85), .B0(n80), .Y(n78) );
  NAND2XL U414 ( .A(n255), .B(A[13]), .Y(n142) );
  INVXL U415 ( .A(B[10]), .Y(n258) );
  NOR2X1 U416 ( .A(n150), .B(n125), .Y(n123) );
  INVXL U417 ( .A(n58), .Y(n56) );
  INVXL U418 ( .A(n180), .Y(n231) );
  AO21X1 U419 ( .A0(n71), .A1(n64), .B0(n65), .Y(n380) );
  INVXL U420 ( .A(n203), .Y(n236) );
  INVXL U421 ( .A(B[15]), .Y(n253) );
  INVXL U422 ( .A(n89), .Y(n87) );
  INVX1 U423 ( .A(n90), .Y(n88) );
  NAND2X2 U424 ( .A(n139), .B(n127), .Y(n125) );
  INVXL U425 ( .A(n102), .Y(n100) );
  INVXL U426 ( .A(n103), .Y(n101) );
  XNOR2X1 U427 ( .A(n379), .B(n19), .Y(DIFF[13]) );
  AO21XL U428 ( .A0(n375), .A1(n225), .B0(n145), .Y(n379) );
  INVXL U429 ( .A(n202), .Y(n201) );
  INVXL U430 ( .A(n57), .Y(n55) );
  OAI21X1 U431 ( .A0(n58), .A1(n52), .B0(n53), .Y(n51) );
  NAND2XL U432 ( .A(n223), .B(n135), .Y(n18) );
  XNOR2XL U433 ( .A(n161), .B(n22), .Y(DIFF[10]) );
  XNOR2X1 U434 ( .A(n380), .B(n6), .Y(DIFF[26]) );
  XNOR2X1 U435 ( .A(n381), .B(n9), .Y(DIFF[23]) );
  AO21X1 U436 ( .A0(n86), .A1(n82), .B0(n83), .Y(n381) );
  XOR2XL U437 ( .A(n148), .B(n20), .Y(DIFF[12]) );
  XOR2XL U438 ( .A(n111), .B(n14), .Y(DIFF[18]) );
  NAND2XL U439 ( .A(n219), .B(n110), .Y(n14) );
  INVXL U440 ( .A(n109), .Y(n219) );
  INVXL U441 ( .A(n91), .Y(n216) );
  XNOR2X1 U442 ( .A(n382), .B(n15), .Y(DIFF[17]) );
  AO21XL U443 ( .A0(n121), .A1(n221), .B0(n118), .Y(n382) );
  NAND2XL U444 ( .A(n226), .B(n155), .Y(n21) );
  INVXL U445 ( .A(n154), .Y(n226) );
  XNOR2X1 U446 ( .A(n383), .B(n17), .Y(DIFF[15]) );
  INVXL U447 ( .A(n69), .Y(n213) );
  XNOR2XL U448 ( .A(n47), .B(n4), .Y(DIFF[28]) );
  XNOR2XL U449 ( .A(n98), .B(n12), .Y(DIFF[20]) );
  NAND2XL U450 ( .A(n94), .B(n97), .Y(n12) );
  XNOR2XL U451 ( .A(n121), .B(n16), .Y(DIFF[16]) );
  NAND2XL U452 ( .A(n238), .B(A[30]), .Y(n38) );
  XOR2XL U453 ( .A(n31), .B(n205), .Y(DIFF[1]) );
  INVXL U454 ( .A(n134), .Y(n223) );
  OR2XL U455 ( .A(n238), .B(A[30]), .Y(n385) );
  XOR2XL U456 ( .A(n171), .B(n24), .Y(DIFF[8]) );
  INVXL U457 ( .A(n169), .Y(n229) );
  XOR2XL U458 ( .A(n182), .B(n26), .Y(DIFF[6]) );
  XOR2XL U459 ( .A(n201), .B(n30), .Y(DIFF[2]) );
  NAND2XL U460 ( .A(n235), .B(n200), .Y(n30) );
  INVXL U461 ( .A(n372), .Y(n235) );
  XNOR2X1 U462 ( .A(n384), .B(n27), .Y(DIFF[5]) );
  AO21XL U463 ( .A0(n192), .A1(n233), .B0(n189), .Y(n384) );
  XNOR2XL U464 ( .A(n192), .B(n28), .Y(DIFF[4]) );
  INVXL U465 ( .A(n166), .Y(n228) );
  INVXL U466 ( .A(n196), .Y(n234) );
  INVXL U467 ( .A(n96), .Y(n94) );
  INVXL U468 ( .A(n97), .Y(n95) );
  NAND2XL U469 ( .A(n258), .B(A[10]), .Y(n160) );
  NAND2XL U470 ( .A(n246), .B(A[22]), .Y(n85) );
  OR2XL U471 ( .A(n242), .B(A[26]), .Y(n386) );
  NAND2XL U472 ( .A(n244), .B(A[24]), .Y(n70) );
  NOR2XL U473 ( .A(n252), .B(A[16]), .Y(n119) );
  NOR2X1 U474 ( .A(n394), .B(A[5]), .Y(n185) );
  NAND2XL U475 ( .A(n247), .B(A[21]), .Y(n92) );
  NAND2XL U476 ( .A(n394), .B(A[5]), .Y(n186) );
  NAND2XL U477 ( .A(n259), .B(A[9]), .Y(n167) );
  NAND2XL U478 ( .A(n390), .B(A[1]), .Y(n204) );
  NOR2X1 U479 ( .A(n262), .B(A[6]), .Y(n180) );
  NAND2XL U480 ( .A(n392), .B(A[3]), .Y(n197) );
  NAND2XL U481 ( .A(n261), .B(A[7]), .Y(n178) );
  NAND2XL U482 ( .A(n249), .B(A[19]), .Y(n107) );
  NAND2XL U483 ( .A(n237), .B(A[31]), .Y(n33) );
  INVX1 U484 ( .A(B[14]), .Y(n254) );
  NOR2XL U485 ( .A(n239), .B(A[29]), .Y(n40) );
  XNOR2XL U486 ( .A(n389), .B(A[0]), .Y(DIFF[0]) );
  NAND2XL U487 ( .A(n240), .B(A[28]), .Y(n46) );
  NAND2XL U488 ( .A(n241), .B(A[27]), .Y(n53) );
  OR2XL U489 ( .A(n240), .B(A[28]), .Y(n387) );
  INVXL U490 ( .A(B[28]), .Y(n240) );
  INVXL U491 ( .A(B[30]), .Y(n238) );
  INVXL U492 ( .A(B[29]), .Y(n239) );
  INVXL U493 ( .A(B[31]), .Y(n237) );
  OR2XL U494 ( .A(n237), .B(A[31]), .Y(n388) );
  OAI21X1 U495 ( .A0(n171), .A1(n150), .B0(n151), .Y(n149) );
  NAND2X1 U496 ( .A(n385), .B(n38), .Y(n2) );
  NAND2X1 U497 ( .A(n224), .B(n142), .Y(n19) );
  CLKINVX1 U498 ( .A(n141), .Y(n224) );
  CLKINVX1 U499 ( .A(n164), .Y(n162) );
  CLKINVX1 U500 ( .A(n165), .Y(n163) );
  CLKINVX1 U501 ( .A(n38), .Y(n36) );
  CLKINVX1 U502 ( .A(n46), .Y(n44) );
  AOI21X1 U503 ( .A0(n65), .A1(n386), .B0(n60), .Y(n58) );
  CLKINVX1 U504 ( .A(n62), .Y(n60) );
  AOI21X1 U505 ( .A0(n113), .A1(n104), .B0(n105), .Y(n103) );
  OAI21XL U506 ( .A0(n106), .A1(n110), .B0(n107), .Y(n105) );
  NAND2X1 U507 ( .A(n183), .B(n175), .Y(n173) );
  AOI21X1 U508 ( .A0(n184), .A1(n175), .B0(n176), .Y(n174) );
  NOR2X1 U509 ( .A(n374), .B(n180), .Y(n175) );
  NOR2X1 U510 ( .A(n372), .B(n196), .Y(n194) );
  OAI21X1 U511 ( .A0(n103), .A1(n75), .B0(n76), .Y(n74) );
  NAND2X1 U512 ( .A(n73), .B(n50), .Y(n48) );
  AOI21X1 U513 ( .A0(n74), .A1(n50), .B0(n51), .Y(n49) );
  NOR2X1 U514 ( .A(n57), .B(n52), .Y(n50) );
  NOR2X1 U515 ( .A(n119), .B(n114), .Y(n112) );
  NOR2X1 U516 ( .A(n106), .B(n109), .Y(n104) );
  XNOR2X1 U517 ( .A(n68), .B(n7), .Y(DIFF[25]) );
  OAI21XL U518 ( .A0(n72), .A1(n69), .B0(n70), .Y(n68) );
  NAND2X1 U519 ( .A(n64), .B(n386), .Y(n57) );
  NAND2X1 U520 ( .A(n221), .B(n120), .Y(n16) );
  NAND2X1 U521 ( .A(n387), .B(n46), .Y(n4) );
  NAND2X1 U522 ( .A(n213), .B(n70), .Y(n8) );
  XNOR2X1 U523 ( .A(n86), .B(n10), .Y(DIFF[22]) );
  NAND2X1 U524 ( .A(n82), .B(n85), .Y(n10) );
  NAND2X1 U525 ( .A(n218), .B(n107), .Y(n13) );
  CLKINVX1 U526 ( .A(n106), .Y(n218) );
  OAI21XL U527 ( .A0(n129), .A1(n135), .B0(n130), .Y(n128) );
  XOR2X1 U528 ( .A(n54), .B(n5), .Y(DIFF[27]) );
  NAND2X1 U529 ( .A(n210), .B(n53), .Y(n5) );
  AOI21X1 U530 ( .A0(n71), .A1(n55), .B0(n56), .Y(n54) );
  CLKINVX1 U531 ( .A(n52), .Y(n210) );
  NAND2X1 U532 ( .A(n214), .B(n80), .Y(n9) );
  CLKINVX1 U533 ( .A(n79), .Y(n214) );
  NAND2X1 U534 ( .A(n208), .B(n41), .Y(n3) );
  CLKINVX1 U535 ( .A(n40), .Y(n208) );
  XOR2X1 U536 ( .A(n93), .B(n11), .Y(DIFF[21]) );
  NAND2X1 U537 ( .A(n216), .B(n92), .Y(n11) );
  AOI21X1 U538 ( .A0(n98), .A1(n94), .B0(n95), .Y(n93) );
  NAND2X1 U539 ( .A(n220), .B(n115), .Y(n15) );
  CLKINVX1 U540 ( .A(n114), .Y(n220) );
  NAND2X1 U541 ( .A(n386), .B(n62), .Y(n6) );
  NAND2X1 U542 ( .A(n222), .B(n130), .Y(n17) );
  CLKINVX1 U543 ( .A(n129), .Y(n222) );
  OAI21X1 U544 ( .A0(n203), .A1(n205), .B0(n204), .Y(n202) );
  INVXL U545 ( .A(n135), .Y(n133) );
  NOR2X1 U546 ( .A(n91), .B(n96), .Y(n89) );
  NAND2X1 U547 ( .A(n227), .B(n160), .Y(n22) );
  XNOR2X1 U548 ( .A(n168), .B(n23), .Y(DIFF[9]) );
  NAND2X1 U549 ( .A(n228), .B(n167), .Y(n23) );
  OAI21XL U550 ( .A0(n171), .A1(n169), .B0(n170), .Y(n168) );
  NAND2X1 U551 ( .A(n233), .B(n191), .Y(n28) );
  CLKINVX1 U552 ( .A(n119), .Y(n221) );
  CLKINVX1 U553 ( .A(n159), .Y(n227) );
  CLKINVX1 U554 ( .A(n84), .Y(n82) );
  NOR2X1 U555 ( .A(n84), .B(n79), .Y(n77) );
  XNOR2X1 U556 ( .A(n198), .B(n29), .Y(DIFF[3]) );
  NAND2X1 U557 ( .A(n234), .B(n373), .Y(n29) );
  OAI21XL U558 ( .A0(n201), .A1(n372), .B0(n200), .Y(n198) );
  NAND2X1 U559 ( .A(n232), .B(n186), .Y(n27) );
  NOR2X1 U560 ( .A(n190), .B(n185), .Y(n183) );
  XNOR2X1 U561 ( .A(n179), .B(n25), .Y(DIFF[7]) );
  NAND2X1 U562 ( .A(n230), .B(n178), .Y(n25) );
  OAI21XL U563 ( .A0(n182), .A1(n180), .B0(n181), .Y(n179) );
  CLKINVX1 U564 ( .A(n374), .Y(n230) );
  CLKINVX1 U565 ( .A(n190), .Y(n233) );
  CLKINVX1 U566 ( .A(n146), .Y(n225) );
  CLKINVX1 U567 ( .A(n120), .Y(n118) );
  CLKINVX1 U568 ( .A(n160), .Y(n158) );
  CLKINVX1 U569 ( .A(n85), .Y(n83) );
  NAND2X1 U570 ( .A(n236), .B(n204), .Y(n31) );
  CLKINVX1 U571 ( .A(n191), .Y(n189) );
  CLKINVX1 U572 ( .A(n147), .Y(n145) );
  XOR2X1 U573 ( .A(n156), .B(n21), .Y(DIFF[11]) );
  AOI21X1 U574 ( .A0(n161), .A1(n227), .B0(n158), .Y(n156) );
  NAND2X1 U575 ( .A(n225), .B(n147), .Y(n20) );
  NAND2X1 U576 ( .A(n229), .B(n170), .Y(n24) );
  CLKINVX1 U577 ( .A(B[4]), .Y(n393) );
  NOR2X1 U578 ( .A(n244), .B(A[24]), .Y(n69) );
  XOR2X1 U579 ( .A(n34), .B(n1), .Y(DIFF[31]) );
  NAND2X1 U580 ( .A(n388), .B(n33), .Y(n1) );
  NAND2X1 U581 ( .A(n253), .B(A[15]), .Y(n130) );
  NOR2X1 U582 ( .A(n389), .B(A[0]), .Y(n205) );
  CLKINVX1 U583 ( .A(B[26]), .Y(n242) );
  CLKINVX1 U584 ( .A(B[0]), .Y(n389) );
  NAND2X1 U585 ( .A(n212), .B(n67), .Y(n7) );
  INVXL U586 ( .A(n66), .Y(n212) );
  NOR2X1 U587 ( .A(n248), .B(A[20]), .Y(n96) );
  NAND2X1 U588 ( .A(n248), .B(A[20]), .Y(n97) );
  NAND2XL U589 ( .A(n243), .B(A[25]), .Y(n67) );
  NAND2XL U590 ( .A(n254), .B(A[14]), .Y(n135) );
  NAND2X1 U591 ( .A(n242), .B(A[26]), .Y(n62) );
  NOR2X1 U592 ( .A(n250), .B(A[18]), .Y(n109) );
  NAND2X1 U593 ( .A(n257), .B(A[11]), .Y(n155) );
  NAND2X1 U594 ( .A(n251), .B(A[17]), .Y(n115) );
  NOR2X2 U595 ( .A(n260), .B(A[8]), .Y(n169) );
  NOR2X2 U596 ( .A(n253), .B(A[15]), .Y(n129) );
endmodule


module ALU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n37, n39, n40, n41, n42, n43, n45, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n210, n212, n214, n215, n216,
         n218, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357;

  OAI21X1 U275 ( .A0(n92), .A1(n98), .B0(n93), .Y(n91) );
  OAI21X1 U276 ( .A0(n172), .A1(n163), .B0(n164), .Y(n162) );
  INVX3 U277 ( .A(n173), .Y(n172) );
  INVX1 U278 ( .A(n194), .Y(n193) );
  AOI21X2 U279 ( .A0(n203), .A1(n195), .B0(n196), .Y(n194) );
  AOI21X2 U280 ( .A0(n122), .A1(n101), .B0(n102), .Y(n100) );
  CLKBUFX3 U281 ( .A(n85), .Y(n342) );
  NOR2X2 U282 ( .A(n343), .B(n155), .Y(n153) );
  OAI21X2 U283 ( .A0(n155), .A1(n161), .B0(n156), .Y(n154) );
  NOR2X2 U284 ( .A(B[11]), .B(A[11]), .Y(n155) );
  AOI21X2 U285 ( .A0(n66), .A1(n351), .B0(n61), .Y(n59) );
  OAI21X1 U286 ( .A0(n67), .A1(n71), .B0(n68), .Y(n66) );
  OAI21X2 U287 ( .A0(n142), .A1(n148), .B0(n143), .Y(n141) );
  NOR2X2 U288 ( .A(B[13]), .B(A[13]), .Y(n142) );
  NAND2X2 U289 ( .A(n74), .B(n51), .Y(n49) );
  NOR2X2 U290 ( .A(n58), .B(n53), .Y(n51) );
  BUFX3 U291 ( .A(n160), .Y(n343) );
  BUFX8 U292 ( .A(n197), .Y(n344) );
  OAI21X2 U293 ( .A0(n186), .A1(n192), .B0(n187), .Y(n185) );
  NAND2X2 U294 ( .A(n357), .B(A[4]), .Y(n192) );
  BUFX6 U295 ( .A(n171), .Y(n345) );
  OAI21X2 U296 ( .A0(n172), .A1(n151), .B0(n152), .Y(n150) );
  NAND2X1 U297 ( .A(n105), .B(n113), .Y(n103) );
  XNOR2X2 U298 ( .A(n48), .B(n4), .Y(SUM[28]) );
  NOR2X1 U299 ( .A(n130), .B(n135), .Y(n128) );
  CLKBUFX3 U300 ( .A(B[4]), .Y(n357) );
  OAI21X2 U301 ( .A0(n194), .A1(n174), .B0(n175), .Y(n173) );
  AOI21X1 U302 ( .A0(n166), .A1(n153), .B0(n154), .Y(n152) );
  NOR2X1 U303 ( .A(B[12]), .B(A[12]), .Y(n147) );
  NOR2X1 U304 ( .A(B[16]), .B(A[16]), .Y(n120) );
  NOR2X1 U305 ( .A(n103), .B(n76), .Y(n74) );
  NOR2X1 U306 ( .A(B[15]), .B(A[15]), .Y(n130) );
  NOR2X1 U307 ( .A(B[5]), .B(A[5]), .Y(n186) );
  NOR2X1 U308 ( .A(B[23]), .B(A[23]), .Y(n80) );
  NAND2X1 U309 ( .A(B[18]), .B(A[18]), .Y(n111) );
  NOR2X1 U310 ( .A(B[18]), .B(A[18]), .Y(n110) );
  NOR2X1 U311 ( .A(n67), .B(n70), .Y(n65) );
  NOR2X1 U312 ( .A(n356), .B(A[3]), .Y(n197) );
  NOR2X1 U313 ( .A(B[2]), .B(A[2]), .Y(n200) );
  NOR2X1 U314 ( .A(B[8]), .B(A[8]), .Y(n170) );
  NOR2X1 U315 ( .A(B[7]), .B(A[7]), .Y(n178) );
  AOI21X1 U316 ( .A0(n193), .A1(n184), .B0(n185), .Y(n183) );
  NAND2X1 U317 ( .A(B[16]), .B(A[16]), .Y(n121) );
  CLKINVX1 U318 ( .A(n100), .Y(n99) );
  NOR2X1 U319 ( .A(B[25]), .B(A[25]), .Y(n67) );
  NAND2X1 U320 ( .A(B[25]), .B(A[25]), .Y(n68) );
  NOR2X1 U321 ( .A(B[9]), .B(A[9]), .Y(n167) );
  NOR2X1 U322 ( .A(n357), .B(A[4]), .Y(n191) );
  NAND2X1 U323 ( .A(B[17]), .B(A[17]), .Y(n116) );
  NOR2X2 U324 ( .A(B[17]), .B(A[17]), .Y(n115) );
  XNOR2X2 U325 ( .A(n72), .B(n8), .Y(SUM[24]) );
  AOI21X4 U326 ( .A0(n122), .A1(n113), .B0(n114), .Y(n112) );
  INVX8 U327 ( .A(n123), .Y(n122) );
  XNOR2X1 U328 ( .A(n99), .B(n12), .Y(SUM[20]) );
  NOR2X1 U329 ( .A(n151), .B(n126), .Y(n124) );
  XOR2X4 U330 ( .A(n64), .B(n6), .Y(SUM[26]) );
  AOI21X2 U331 ( .A0(n72), .A1(n65), .B0(n66), .Y(n64) );
  OAI21X1 U332 ( .A0(n152), .A1(n126), .B0(n127), .Y(n125) );
  OR2XL U333 ( .A(n123), .B(n49), .Y(n346) );
  NAND2X2 U334 ( .A(n346), .B(n50), .Y(n48) );
  AOI21X1 U335 ( .A0(n75), .A1(n51), .B0(n52), .Y(n50) );
  AOI21X4 U336 ( .A0(n48), .A1(n353), .B0(n45), .Y(n43) );
  AOI21X4 U337 ( .A0(n173), .A1(n124), .B0(n125), .Y(n123) );
  OAI21X1 U338 ( .A0(n344), .A1(n201), .B0(n198), .Y(n196) );
  NAND2X1 U339 ( .A(B[2]), .B(A[2]), .Y(n201) );
  BUFX4 U340 ( .A(n87), .Y(n347) );
  NOR2X1 U341 ( .A(B[14]), .B(A[14]), .Y(n135) );
  AOI21X4 U342 ( .A0(n40), .A1(n352), .B0(n37), .Y(n35) );
  OAI21X4 U343 ( .A0(n43), .A1(n41), .B0(n42), .Y(n40) );
  NAND2X1 U344 ( .A(n356), .B(A[3]), .Y(n198) );
  AOI21X2 U345 ( .A0(n347), .A1(n83), .B0(n84), .Y(n82) );
  XNOR2X1 U346 ( .A(n347), .B(n10), .Y(SUM[22]) );
  OAI21X2 U347 ( .A0(n204), .A1(n207), .B0(n205), .Y(n203) );
  NOR2X1 U348 ( .A(B[1]), .B(A[1]), .Y(n204) );
  OAI21X4 U349 ( .A0(n149), .A1(n138), .B0(n139), .Y(n137) );
  INVX3 U350 ( .A(n150), .Y(n149) );
  NOR2X1 U351 ( .A(n120), .B(n115), .Y(n113) );
  NAND2XL U352 ( .A(B[13]), .B(A[13]), .Y(n143) );
  NAND2X1 U353 ( .A(n165), .B(n153), .Y(n151) );
  INVXL U354 ( .A(n103), .Y(n101) );
  INVXL U355 ( .A(n58), .Y(n56) );
  XNOR2X1 U356 ( .A(n40), .B(n2), .Y(SUM[30]) );
  INVXL U357 ( .A(n70), .Y(n215) );
  NAND2XL U358 ( .A(n355), .B(A[0]), .Y(n207) );
  INVX3 U359 ( .A(n73), .Y(n72) );
  INVXL U360 ( .A(n90), .Y(n88) );
  INVXL U361 ( .A(n91), .Y(n89) );
  INVXL U362 ( .A(n104), .Y(n102) );
  INVXL U363 ( .A(n59), .Y(n57) );
  NAND2XL U364 ( .A(n225), .B(n136), .Y(n18) );
  NAND2XL U365 ( .A(n221), .B(n111), .Y(n14) );
  INVXL U366 ( .A(n110), .Y(n221) );
  INVXL U367 ( .A(n80), .Y(n216) );
  NAND2XL U368 ( .A(n351), .B(n63), .Y(n6) );
  NAND2XL U369 ( .A(n224), .B(n131), .Y(n17) );
  INVXL U370 ( .A(n130), .Y(n224) );
  XNOR2X1 U371 ( .A(n348), .B(n15), .Y(SUM[17]) );
  AO21XL U372 ( .A0(n122), .A1(n223), .B0(n119), .Y(n348) );
  NAND2XL U373 ( .A(n228), .B(n156), .Y(n21) );
  INVXL U374 ( .A(n155), .Y(n228) );
  NAND2XL U375 ( .A(n95), .B(n98), .Y(n12) );
  XNOR2XL U376 ( .A(n122), .B(n16), .Y(SUM[16]) );
  NAND2XL U377 ( .A(n229), .B(n161), .Y(n22) );
  XOR2XL U378 ( .A(n149), .B(n20), .Y(SUM[12]) );
  XOR2XL U379 ( .A(n172), .B(n24), .Y(SUM[8]) );
  INVXL U380 ( .A(n170), .Y(n231) );
  XOR2XL U381 ( .A(n202), .B(n30), .Y(SUM[2]) );
  INVXL U382 ( .A(n200), .Y(n237) );
  XNOR2X1 U383 ( .A(n349), .B(n19), .Y(SUM[13]) );
  AO21XL U384 ( .A0(n150), .A1(n227), .B0(n146), .Y(n349) );
  XNOR2X1 U385 ( .A(n350), .B(n27), .Y(SUM[5]) );
  AO21XL U386 ( .A0(n193), .A1(n235), .B0(n190), .Y(n350) );
  XNOR2XL U387 ( .A(n193), .B(n28), .Y(SUM[4]) );
  INVXL U388 ( .A(n167), .Y(n230) );
  INVXL U389 ( .A(n178), .Y(n232) );
  INVXL U390 ( .A(n344), .Y(n236) );
  INVXL U391 ( .A(n135), .Y(n225) );
  INVXL U392 ( .A(n97), .Y(n95) );
  INVXL U393 ( .A(n98), .Y(n96) );
  NAND2XL U394 ( .A(B[12]), .B(A[12]), .Y(n148) );
  NAND2XL U395 ( .A(B[31]), .B(A[31]), .Y(n34) );
  NAND2XL U396 ( .A(B[8]), .B(A[8]), .Y(n171) );
  NAND2XL U397 ( .A(B[10]), .B(A[10]), .Y(n161) );
  NAND2XL U398 ( .A(B[22]), .B(A[22]), .Y(n86) );
  NOR2XL U399 ( .A(B[10]), .B(A[10]), .Y(n160) );
  NOR2XL U400 ( .A(B[22]), .B(A[22]), .Y(n85) );
  NAND2XL U401 ( .A(B[24]), .B(A[24]), .Y(n71) );
  NAND2XL U402 ( .A(B[6]), .B(A[6]), .Y(n182) );
  NOR2X1 U403 ( .A(B[21]), .B(A[21]), .Y(n92) );
  NOR2X1 U404 ( .A(B[19]), .B(A[19]), .Y(n107) );
  NAND2XL U405 ( .A(B[23]), .B(A[23]), .Y(n81) );
  NOR2X1 U406 ( .A(B[6]), .B(A[6]), .Y(n181) );
  NAND2XL U407 ( .A(B[9]), .B(A[9]), .Y(n168) );
  NAND2XL U408 ( .A(B[21]), .B(A[21]), .Y(n93) );
  NAND2XL U409 ( .A(B[7]), .B(A[7]), .Y(n179) );
  NAND2XL U410 ( .A(B[19]), .B(A[19]), .Y(n108) );
  NAND2XL U411 ( .A(B[5]), .B(A[5]), .Y(n187) );
  NAND2XL U412 ( .A(B[1]), .B(A[1]), .Y(n205) );
  OR2XL U413 ( .A(B[26]), .B(A[26]), .Y(n351) );
  NOR2XL U414 ( .A(B[29]), .B(A[29]), .Y(n41) );
  NAND2XL U415 ( .A(B[28]), .B(A[28]), .Y(n47) );
  NAND2XL U416 ( .A(B[30]), .B(A[30]), .Y(n39) );
  NOR2X1 U417 ( .A(B[27]), .B(A[27]), .Y(n53) );
  NAND2XL U418 ( .A(B[27]), .B(A[27]), .Y(n54) );
  NAND2XL U419 ( .A(B[29]), .B(A[29]), .Y(n42) );
  OR2XL U420 ( .A(B[28]), .B(A[28]), .Y(n353) );
  OR2XL U421 ( .A(B[30]), .B(A[30]), .Y(n352) );
  NAND2BXL U422 ( .AN(n206), .B(n207), .Y(n32) );
  NOR2XL U423 ( .A(n355), .B(A[0]), .Y(n206) );
  OR2XL U424 ( .A(B[31]), .B(A[31]), .Y(n354) );
  NAND2X1 U425 ( .A(n140), .B(n128), .Y(n126) );
  AOI21X1 U426 ( .A0(n122), .A1(n74), .B0(n75), .Y(n73) );
  CLKINVX1 U427 ( .A(n165), .Y(n163) );
  CLKINVX1 U428 ( .A(n166), .Y(n164) );
  CLKINVX1 U429 ( .A(n141), .Y(n139) );
  CLKINVX1 U430 ( .A(n140), .Y(n138) );
  OAI21XL U431 ( .A0(n100), .A1(n88), .B0(n89), .Y(n87) );
  NAND2X1 U432 ( .A(n90), .B(n78), .Y(n76) );
  CLKINVX1 U433 ( .A(n203), .Y(n202) );
  OAI21X1 U434 ( .A0(n115), .A1(n121), .B0(n116), .Y(n114) );
  XNOR2X1 U435 ( .A(n69), .B(n7), .Y(SUM[25]) );
  OAI21XL U436 ( .A0(n73), .A1(n70), .B0(n71), .Y(n69) );
  OAI21X1 U437 ( .A0(n167), .A1(n345), .B0(n168), .Y(n166) );
  CLKINVX1 U438 ( .A(n47), .Y(n45) );
  CLKINVX1 U439 ( .A(n63), .Y(n61) );
  XNOR2X1 U440 ( .A(n137), .B(n18), .Y(SUM[14]) );
  AOI21X1 U441 ( .A0(n114), .A1(n105), .B0(n106), .Y(n104) );
  OAI21XL U442 ( .A0(n107), .A1(n111), .B0(n108), .Y(n106) );
  NAND2X1 U443 ( .A(n184), .B(n176), .Y(n174) );
  AOI21X1 U444 ( .A0(n185), .A1(n176), .B0(n177), .Y(n175) );
  NOR2X1 U445 ( .A(n178), .B(n181), .Y(n176) );
  NOR2X1 U446 ( .A(n200), .B(n344), .Y(n195) );
  OAI21X1 U447 ( .A0(n104), .A1(n76), .B0(n77), .Y(n75) );
  AOI21X1 U448 ( .A0(n91), .A1(n78), .B0(n79), .Y(n77) );
  OAI21XL U449 ( .A0(n80), .A1(n86), .B0(n81), .Y(n79) );
  NAND2X1 U450 ( .A(n352), .B(n39), .Y(n2) );
  NAND2X1 U451 ( .A(n223), .B(n121), .Y(n16) );
  NAND2X1 U452 ( .A(n215), .B(n71), .Y(n8) );
  NAND2X1 U453 ( .A(n353), .B(n47), .Y(n4) );
  XNOR2X1 U454 ( .A(n180), .B(n25), .Y(SUM[7]) );
  NAND2X1 U455 ( .A(n232), .B(n179), .Y(n25) );
  OAI21XL U456 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  XNOR2X1 U457 ( .A(n109), .B(n13), .Y(SUM[19]) );
  NAND2X1 U458 ( .A(n220), .B(n108), .Y(n13) );
  OAI21XL U459 ( .A0(n112), .A1(n110), .B0(n111), .Y(n109) );
  CLKINVX1 U460 ( .A(n107), .Y(n220) );
  NAND2X1 U461 ( .A(n83), .B(n86), .Y(n10) );
  NOR2X1 U462 ( .A(n107), .B(n110), .Y(n105) );
  NOR2X1 U463 ( .A(n147), .B(n142), .Y(n140) );
  NAND2X1 U464 ( .A(n65), .B(n351), .Y(n58) );
  NOR2X1 U465 ( .A(n92), .B(n97), .Y(n90) );
  OAI21XL U466 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U467 ( .A(n170), .B(n167), .Y(n165) );
  AOI21X1 U468 ( .A0(n141), .A1(n128), .B0(n129), .Y(n127) );
  OAI21XL U469 ( .A0(n130), .A1(n136), .B0(n131), .Y(n129) );
  OAI21XL U470 ( .A0(n59), .A1(n53), .B0(n54), .Y(n52) );
  NOR2X1 U471 ( .A(n342), .B(n80), .Y(n78) );
  NAND2X1 U472 ( .A(n226), .B(n143), .Y(n19) );
  CLKINVX1 U473 ( .A(n142), .Y(n226) );
  NOR2X1 U474 ( .A(n191), .B(n186), .Y(n184) );
  XOR2X1 U475 ( .A(n55), .B(n5), .Y(SUM[27]) );
  NAND2X1 U476 ( .A(n212), .B(n54), .Y(n5) );
  AOI21X1 U477 ( .A0(n72), .A1(n56), .B0(n57), .Y(n55) );
  CLKINVX1 U478 ( .A(n53), .Y(n212) );
  XOR2X1 U479 ( .A(n94), .B(n11), .Y(SUM[21]) );
  NAND2X1 U480 ( .A(n218), .B(n93), .Y(n11) );
  AOI21X1 U481 ( .A0(n99), .A1(n95), .B0(n96), .Y(n94) );
  CLKINVX1 U482 ( .A(n92), .Y(n218) );
  NAND2X1 U483 ( .A(n222), .B(n116), .Y(n15) );
  CLKINVX1 U484 ( .A(n115), .Y(n222) );
  XOR2X1 U485 ( .A(n157), .B(n21), .Y(SUM[11]) );
  AOI21X1 U486 ( .A0(n162), .A1(n229), .B0(n159), .Y(n157) );
  NAND2X1 U487 ( .A(n227), .B(n148), .Y(n20) );
  XOR2X1 U488 ( .A(n132), .B(n17), .Y(SUM[15]) );
  AOI21X1 U489 ( .A0(n137), .A1(n225), .B0(n134), .Y(n132) );
  XOR2X1 U490 ( .A(n82), .B(n9), .Y(SUM[23]) );
  NAND2X1 U491 ( .A(n216), .B(n81), .Y(n9) );
  XOR2X1 U492 ( .A(n112), .B(n14), .Y(SUM[18]) );
  XOR2X1 U493 ( .A(n43), .B(n3), .Y(SUM[29]) );
  NAND2X1 U494 ( .A(n210), .B(n42), .Y(n3) );
  CLKINVX1 U495 ( .A(n41), .Y(n210) );
  CLKBUFX3 U496 ( .A(B[3]), .Y(n356) );
  INVXL U497 ( .A(n136), .Y(n134) );
  NAND2X1 U498 ( .A(n235), .B(n192), .Y(n28) );
  XNOR2X1 U499 ( .A(n199), .B(n29), .Y(SUM[3]) );
  NAND2X1 U500 ( .A(n236), .B(n198), .Y(n29) );
  OAI21XL U501 ( .A0(n202), .A1(n200), .B0(n201), .Y(n199) );
  XNOR2X1 U502 ( .A(n162), .B(n22), .Y(SUM[10]) );
  CLKINVX1 U503 ( .A(n120), .Y(n223) );
  CLKINVX1 U504 ( .A(n343), .Y(n229) );
  CLKINVX1 U505 ( .A(n342), .Y(n83) );
  XNOR2X1 U506 ( .A(n169), .B(n23), .Y(SUM[9]) );
  NAND2X1 U507 ( .A(n230), .B(n168), .Y(n23) );
  OAI21XL U508 ( .A0(n172), .A1(n170), .B0(n345), .Y(n169) );
  NAND2X1 U509 ( .A(n234), .B(n187), .Y(n27) );
  CLKINVX1 U510 ( .A(n186), .Y(n234) );
  CLKINVX1 U511 ( .A(n39), .Y(n37) );
  CLKINVX1 U512 ( .A(n191), .Y(n235) );
  CLKINVX1 U513 ( .A(n147), .Y(n227) );
  CLKINVX1 U514 ( .A(n121), .Y(n119) );
  CLKINVX1 U515 ( .A(n161), .Y(n159) );
  CLKINVX1 U516 ( .A(n86), .Y(n84) );
  XOR2X1 U517 ( .A(n31), .B(n207), .Y(SUM[1]) );
  NAND2X1 U518 ( .A(n238), .B(n205), .Y(n31) );
  CLKINVX1 U519 ( .A(n204), .Y(n238) );
  CLKINVX1 U520 ( .A(n192), .Y(n190) );
  NAND2X1 U521 ( .A(n237), .B(n201), .Y(n30) );
  XOR2X1 U522 ( .A(n183), .B(n26), .Y(SUM[6]) );
  NAND2X1 U523 ( .A(n233), .B(n182), .Y(n26) );
  CLKINVX1 U524 ( .A(n181), .Y(n233) );
  NAND2X1 U525 ( .A(n231), .B(n345), .Y(n24) );
  CLKINVX1 U526 ( .A(n148), .Y(n146) );
  NAND2X1 U527 ( .A(B[15]), .B(A[15]), .Y(n131) );
  XOR2X1 U528 ( .A(n35), .B(n1), .Y(SUM[31]) );
  NAND2X1 U529 ( .A(n354), .B(n34), .Y(n1) );
  CLKBUFX3 U530 ( .A(B[0]), .Y(n355) );
  NOR2X1 U531 ( .A(B[24]), .B(A[24]), .Y(n70) );
  CLKINVX1 U532 ( .A(n32), .Y(SUM[0]) );
  INVXL U533 ( .A(n67), .Y(n214) );
  NAND2X1 U534 ( .A(n214), .B(n68), .Y(n7) );
  NOR2X1 U535 ( .A(B[20]), .B(A[20]), .Y(n97) );
  NAND2X1 U536 ( .A(B[20]), .B(A[20]), .Y(n98) );
  NAND2XL U537 ( .A(B[14]), .B(A[14]), .Y(n136) );
  NAND2X1 U538 ( .A(B[26]), .B(A[26]), .Y(n63) );
  NAND2X1 U539 ( .A(B[11]), .B(A[11]), .Y(n156) );
endmodule


module ALU ( ALUOp_regD, funct_regD, ALUinA, ALUinB, ALUout );
  input [5:0] ALUOp_regD;
  input [5:0] funct_regD;
  input [31:0] ALUinA;
  input [31:0] ALUinB;
  output [31:0] ALUout;
  wire   N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N441, n110, n111, n112,
         n117, n119, n120, n130, n131, n140, n141, n150, n151, n160, n161,
         n170, n171, n180, n181, n210, n211, n290, n291, n300, n301, n310,
         n311, n320, n321, n330, n331, n340, n341, n350, n351, n360, n361,
         n370, n371, n380, n381, n390, n391, n400, n401, n410, n411, n420,
         n422, n426, n427, n429, n430, n432, n441, n442, n444, n445, n447, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n113, n114, n115, n116, n118, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n132, n133, n134,
         n135, n136, n137, n138, n139, n142, n143, n144, n145, n146, n147,
         n148, n149, n152, n153, n154, n155, n156, n157, n158, n159, n162,
         n163, n164, n165, n166, n167, n168, n169, n172, n173, n174, n175,
         n176, n177, n178, n179, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n292, n293, n294, n295, n296, n297, n298, n299, n302, n303, n304,
         n305, n306, n307, n308, n309, n312, n313, n314, n315, n316, n317,
         n318, n319, n322, n323, n324, n325, n326, n327, n328, n329, n332,
         n333, n334, n335, n336, n337, n338, n339, n342, n343, n344, n345,
         n346, n347, n348, n349, n352, n353, n354, n355, n356, n357, n358,
         n359, n362, n363, n364, n365, n366, n367, n368, n369, n372, n373,
         n374, n375, n376, n377, n378, n379, n382, n383, n384, n385, n386,
         n387, n388, n389, n392, n393, n394, n395, n396, n397, n398, n399,
         n402, n403, n404, n405, n406, n407, n408, n409, n412, n413, n414,
         n415, n416, n417, n418, n419, n421, n423, n424, n425, n428, n431,
         n433, n434, n435, n436, n437, n438, n439, n440, n443, n446, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560;

  ALU_DW_leftsh_0 sll_1160 ( .A(ALUinA), .SH({ALUinB[31:27], n4, ALUinB[25:23], 
        n56, n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, 
        n42, n41, n40, n90, n88, n86, n2, n82, n81}), .B({N376, N375, N374, 
        N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, 
        N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, 
        N349, N348, N347, N346, N345}) );
  ALU_DW_cmp_0 r323 ( .A(ALUinA), .B({ALUinB[31:27], n5, ALUinB[25:23], n56, 
        n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, n42, 
        n41, n40, n90, n88, n86, n2, n82, n81}), .TC(1'b0), .GE_LT(1'b1), 
        .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N441) );
  ALU_DW_rightsh_0 r322 ( .A(ALUinA), .DATA_TC(1'b0), .SH({ALUinB[31:27], n5, 
        ALUinB[25:23], n56, n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, 
        n45, n44, n43, n42, n41, n40, n90, n88, n86, n2, n82, n81}), .B({N408, 
        N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, 
        N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, 
        N383, N382, N381, N380, N379, N378, N377}) );
  ALU_DW01_sub_1 sub_1145 ( .A(ALUinA), .B({ALUinB[31:27], n4, ALUinB[25:23], 
        n56, n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, 
        n42, n41, n40, n90, n88, n86, n1, n82, n81}), .CI(1'b0), .DIFF({N312, 
        N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, 
        N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, 
        N287, N286, N285, N284, N283, N282, N281}) );
  ALU_DW01_add_1 r319 ( .A(ALUinA), .B({ALUinB[31:27], n4, ALUinB[25:23], n56, 
        n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, n42, 
        n41, n40, n90, n88, n86, n2, n82, n81}), .CI(1'b0), .SUM({N280, N279, 
        N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, 
        N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, 
        N254, N253, N252, N251, N250, N249}) );
  OAI221X1 U8 ( .A0(n75), .A1(n389), .B0(n388), .B1(n74), .C0(n387), .Y(
        ALUout[22]) );
  CLKBUFX20 U9 ( .A(n84), .Y(n1) );
  CLKBUFX20 U10 ( .A(n84), .Y(n2) );
  BUFX12 U11 ( .A(ALUinB[9]), .Y(n43) );
  OAI221X2 U12 ( .A0(n75), .A1(n303), .B0(n302), .B1(n74), .C0(n299), .Y(
        ALUout[15]) );
  OAI221X2 U13 ( .A0(n75), .A1(n404), .B0(n403), .B1(n74), .C0(n402), .Y(
        ALUout[23]) );
  OAI221X2 U14 ( .A0(n76), .A1(n451), .B0(n450), .B1(n74), .C0(n449), .Y(
        ALUout[26]) );
  BUFX16 U15 ( .A(ALUinB[6]), .Y(n40) );
  BUFX4 U16 ( .A(ALUinB[16]), .Y(n50) );
  CLKINVX1 U17 ( .A(ALUOp_regD[4]), .Y(n138) );
  AO22X2 U18 ( .A0(N361), .A1(n63), .B0(n361), .B1(n70), .Y(n306) );
  NOR4X1 U19 ( .A(n334), .B(n333), .C(n332), .D(n329), .Y(n338) );
  NOR4X1 U20 ( .A(n446), .B(n443), .C(n440), .D(n439), .Y(n450) );
  NOR4X2 U21 ( .A(n372), .B(n369), .C(n368), .D(n367), .Y(n376) );
  NOR4X2 U22 ( .A(n458), .B(n457), .C(n456), .D(n455), .Y(n461) );
  NOR4X2 U23 ( .A(n508), .B(n507), .C(n506), .D(n505), .Y(n513) );
  AND2X2 U24 ( .A(N249), .B(n38), .Y(n8) );
  CLKINVX1 U25 ( .A(n120), .Y(n108) );
  INVX3 U26 ( .A(n85), .Y(n84) );
  CLKINVX1 U27 ( .A(N441), .Y(n519) );
  CLKINVX1 U28 ( .A(n119), .Y(n139) );
  NAND2X1 U29 ( .A(n429), .B(ALUOp_regD[1]), .Y(n113) );
  NOR4X2 U30 ( .A(n491), .B(n490), .C(n489), .D(n488), .Y(n494) );
  AO22X1 U31 ( .A0(N311), .A1(n64), .B0(N375), .B1(n62), .Y(n490) );
  OR2X2 U32 ( .A(n352), .B(n74), .Y(n7) );
  NOR4X1 U33 ( .A(n346), .B(n345), .C(n344), .D(n343), .Y(n352) );
  AO22X1 U34 ( .A0(n330), .A1(n53), .B0(N300), .B1(n64), .Y(n345) );
  OAI221XL U35 ( .A0(n75), .A1(n339), .B0(n338), .B1(n74), .C0(n337), .Y(
        ALUout[18]) );
  OAI221XL U36 ( .A0(n75), .A1(n175), .B0(n174), .B1(n74), .C0(n173), .Y(
        ALUout[3]) );
  OAI221XL U37 ( .A0(n75), .A1(n289), .B0(n288), .B1(n74), .C0(n287), .Y(
        ALUout[14]) );
  OAI221XL U38 ( .A0(n76), .A1(n229), .B0(n228), .B1(n74), .C0(n227), .Y(
        ALUout[8]) );
  OAI221XL U39 ( .A0(n75), .A1(n187), .B0(n186), .B1(n74), .C0(n185), .Y(
        ALUout[4]) );
  OAI221X1 U40 ( .A0(n75), .A1(n417), .B0(n416), .B1(n74), .C0(n415), .Y(
        ALUout[24]) );
  OAI221XL U41 ( .A0(n76), .A1(n473), .B0(n472), .B1(n74), .C0(n471), .Y(
        ALUout[28]) );
  OAI221X1 U42 ( .A0(n76), .A1(n259), .B0(n258), .B1(n74), .C0(n257), .Y(
        ALUout[11]) );
  OAI221XL U43 ( .A0(n76), .A1(n219), .B0(n218), .B1(n74), .C0(n217), .Y(
        ALUout[7]) );
  OAI221X1 U44 ( .A0(n75), .A1(n279), .B0(n278), .B1(n74), .C0(n277), .Y(
        ALUout[13]) );
  OAI221XL U45 ( .A0(n75), .A1(n315), .B0(n314), .B1(n74), .C0(n313), .Y(
        ALUout[16]) );
  OAI221X1 U46 ( .A0(n75), .A1(n377), .B0(n376), .B1(n74), .C0(n375), .Y(
        ALUout[21]) );
  OAI221XL U47 ( .A0(n76), .A1(n484), .B0(n483), .B1(n74), .C0(n482), .Y(
        ALUout[29]) );
  NOR3X4 U48 ( .A(n8), .B(n9), .C(n10), .Y(n125) );
  OAI221XL U49 ( .A0(n75), .A1(n147), .B0(n146), .B1(n74), .C0(n145), .Y(
        ALUout[1]) );
  INVX6 U50 ( .A(n83), .Y(n82) );
  CLKBUFX6 U51 ( .A(n512), .Y(n74) );
  CLKINVX3 U52 ( .A(n87), .Y(n86) );
  INVXL U53 ( .A(ALUinA[0]), .Y(n126) );
  BUFX4 U54 ( .A(ALUinB[26]), .Y(n4) );
  CLKINVX1 U55 ( .A(n132), .Y(n499) );
  INVX4 U56 ( .A(n91), .Y(n90) );
  CLKINVX1 U57 ( .A(n133), .Y(n504) );
  AND4X1 U58 ( .A(n442), .B(funct_regD[5]), .C(funct_regD[0]), .D(
        funct_regD[1]), .Y(n3) );
  CLKINVX1 U59 ( .A(n96), .Y(n498) );
  CLKINVX1 U60 ( .A(n112), .Y(n80) );
  AND2X2 U61 ( .A(n426), .B(n72), .Y(n10) );
  XOR2X1 U62 ( .A(n81), .B(ALUinA[0]), .Y(n426) );
  OAI221X1 U63 ( .A0(n76), .A1(n462), .B0(n461), .B1(n74), .C0(n460), .Y(
        ALUout[27]) );
  OAI221X1 U64 ( .A0(n76), .A1(n514), .B0(n513), .B1(n74), .C0(n511), .Y(
        ALUout[31]) );
  OAI221X1 U65 ( .A0(n76), .A1(n495), .B0(n494), .B1(n74), .C0(n493), .Y(
        ALUout[30]) );
  INVX3 U66 ( .A(n38), .Y(n76) );
  CLKBUFX2 U67 ( .A(ALUinB[26]), .Y(n5) );
  AO22X4 U68 ( .A0(N408), .A1(n501), .B0(n66), .B1(N280), .Y(n506) );
  NOR4X4 U69 ( .A(n274), .B(n273), .C(n272), .D(n271), .Y(n278) );
  AO22X4 U70 ( .A0(N404), .A1(n501), .B0(N276), .B1(n66), .Y(n456) );
  BUFX4 U71 ( .A(ALUinB[7]), .Y(n41) );
  OAI31X2 U72 ( .A0(n519), .A1(ALUOp_regD[5]), .A2(ALUOp_regD[0]), .B0(n560), 
        .Y(n430) );
  OAI221X2 U73 ( .A0(n75), .A1(n197), .B0(n196), .B1(n74), .C0(n195), .Y(
        ALUout[5]) );
  NOR4X2 U74 ( .A(n308), .B(n307), .C(n306), .D(n305), .Y(n314) );
  BUFX16 U75 ( .A(ALUinB[22]), .Y(n56) );
  BUFX12 U76 ( .A(ALUinB[20]), .Y(n54) );
  OAI221X2 U77 ( .A0(n76), .A1(n162), .B0(n159), .B1(n74), .C0(n158), .Y(
        ALUout[2]) );
  BUFX20 U78 ( .A(ALUinB[13]), .Y(n47) );
  BUFX6 U79 ( .A(ALUinB[11]), .Y(n45) );
  NOR4X4 U80 ( .A(n413), .B(n412), .C(n409), .D(n408), .Y(n416) );
  CLKBUFX6 U81 ( .A(ALUinB[18]), .Y(n52) );
  BUFX20 U82 ( .A(ALUinB[21]), .Y(n55) );
  NOR4X2 U83 ( .A(n480), .B(n479), .C(n478), .D(n477), .Y(n483) );
  BUFX20 U84 ( .A(ALUinB[19]), .Y(n53) );
  OAI221X1 U85 ( .A0(n75), .A1(n365), .B0(n364), .B1(n74), .C0(n363), .Y(
        ALUout[20]) );
  AO22X4 U86 ( .A0(N312), .A1(n64), .B0(N376), .B1(n498), .Y(n507) );
  BUFX16 U87 ( .A(ALUinB[14]), .Y(n48) );
  NOR4X4 U88 ( .A(n254), .B(n253), .C(n252), .D(n251), .Y(n258) );
  OR2X6 U89 ( .A(n75), .B(n353), .Y(n6) );
  NAND3X8 U90 ( .A(n6), .B(n7), .C(n349), .Y(ALUout[19]) );
  AOI211X4 U91 ( .A0(n331), .A1(n73), .B0(n348), .C0(n347), .Y(n349) );
  INVXL U92 ( .A(ALUinA[23]), .Y(n394) );
  AND2X8 U93 ( .A(n124), .B(n138), .Y(n9) );
  OAI2BB1X4 U94 ( .A0N(n81), .A1N(n432), .B0(n122), .Y(n124) );
  OAI221X2 U95 ( .A0(n127), .A1(n74), .B0(n58), .B1(n126), .C0(n125), .Y(
        ALUout[0]) );
  BUFX12 U96 ( .A(ALUinB[0]), .Y(n81) );
  BUFX12 U97 ( .A(ALUinB[15]), .Y(n49) );
  BUFX12 U98 ( .A(ALUinB[8]), .Y(n42) );
  BUFX12 U99 ( .A(ALUinB[10]), .Y(n44) );
  BUFX12 U100 ( .A(ALUinB[12]), .Y(n46) );
  INVX4 U101 ( .A(ALUinB[3]), .Y(n87) );
  INVXL U102 ( .A(N250), .Y(n147) );
  INVXL U103 ( .A(N251), .Y(n162) );
  INVX12 U104 ( .A(n89), .Y(n88) );
  INVXL U105 ( .A(N270), .Y(n377) );
  INVXL U106 ( .A(N264), .Y(n303) );
  INVXL U107 ( .A(N276), .Y(n462) );
  INVXL U108 ( .A(N278), .Y(n484) );
  INVXL U109 ( .A(N274), .Y(n435) );
  INVXL U110 ( .A(N268), .Y(n353) );
  INVXL U111 ( .A(N259), .Y(n249) );
  INVXL U112 ( .A(N255), .Y(n207) );
  INVXL U113 ( .A(N260), .Y(n259) );
  INVXL U114 ( .A(N256), .Y(n219) );
  INVXL U115 ( .A(N258), .Y(n239) );
  INVXL U116 ( .A(N280), .Y(n514) );
  INVXL U117 ( .A(ALUinA[13]), .Y(n538) );
  INVXL U118 ( .A(ALUinA[30]), .Y(n487) );
  INVXL U119 ( .A(N267), .Y(n339) );
  INVXL U120 ( .A(N272), .Y(n404) );
  INVXL U121 ( .A(N275), .Y(n451) );
  INVXL U122 ( .A(N266), .Y(n327) );
  INVXL U123 ( .A(N263), .Y(n289) );
  INVXL U124 ( .A(N257), .Y(n229) );
  INVXL U125 ( .A(N252), .Y(n175) );
  XOR2XL U126 ( .A(n47), .B(ALUinA[13]), .Y(n391) );
  XOR2XL U127 ( .A(n40), .B(ALUinA[6]), .Y(n151) );
  XNOR2XL U128 ( .A(n394), .B(ALUinB[23]), .Y(n27) );
  XOR2XL U129 ( .A(n86), .B(ALUinA[3]), .Y(n181) );
  XOR2XL U130 ( .A(n41), .B(ALUinA[7]), .Y(n141) );
  XOR2XL U131 ( .A(n55), .B(ALUinA[21]), .Y(n301) );
  XOR2XL U132 ( .A(n54), .B(ALUinA[20]), .Y(n311) );
  XNOR2XL U133 ( .A(n465), .B(ALUinB[28]), .Y(n14) );
  XOR2XL U134 ( .A(n90), .B(ALUinA[5]), .Y(n161) );
  XOR2XL U135 ( .A(n52), .B(ALUinA[18]), .Y(n341) );
  XOR2XL U136 ( .A(n50), .B(ALUinA[16]), .Y(n361) );
  XOR2XL U137 ( .A(n51), .B(ALUinA[17]), .Y(n351) );
  XOR2XL U138 ( .A(n2), .B(ALUinA[2]), .Y(n211) );
  XOR2XL U139 ( .A(n43), .B(ALUinA[9]), .Y(n117) );
  XNOR2XL U140 ( .A(n421), .B(ALUinB[25]), .Y(n32) );
  XOR2XL U141 ( .A(n48), .B(ALUinA[14]), .Y(n381) );
  XOR2XL U142 ( .A(n45), .B(ALUinA[11]), .Y(n411) );
  XOR2XL U143 ( .A(n42), .B(ALUinA[8]), .Y(n131) );
  XOR2XL U144 ( .A(n88), .B(ALUinA[4]), .Y(n171) );
  XOR2XL U145 ( .A(n53), .B(ALUinA[19]), .Y(n331) );
  XOR2XL U146 ( .A(n82), .B(ALUinA[1]), .Y(n321) );
  XOR2XL U147 ( .A(n46), .B(ALUinA[12]), .Y(n401) );
  XNOR2XL U148 ( .A(n487), .B(ALUinB[30]), .Y(n15) );
  XNOR2XL U149 ( .A(n438), .B(ALUinB[26]), .Y(n28) );
  XOR2XL U150 ( .A(n49), .B(ALUinA[15]), .Y(n371) );
  XOR2XL U151 ( .A(n44), .B(ALUinA[10]), .Y(n422) );
  XOR2XL U152 ( .A(n56), .B(ALUinA[22]), .Y(n291) );
  XNOR2XL U153 ( .A(n454), .B(ALUinB[27]), .Y(n13) );
  XNOR2XL U154 ( .A(n502), .B(ALUinB[31]), .Y(n12) );
  XNOR2XL U155 ( .A(n407), .B(ALUinB[24]), .Y(n26) );
  MX2XL U156 ( .A(n95), .B(n94), .S0(n81), .Y(n99) );
  INVXL U157 ( .A(ALUinB[23]), .Y(n392) );
  INVXL U158 ( .A(ALUinB[25]), .Y(n418) );
  INVXL U159 ( .A(n5), .Y(n436) );
  INVXL U160 ( .A(ALUinB[24]), .Y(n405) );
  INVXL U161 ( .A(ALUinB[27]), .Y(n452) );
  INVXL U162 ( .A(ALUinB[29]), .Y(n474) );
  INVXL U163 ( .A(ALUinB[31]), .Y(n496) );
  AOI2BB1XL U164 ( .A0N(n42), .A1N(ALUinA[8]), .B0(n58), .Y(n225) );
  AOI2BB1XL U165 ( .A0N(n43), .A1N(ALUinA[9]), .B0(n58), .Y(n235) );
  AOI2BB1XL U166 ( .A0N(n41), .A1N(ALUinA[7]), .B0(n58), .Y(n215) );
  AOI2BB1XL U167 ( .A0N(n44), .A1N(ALUinA[10]), .B0(n58), .Y(n245) );
  AOI2BB1XL U168 ( .A0N(n46), .A1N(ALUinA[12]), .B0(n58), .Y(n265) );
  AOI2BB1XL U169 ( .A0N(n48), .A1N(ALUinA[14]), .B0(n59), .Y(n285) );
  AOI2BB1XL U170 ( .A0N(n51), .A1N(ALUinA[17]), .B0(n59), .Y(n323) );
  AOI2BB1XL U171 ( .A0N(n47), .A1N(ALUinA[13]), .B0(n59), .Y(n275) );
  AOI2BB1XL U172 ( .A0N(n49), .A1N(ALUinA[15]), .B0(n59), .Y(n297) );
  AOI2BB1XL U173 ( .A0N(n50), .A1N(ALUinA[16]), .B0(n59), .Y(n309) );
  AOI2BB1XL U174 ( .A0N(n53), .A1N(ALUinA[19]), .B0(n59), .Y(n347) );
  AOI2BB1XL U175 ( .A0N(n54), .A1N(ALUinA[20]), .B0(n59), .Y(n359) );
  AOI2BB1XL U176 ( .A0N(n55), .A1N(ALUinA[21]), .B0(n59), .Y(n373) );
  INVXL U177 ( .A(ALUinB[28]), .Y(n463) );
  INVXL U178 ( .A(ALUinB[30]), .Y(n485) );
  INVXL U179 ( .A(n43), .Y(n547) );
  INVXL U180 ( .A(n49), .Y(n535) );
  INVXL U181 ( .A(n44), .Y(n545) );
  INVXL U182 ( .A(n47), .Y(n539) );
  INVXL U183 ( .A(n55), .Y(n523) );
  INVXL U184 ( .A(n40), .Y(n553) );
  INVXL U185 ( .A(n52), .Y(n529) );
  AND2XL U186 ( .A(ALUinB[23]), .B(ALUinA[23]), .Y(n29) );
  AND2XL U187 ( .A(ALUinB[28]), .B(ALUinA[28]), .Y(n30) );
  AND2XL U188 ( .A(ALUinB[25]), .B(ALUinA[25]), .Y(n11) );
  AND2XL U189 ( .A(ALUinB[30]), .B(ALUinA[30]), .Y(n18) );
  AND2XL U190 ( .A(n5), .B(ALUinA[26]), .Y(n24) );
  AND2XL U191 ( .A(ALUinB[27]), .B(ALUinA[27]), .Y(n31) );
  AND2XL U192 ( .A(ALUinB[31]), .B(ALUinA[31]), .Y(n16) );
  AND3XL U193 ( .A(n42), .B(n71), .C(ALUinA[8]), .Y(n226) );
  AND3XL U194 ( .A(n48), .B(n71), .C(ALUinA[14]), .Y(n286) );
  AND3XL U195 ( .A(n51), .B(n34), .C(ALUinA[17]), .Y(n324) );
  AND3XL U196 ( .A(n46), .B(n34), .C(ALUinA[12]), .Y(n266) );
  AND3XL U197 ( .A(n47), .B(n34), .C(ALUinA[13]), .Y(n276) );
  AND3XL U198 ( .A(n50), .B(n34), .C(ALUinA[16]), .Y(n312) );
  AND3XL U199 ( .A(n53), .B(n71), .C(ALUinA[19]), .Y(n348) );
  AND3XL U200 ( .A(n54), .B(n71), .C(ALUinA[20]), .Y(n362) );
  AND3XL U201 ( .A(n55), .B(n71), .C(ALUinA[21]), .Y(n374) );
  INVXL U202 ( .A(n54), .Y(n525) );
  INVXL U203 ( .A(n56), .Y(n521) );
  INVXL U204 ( .A(n42), .Y(n549) );
  INVXL U205 ( .A(n48), .Y(n537) );
  INVXL U206 ( .A(n51), .Y(n531) );
  INVXL U207 ( .A(n45), .Y(n543) );
  INVXL U208 ( .A(n41), .Y(n551) );
  INVXL U209 ( .A(n46), .Y(n541) );
  INVXL U210 ( .A(n50), .Y(n533) );
  INVXL U211 ( .A(n53), .Y(n527) );
  XNOR2XL U212 ( .A(n476), .B(ALUinB[29]), .Y(n25) );
  INVXL U213 ( .A(ALUinA[6]), .Y(n552) );
  INVXL U214 ( .A(ALUinA[3]), .Y(n556) );
  INVXL U215 ( .A(ALUinA[7]), .Y(n550) );
  INVXL U216 ( .A(ALUinA[21]), .Y(n522) );
  INVXL U217 ( .A(ALUinA[20]), .Y(n524) );
  INVXL U218 ( .A(ALUinA[5]), .Y(n554) );
  INVXL U219 ( .A(ALUinA[18]), .Y(n528) );
  INVXL U220 ( .A(ALUinA[16]), .Y(n532) );
  INVXL U221 ( .A(ALUinA[17]), .Y(n530) );
  INVXL U222 ( .A(ALUinA[9]), .Y(n546) );
  INVXL U223 ( .A(ALUinA[14]), .Y(n536) );
  INVXL U224 ( .A(ALUinA[11]), .Y(n542) );
  INVXL U225 ( .A(ALUinA[8]), .Y(n548) );
  INVXL U226 ( .A(ALUinA[4]), .Y(n555) );
  INVXL U227 ( .A(ALUinA[19]), .Y(n526) );
  INVXL U228 ( .A(ALUinA[1]), .Y(n558) );
  INVXL U229 ( .A(ALUinA[12]), .Y(n540) );
  INVXL U230 ( .A(ALUinA[10]), .Y(n544) );
  INVXL U231 ( .A(ALUinA[22]), .Y(n520) );
  AOI2BB1XL U232 ( .A0N(n45), .A1N(ALUinA[11]), .B0(n58), .Y(n255) );
  AOI2BB1XL U233 ( .A0N(n40), .A1N(ALUinA[6]), .B0(n58), .Y(n203) );
  AOI2BB1XL U234 ( .A0N(n81), .A1N(ALUinA[0]), .B0(n77), .Y(n103) );
  AOI2BB1XL U235 ( .A0N(n52), .A1N(ALUinA[18]), .B0(n59), .Y(n335) );
  AOI2BB1XL U236 ( .A0N(n56), .A1N(ALUinA[22]), .B0(n59), .Y(n385) );
  INVXL U237 ( .A(ALUinA[27]), .Y(n454) );
  INVXL U238 ( .A(ALUinA[26]), .Y(n438) );
  INVXL U239 ( .A(ALUinA[24]), .Y(n407) );
  INVXL U240 ( .A(ALUinA[29]), .Y(n476) );
  INVXL U241 ( .A(ALUinA[28]), .Y(n465) );
  INVXL U242 ( .A(ALUinA[31]), .Y(n502) );
  AND2XL U243 ( .A(ALUinB[24]), .B(ALUinA[24]), .Y(n33) );
  AND2XL U244 ( .A(ALUinB[29]), .B(ALUinA[29]), .Y(n17) );
  AND3XL U245 ( .A(n43), .B(n34), .C(ALUinA[9]), .Y(n236) );
  AND3XL U246 ( .A(n45), .B(n34), .C(ALUinA[11]), .Y(n256) );
  AND3XL U247 ( .A(n52), .B(n34), .C(ALUinA[18]), .Y(n336) );
  AND3XL U248 ( .A(n41), .B(n34), .C(ALUinA[7]), .Y(n216) );
  AND3XL U249 ( .A(n40), .B(n34), .C(ALUinA[6]), .Y(n204) );
  AND3XL U250 ( .A(n44), .B(n34), .C(ALUinA[10]), .Y(n246) );
  AND3XL U251 ( .A(n49), .B(n34), .C(ALUinA[15]), .Y(n298) );
  AND3XL U252 ( .A(n56), .B(n71), .C(ALUinA[22]), .Y(n386) );
  AND2XL U253 ( .A(n83), .B(n60), .Y(n129) );
  AND2XL U254 ( .A(n85), .B(n61), .Y(n148) );
  AND2XL U255 ( .A(n89), .B(n60), .Y(n176) );
  AND2XL U256 ( .A(n91), .B(n61), .Y(n188) );
  AOI21X1 U257 ( .A0(n444), .A1(n102), .B0(funct_regD[1]), .Y(n500) );
  BUFX4 U258 ( .A(n111), .Y(n57) );
  NOR2X1 U259 ( .A(ALUOp_regD[4]), .B(n123), .Y(n510) );
  CLKINVX1 U260 ( .A(N269), .Y(n365) );
  CLKINVX1 U261 ( .A(N279), .Y(n495) );
  CLKINVX1 U262 ( .A(N265), .Y(n315) );
  CLKINVX1 U263 ( .A(N273), .Y(n417) );
  CLKINVX1 U264 ( .A(N277), .Y(n473) );
  CLKINVX1 U265 ( .A(N271), .Y(n389) );
  CLKINVX1 U266 ( .A(N253), .Y(n187) );
  CLKINVX1 U267 ( .A(N262), .Y(n279) );
  CLKINVX1 U268 ( .A(N254), .Y(n197) );
  CLKINVX1 U269 ( .A(N261), .Y(n269) );
  INVX3 U270 ( .A(n35), .Y(n58) );
  INVX3 U271 ( .A(n35), .Y(n59) );
  NOR4X1 U272 ( .A(n469), .B(n468), .C(n467), .D(n466), .Y(n472) );
  CLKMX2X2 U273 ( .A(n80), .B(n60), .S0(n464), .Y(n469) );
  AO22X1 U274 ( .A0(n69), .A1(n14), .B0(n30), .B1(n503), .Y(n466) );
  AO22X1 U275 ( .A0(N309), .A1(n64), .B0(N373), .B1(n63), .Y(n468) );
  CLKMX2X2 U276 ( .A(n79), .B(n60), .S0(n437), .Y(n446) );
  AO22X1 U277 ( .A0(n69), .A1(n28), .B0(n24), .B1(n503), .Y(n439) );
  AO22X1 U278 ( .A0(N307), .A1(n64), .B0(N371), .B1(n63), .Y(n443) );
  NOR4X1 U279 ( .A(n154), .B(n153), .C(n152), .D(n149), .Y(n159) );
  CLKMX2X2 U280 ( .A(n78), .B(n148), .S0(n557), .Y(n154) );
  AO22X1 U281 ( .A0(n210), .A1(n2), .B0(N283), .B1(n65), .Y(n153) );
  AO22X1 U282 ( .A0(N347), .A1(n62), .B0(n211), .B1(n69), .Y(n152) );
  NOR4X1 U283 ( .A(n167), .B(n166), .C(n165), .D(n164), .Y(n174) );
  CLKMX2X2 U284 ( .A(n78), .B(n163), .S0(n556), .Y(n167) );
  AO22X1 U285 ( .A0(n180), .A1(n86), .B0(N284), .B1(n499), .Y(n166) );
  AO22X1 U286 ( .A0(N348), .A1(n62), .B0(n181), .B1(n70), .Y(n165) );
  NOR4X1 U287 ( .A(n398), .B(n397), .C(n396), .D(n395), .Y(n403) );
  CLKMX2X2 U288 ( .A(n78), .B(n60), .S0(n393), .Y(n398) );
  AO22X1 U289 ( .A0(n69), .A1(n27), .B0(n29), .B1(n503), .Y(n395) );
  AO22X1 U290 ( .A0(N304), .A1(n64), .B0(N368), .B1(n63), .Y(n397) );
  NOR4X1 U291 ( .A(n137), .B(n136), .C(n135), .D(n134), .Y(n146) );
  CLKMX2X2 U292 ( .A(n78), .B(n129), .S0(n558), .Y(n137) );
  AO22X1 U293 ( .A0(n320), .A1(n82), .B0(N282), .B1(n64), .Y(n136) );
  AO22X1 U294 ( .A0(N346), .A1(n62), .B0(n321), .B1(n69), .Y(n135) );
  NOR4X1 U295 ( .A(n182), .B(n179), .C(n178), .D(n177), .Y(n186) );
  CLKMX2X2 U296 ( .A(n78), .B(n176), .S0(n555), .Y(n182) );
  AO22X1 U297 ( .A0(n170), .A1(n88), .B0(N285), .B1(n499), .Y(n179) );
  AO22X1 U298 ( .A0(N349), .A1(n62), .B0(n171), .B1(n504), .Y(n178) );
  NOR4X1 U299 ( .A(n192), .B(n191), .C(n190), .D(n189), .Y(n196) );
  CLKMX2X2 U300 ( .A(n78), .B(n188), .S0(n554), .Y(n192) );
  AO22X1 U301 ( .A0(n160), .A1(n90), .B0(N286), .B1(n499), .Y(n191) );
  AO22X1 U302 ( .A0(N350), .A1(n62), .B0(n161), .B1(n504), .Y(n190) );
  CLKMX2X2 U303 ( .A(n80), .B(n60), .S0(n406), .Y(n413) );
  AO22X1 U304 ( .A0(n69), .A1(n26), .B0(n33), .B1(n503), .Y(n408) );
  AO22X1 U305 ( .A0(N305), .A1(n64), .B0(N369), .B1(n63), .Y(n412) );
  NOR4X1 U306 ( .A(n428), .B(n425), .C(n424), .D(n423), .Y(n434) );
  CLKMX2X2 U307 ( .A(n79), .B(n60), .S0(n419), .Y(n428) );
  AO22X1 U308 ( .A0(n69), .A1(n32), .B0(n11), .B1(n503), .Y(n423) );
  AO22X1 U309 ( .A0(N306), .A1(n64), .B0(N370), .B1(n63), .Y(n425) );
  CLKMX2X2 U310 ( .A(n78), .B(n60), .S0(n453), .Y(n458) );
  AO22X1 U311 ( .A0(n69), .A1(n13), .B0(n31), .B1(n503), .Y(n455) );
  AO22X1 U312 ( .A0(N308), .A1(n64), .B0(N372), .B1(n63), .Y(n457) );
  CLKMX2X2 U313 ( .A(n78), .B(n60), .S0(n475), .Y(n480) );
  AO22X1 U314 ( .A0(n69), .A1(n25), .B0(n17), .B1(n503), .Y(n477) );
  AO22X1 U315 ( .A0(N310), .A1(n64), .B0(N374), .B1(n63), .Y(n479) );
  CLKMX2X2 U316 ( .A(n79), .B(n60), .S0(n486), .Y(n491) );
  AO22X1 U317 ( .A0(n69), .A1(n15), .B0(n18), .B1(n503), .Y(n488) );
  CLKMX2X2 U318 ( .A(n79), .B(n60), .S0(n497), .Y(n508) );
  AO22X1 U319 ( .A0(n69), .A1(n12), .B0(n16), .B1(n503), .Y(n505) );
  AO22X1 U320 ( .A0(N389), .A1(n68), .B0(N261), .B1(n67), .Y(n261) );
  AO22X1 U321 ( .A0(N397), .A1(n68), .B0(N269), .B1(n66), .Y(n355) );
  AO22X1 U322 ( .A0(N399), .A1(n68), .B0(N271), .B1(n66), .Y(n379) );
  AO22X1 U323 ( .A0(N394), .A1(n68), .B0(N266), .B1(n67), .Y(n317) );
  AO22X1 U324 ( .A0(N395), .A1(n68), .B0(N267), .B1(n67), .Y(n329) );
  AO22X1 U325 ( .A0(N393), .A1(n68), .B0(N265), .B1(n67), .Y(n305) );
  AO22X1 U326 ( .A0(N396), .A1(n68), .B0(N268), .B1(n66), .Y(n343) );
  AO22X1 U327 ( .A0(N398), .A1(n68), .B0(N270), .B1(n66), .Y(n367) );
  AO22X1 U328 ( .A0(N385), .A1(n501), .B0(N257), .B1(n67), .Y(n221) );
  AO22X1 U329 ( .A0(N391), .A1(n68), .B0(N263), .B1(n67), .Y(n281) );
  AO22X1 U330 ( .A0(N386), .A1(n501), .B0(N258), .B1(n67), .Y(n231) );
  AO22X1 U331 ( .A0(N388), .A1(n501), .B0(N260), .B1(n67), .Y(n251) );
  AO22X1 U332 ( .A0(N379), .A1(n501), .B0(N251), .B1(n67), .Y(n149) );
  AO22X1 U333 ( .A0(N380), .A1(n501), .B0(N252), .B1(n500), .Y(n164) );
  AO22X1 U334 ( .A0(N378), .A1(n501), .B0(N250), .B1(n66), .Y(n134) );
  AO22X1 U335 ( .A0(N382), .A1(n501), .B0(N254), .B1(n66), .Y(n189) );
  AO22X1 U336 ( .A0(N387), .A1(n501), .B0(N259), .B1(n67), .Y(n241) );
  AO22X1 U337 ( .A0(N390), .A1(n68), .B0(N262), .B1(n67), .Y(n271) );
  AO22X1 U338 ( .A0(N392), .A1(n68), .B0(N264), .B1(n67), .Y(n293) );
  AO22X1 U339 ( .A0(N384), .A1(n501), .B0(N256), .B1(n67), .Y(n209) );
  AO22X1 U340 ( .A0(N381), .A1(n501), .B0(N253), .B1(n67), .Y(n177) );
  AO22X1 U341 ( .A0(N383), .A1(n501), .B0(N255), .B1(n67), .Y(n199) );
  AO22X1 U342 ( .A0(N400), .A1(n68), .B0(N272), .B1(n66), .Y(n396) );
  AO22X1 U343 ( .A0(N405), .A1(n501), .B0(N277), .B1(n66), .Y(n467) );
  AO22X1 U344 ( .A0(N403), .A1(n501), .B0(N275), .B1(n66), .Y(n440) );
  AO22X1 U345 ( .A0(N401), .A1(n68), .B0(N273), .B1(n66), .Y(n409) );
  AO22X1 U346 ( .A0(N402), .A1(n501), .B0(N274), .B1(n66), .Y(n424) );
  AO22X1 U347 ( .A0(N406), .A1(n68), .B0(N278), .B1(n66), .Y(n478) );
  AO22X1 U348 ( .A0(N407), .A1(n501), .B0(N279), .B1(n66), .Y(n489) );
  AO22X1 U349 ( .A0(N377), .A1(n501), .B0(N249), .B1(n66), .Y(n105) );
  CLKINVX1 U350 ( .A(n431), .Y(n419) );
  CLKINVX1 U351 ( .A(n426), .Y(n97) );
  CLKINVX1 U352 ( .A(n459), .Y(n453) );
  CLKINVX1 U353 ( .A(n509), .Y(n497) );
  CLKINVX1 U354 ( .A(n414), .Y(n406) );
  CLKINVX1 U355 ( .A(n481), .Y(n475) );
  CLKINVX1 U356 ( .A(n399), .Y(n393) );
  CLKINVX1 U357 ( .A(n470), .Y(n464) );
  CLKINVX1 U358 ( .A(n448), .Y(n437) );
  CLKINVX1 U359 ( .A(n492), .Y(n486) );
  AOI2BB1X1 U360 ( .A0N(n82), .A1N(n142), .B0(n58), .Y(n143) );
  AOI2BB1X1 U361 ( .A0N(n88), .A1N(ALUinA[4]), .B0(n58), .Y(n183) );
  AOI2BB1X1 U362 ( .A0N(n90), .A1N(ALUinA[5]), .B0(n58), .Y(n193) );
  AOI2BB1X1 U363 ( .A0N(n2), .A1N(n155), .B0(n58), .Y(n156) );
  AOI2BB1X1 U364 ( .A0N(n86), .A1N(n168), .B0(n58), .Y(n169) );
  NAND2X1 U365 ( .A(n60), .B(n126), .Y(n95) );
  CLKINVX1 U366 ( .A(n558), .Y(n142) );
  CLKINVX1 U367 ( .A(n556), .Y(n168) );
  CLKINVX1 U368 ( .A(n557), .Y(n155) );
  NAND2X1 U369 ( .A(ALUinA[0]), .B(n503), .Y(n94) );
  CLKBUFX3 U370 ( .A(n499), .Y(n64) );
  CLKBUFX3 U371 ( .A(n499), .Y(n65) );
  AND3X2 U372 ( .A(n82), .B(n71), .C(n142), .Y(n144) );
  AND3X2 U373 ( .A(n88), .B(n71), .C(ALUinA[4]), .Y(n184) );
  AND3X2 U374 ( .A(n90), .B(n71), .C(ALUinA[5]), .Y(n194) );
  AND3X2 U375 ( .A(n2), .B(n34), .C(n155), .Y(n157) );
  AND3X2 U376 ( .A(n86), .B(n34), .C(n168), .Y(n172) );
  CLKBUFX3 U377 ( .A(n34), .Y(n71) );
  INVX3 U378 ( .A(n79), .Y(n77) );
  CLKBUFX3 U379 ( .A(n504), .Y(n69) );
  CLKBUFX3 U380 ( .A(n504), .Y(n70) );
  NOR4X1 U381 ( .A(n224), .B(n223), .C(n222), .D(n221), .Y(n228) );
  CLKMX2X2 U382 ( .A(n78), .B(n220), .S0(n548), .Y(n224) );
  AO22X1 U383 ( .A0(n130), .A1(n42), .B0(N289), .B1(n65), .Y(n223) );
  AO22X1 U384 ( .A0(N353), .A1(n62), .B0(n131), .B1(n70), .Y(n222) );
  NOR4X1 U385 ( .A(n284), .B(n283), .C(n282), .D(n281), .Y(n288) );
  CLKMX2X2 U386 ( .A(n79), .B(n280), .S0(n536), .Y(n284) );
  AO22X1 U387 ( .A0(n380), .A1(n48), .B0(N295), .B1(n65), .Y(n283) );
  AO22X1 U388 ( .A0(N359), .A1(n63), .B0(n381), .B1(n70), .Y(n282) );
  NOR4X1 U389 ( .A(n234), .B(n233), .C(n232), .D(n231), .Y(n238) );
  CLKMX2X2 U390 ( .A(n79), .B(n230), .S0(n546), .Y(n234) );
  AO22X1 U391 ( .A0(n110), .A1(n43), .B0(N290), .B1(n65), .Y(n233) );
  AO22X1 U392 ( .A0(N354), .A1(n62), .B0(n117), .B1(n70), .Y(n232) );
  NOR4X1 U393 ( .A(n322), .B(n319), .C(n318), .D(n317), .Y(n326) );
  CLKMX2X2 U394 ( .A(n79), .B(n316), .S0(n530), .Y(n322) );
  AO22X1 U395 ( .A0(N362), .A1(n63), .B0(n351), .B1(n70), .Y(n318) );
  AO22X1 U396 ( .A0(n350), .A1(n51), .B0(N298), .B1(n65), .Y(n319) );
  CLKMX2X2 U397 ( .A(n79), .B(n250), .S0(n542), .Y(n254) );
  AO22X1 U398 ( .A0(n410), .A1(n45), .B0(N292), .B1(n65), .Y(n253) );
  AO22X1 U399 ( .A0(N356), .A1(n62), .B0(n411), .B1(n70), .Y(n252) );
  CLKMX2X2 U400 ( .A(n80), .B(n328), .S0(n528), .Y(n334) );
  AO22X1 U401 ( .A0(N363), .A1(n63), .B0(n341), .B1(n70), .Y(n332) );
  AO22X1 U402 ( .A0(n340), .A1(n52), .B0(N299), .B1(n65), .Y(n333) );
  NOR4X1 U403 ( .A(n214), .B(n213), .C(n212), .D(n209), .Y(n218) );
  CLKMX2X2 U404 ( .A(n78), .B(n208), .S0(n550), .Y(n214) );
  AO22X1 U405 ( .A0(n140), .A1(n41), .B0(N288), .B1(n65), .Y(n213) );
  AO22X1 U406 ( .A0(N352), .A1(n62), .B0(n141), .B1(n70), .Y(n212) );
  NOR4X1 U407 ( .A(n202), .B(n201), .C(n200), .D(n199), .Y(n206) );
  CLKMX2X2 U408 ( .A(n78), .B(n198), .S0(n552), .Y(n202) );
  AO22X1 U409 ( .A0(n150), .A1(n40), .B0(N287), .B1(n65), .Y(n201) );
  AO22X1 U410 ( .A0(N351), .A1(n62), .B0(n151), .B1(n70), .Y(n200) );
  NOR4X1 U411 ( .A(n244), .B(n243), .C(n242), .D(n241), .Y(n248) );
  CLKMX2X2 U412 ( .A(n79), .B(n240), .S0(n544), .Y(n244) );
  AO22X1 U413 ( .A0(n420), .A1(n44), .B0(N291), .B1(n65), .Y(n243) );
  AO22X1 U414 ( .A0(N355), .A1(n62), .B0(n422), .B1(n70), .Y(n242) );
  NOR4X1 U415 ( .A(n264), .B(n263), .C(n262), .D(n261), .Y(n268) );
  CLKMX2X2 U416 ( .A(n79), .B(n260), .S0(n540), .Y(n264) );
  AO22X1 U417 ( .A0(n400), .A1(n46), .B0(N293), .B1(n65), .Y(n263) );
  AO22X1 U418 ( .A0(N357), .A1(n62), .B0(n401), .B1(n70), .Y(n262) );
  CLKMX2X2 U419 ( .A(n79), .B(n270), .S0(n538), .Y(n274) );
  AO22X1 U420 ( .A0(n390), .A1(n47), .B0(N294), .B1(n65), .Y(n273) );
  AO22X1 U421 ( .A0(N358), .A1(n62), .B0(n391), .B1(n70), .Y(n272) );
  NOR4X1 U422 ( .A(n296), .B(n295), .C(n294), .D(n293), .Y(n302) );
  CLKMX2X2 U423 ( .A(n80), .B(n292), .S0(n534), .Y(n296) );
  AO22X1 U424 ( .A0(n370), .A1(n49), .B0(N296), .B1(n65), .Y(n295) );
  AO22X1 U425 ( .A0(N360), .A1(n63), .B0(n371), .B1(n70), .Y(n294) );
  CLKMX2X2 U426 ( .A(n79), .B(n304), .S0(n532), .Y(n308) );
  AO22X1 U427 ( .A0(n360), .A1(n50), .B0(N297), .B1(n65), .Y(n307) );
  CLKMX2X2 U428 ( .A(n78), .B(n342), .S0(n526), .Y(n346) );
  AO22X1 U429 ( .A0(N364), .A1(n63), .B0(n331), .B1(n69), .Y(n344) );
  NOR4X1 U430 ( .A(n358), .B(n357), .C(n356), .D(n355), .Y(n364) );
  CLKMX2X2 U431 ( .A(n78), .B(n354), .S0(n524), .Y(n358) );
  AO22X1 U432 ( .A0(N365), .A1(n63), .B0(n311), .B1(n69), .Y(n356) );
  AO22X1 U433 ( .A0(n310), .A1(n54), .B0(N301), .B1(n64), .Y(n357) );
  CLKMX2X2 U434 ( .A(n78), .B(n366), .S0(n522), .Y(n372) );
  AO22X1 U435 ( .A0(N366), .A1(n63), .B0(n301), .B1(n69), .Y(n368) );
  AO22X1 U436 ( .A0(n300), .A1(n55), .B0(N302), .B1(n64), .Y(n369) );
  NOR4X1 U437 ( .A(n384), .B(n383), .C(n382), .D(n379), .Y(n388) );
  CLKMX2X2 U438 ( .A(n79), .B(n378), .S0(n520), .Y(n384) );
  AO22X1 U439 ( .A0(N367), .A1(n63), .B0(n291), .B1(n69), .Y(n382) );
  AO22X1 U440 ( .A0(n290), .A1(n56), .B0(N303), .B1(n64), .Y(n383) );
  OAI211X1 U441 ( .A0(n132), .A1(n100), .B0(n99), .C0(n98), .Y(n106) );
  CLKINVX1 U442 ( .A(N281), .Y(n100) );
  AOI2BB2X1 U443 ( .B0(N345), .B1(n62), .A0N(n133), .A1N(n97), .Y(n98) );
  AOI222XL U444 ( .A0(n72), .A1(n27), .B0(n29), .B1(n71), .C0(n35), .C1(n399), 
        .Y(n402) );
  AOI222XL U445 ( .A0(n72), .A1(n28), .B0(n24), .B1(n71), .C0(n35), .C1(n448), 
        .Y(n449) );
  AOI211X1 U446 ( .A0(n341), .A1(n73), .B0(n336), .C0(n335), .Y(n337) );
  OAI221XL U447 ( .A0(n75), .A1(n327), .B0(n326), .B1(n74), .C0(n325), .Y(
        ALUout[17]) );
  AOI211X1 U448 ( .A0(n351), .A1(n73), .B0(n324), .C0(n323), .Y(n325) );
  AOI211X1 U449 ( .A0(n131), .A1(n73), .B0(n226), .C0(n225), .Y(n227) );
  AOI211X1 U450 ( .A0(n381), .A1(n73), .B0(n286), .C0(n285), .Y(n287) );
  AOI211X1 U451 ( .A0(n181), .A1(n73), .B0(n172), .C0(n169), .Y(n173) );
  NAND2X1 U452 ( .A(n454), .B(n452), .Y(n459) );
  NAND2X1 U453 ( .A(n476), .B(n474), .Y(n481) );
  NAND2X1 U454 ( .A(n407), .B(n405), .Y(n414) );
  NAND2X1 U455 ( .A(n394), .B(n392), .Y(n399) );
  NAND2X1 U456 ( .A(n465), .B(n463), .Y(n470) );
  NAND2X1 U457 ( .A(n438), .B(n436), .Y(n448) );
  NAND2X1 U458 ( .A(n487), .B(n485), .Y(n492) );
  NAND2X1 U459 ( .A(n502), .B(n496), .Y(n509) );
  CLKINVX1 U460 ( .A(ALUinA[2]), .Y(n557) );
  CLKINVX1 U461 ( .A(ALUinA[15]), .Y(n534) );
  OAI21XL U462 ( .A0(n57), .A1(n536), .B0(n112), .Y(n380) );
  OAI21XL U463 ( .A0(n57), .A1(n538), .B0(n112), .Y(n390) );
  OAI21XL U464 ( .A0(n57), .A1(n524), .B0(n77), .Y(n310) );
  OAI21XL U465 ( .A0(n57), .A1(n530), .B0(n77), .Y(n350) );
  OAI21XL U466 ( .A0(n57), .A1(n528), .B0(n112), .Y(n340) );
  OAI21XL U467 ( .A0(n57), .A1(n542), .B0(n112), .Y(n410) );
  OAI21XL U468 ( .A0(n57), .A1(n558), .B0(n77), .Y(n320) );
  OAI21XL U469 ( .A0(n57), .A1(n552), .B0(n77), .Y(n150) );
  OAI21XL U470 ( .A0(n57), .A1(n554), .B0(n77), .Y(n160) );
  OAI21XL U471 ( .A0(n57), .A1(n555), .B0(n77), .Y(n170) );
  OAI21XL U472 ( .A0(n57), .A1(n540), .B0(n77), .Y(n400) );
  OAI21XL U473 ( .A0(n57), .A1(n522), .B0(n77), .Y(n300) );
  OAI21XL U474 ( .A0(n57), .A1(n548), .B0(n77), .Y(n130) );
  OAI21XL U475 ( .A0(n57), .A1(n557), .B0(n77), .Y(n210) );
  OAI21XL U476 ( .A0(n57), .A1(n556), .B0(n77), .Y(n180) );
  OAI21XL U477 ( .A0(n57), .A1(n550), .B0(n77), .Y(n140) );
  OAI21XL U478 ( .A0(n57), .A1(n544), .B0(n77), .Y(n420) );
  OAI21XL U479 ( .A0(n57), .A1(n534), .B0(n112), .Y(n370) );
  OAI21XL U480 ( .A0(n57), .A1(n532), .B0(n112), .Y(n360) );
  OAI21XL U481 ( .A0(n57), .A1(n526), .B0(n77), .Y(n330) );
  OAI21XL U482 ( .A0(n57), .A1(n520), .B0(n77), .Y(n290) );
  OAI21XL U483 ( .A0(n546), .A1(n57), .B0(n77), .Y(n110) );
  CLKBUFX3 U484 ( .A(n498), .Y(n63) );
  CLKBUFX3 U485 ( .A(n498), .Y(n62) );
  CLKBUFX3 U486 ( .A(n500), .Y(n66) );
  CLKBUFX3 U487 ( .A(n500), .Y(n67) );
  AND2X2 U488 ( .A(n541), .B(n61), .Y(n260) );
  AND2X2 U489 ( .A(n553), .B(n61), .Y(n198) );
  AND2X2 U490 ( .A(n527), .B(n61), .Y(n342) );
  AND2X2 U491 ( .A(n551), .B(n61), .Y(n208) );
  AND2X2 U492 ( .A(n535), .B(n61), .Y(n292) );
  AND2X2 U493 ( .A(n549), .B(n61), .Y(n220) );
  AND2X2 U494 ( .A(n543), .B(n61), .Y(n250) );
  AND2X2 U495 ( .A(n533), .B(n61), .Y(n304) );
  AND2X2 U496 ( .A(n531), .B(n61), .Y(n316) );
  AND2X2 U497 ( .A(n521), .B(n60), .Y(n378) );
  AND2X2 U498 ( .A(n537), .B(n61), .Y(n280) );
  AND2X2 U499 ( .A(n525), .B(n60), .Y(n354) );
  AND2X2 U500 ( .A(n87), .B(n61), .Y(n163) );
  AND2X2 U501 ( .A(n523), .B(n60), .Y(n366) );
  AND2X2 U502 ( .A(n547), .B(n61), .Y(n230) );
  AND2X2 U503 ( .A(n545), .B(n61), .Y(n240) );
  AND2X2 U504 ( .A(n539), .B(n61), .Y(n270) );
  AND2X2 U505 ( .A(n529), .B(n61), .Y(n328) );
  AND2X2 U506 ( .A(n139), .B(n138), .Y(n34) );
  CLKINVX1 U507 ( .A(n560), .Y(n116) );
  NAND2X1 U508 ( .A(n128), .B(n109), .Y(n114) );
  CLKINVX1 U509 ( .A(n429), .Y(n109) );
  CLKBUFX3 U510 ( .A(n80), .Y(n78) );
  CLKBUFX3 U511 ( .A(n80), .Y(n79) );
  AND2X2 U512 ( .A(n108), .B(n138), .Y(n35) );
  CLKBUFX3 U513 ( .A(n510), .Y(n72) );
  CLKBUFX3 U514 ( .A(n510), .Y(n73) );
  CLKBUFX3 U515 ( .A(n3), .Y(n60) );
  CLKBUFX3 U516 ( .A(n3), .Y(n61) );
  CLKBUFX3 U517 ( .A(n501), .Y(n68) );
  INVX3 U518 ( .A(n57), .Y(n503) );
  INVX3 U519 ( .A(n38), .Y(n75) );
  NOR4X1 U520 ( .A(n441), .B(n559), .C(funct_regD[0]), .D(funct_regD[2]), .Y(
        n104) );
  AOI32X1 U521 ( .A0(funct_regD[5]), .A1(funct_regD[1]), .A2(N441), .B0(n518), 
        .B1(n516), .Y(n441) );
  OAI21XL U522 ( .A0(n119), .A1(n126), .B0(n120), .Y(n432) );
  CLKMX2X2 U523 ( .A(n121), .B(n118), .S0(ALUOp_regD[1]), .Y(n122) );
  NOR4X1 U524 ( .A(n106), .B(n105), .C(n104), .D(n103), .Y(n127) );
  AOI211X1 U525 ( .A0(n361), .A1(n73), .B0(n312), .C0(n309), .Y(n313) );
  AOI211X1 U526 ( .A0(n311), .A1(n73), .B0(n362), .C0(n359), .Y(n363) );
  AOI211X1 U527 ( .A0(n301), .A1(n72), .B0(n374), .C0(n373), .Y(n375) );
  AOI211X1 U528 ( .A0(n291), .A1(n72), .B0(n386), .C0(n385), .Y(n387) );
  NAND2X1 U529 ( .A(n115), .B(n430), .Y(n118) );
  AOI211X1 U530 ( .A0(n161), .A1(n73), .B0(n194), .C0(n193), .Y(n195) );
  OAI221XL U531 ( .A0(n76), .A1(n207), .B0(n206), .B1(n74), .C0(n205), .Y(
        ALUout[6]) );
  AOI211X1 U532 ( .A0(n151), .A1(n73), .B0(n204), .C0(n203), .Y(n205) );
  OAI221XL U533 ( .A0(n76), .A1(n249), .B0(n248), .B1(n74), .C0(n247), .Y(
        ALUout[10]) );
  AOI211X1 U534 ( .A0(n422), .A1(n73), .B0(n246), .C0(n245), .Y(n247) );
  OAI221XL U535 ( .A0(n76), .A1(n269), .B0(n268), .B1(n74), .C0(n267), .Y(
        ALUout[12]) );
  AOI211X1 U536 ( .A0(n401), .A1(n73), .B0(n266), .C0(n265), .Y(n267) );
  AOI211X1 U537 ( .A0(n391), .A1(n73), .B0(n276), .C0(n275), .Y(n277) );
  AOI211X1 U538 ( .A0(n371), .A1(n73), .B0(n298), .C0(n297), .Y(n299) );
  AOI222XL U539 ( .A0(n72), .A1(n26), .B0(n33), .B1(n71), .C0(n35), .C1(n414), 
        .Y(n415) );
  OAI221XL U540 ( .A0(n76), .A1(n435), .B0(n434), .B1(n74), .C0(n433), .Y(
        ALUout[25]) );
  AOI222XL U541 ( .A0(n72), .A1(n32), .B0(n11), .B1(n71), .C0(n35), .C1(n431), 
        .Y(n433) );
  AOI222XL U542 ( .A0(n72), .A1(n13), .B0(n31), .B1(n71), .C0(n35), .C1(n459), 
        .Y(n460) );
  AOI222XL U543 ( .A0(n72), .A1(n25), .B0(n17), .B1(n71), .C0(n35), .C1(n481), 
        .Y(n482) );
  AOI222XL U544 ( .A0(n72), .A1(n15), .B0(n18), .B1(n71), .C0(n35), .C1(n492), 
        .Y(n493) );
  AOI222XL U545 ( .A0(n72), .A1(n12), .B0(n16), .B1(n71), .C0(n35), .C1(n509), 
        .Y(n511) );
  AOI211X1 U546 ( .A0(n321), .A1(n72), .B0(n144), .C0(n143), .Y(n145) );
  AOI211X1 U547 ( .A0(n171), .A1(n73), .B0(n184), .C0(n183), .Y(n185) );
  CLKBUFX3 U548 ( .A(ALUinB[17]), .Y(n51) );
  AOI222XL U549 ( .A0(n72), .A1(n14), .B0(n30), .B1(n71), .C0(n35), .C1(n470), 
        .Y(n471) );
  OAI221XL U550 ( .A0(n76), .A1(n239), .B0(n238), .B1(n74), .C0(n237), .Y(
        ALUout[9]) );
  AOI211X1 U551 ( .A0(n117), .A1(n73), .B0(n236), .C0(n235), .Y(n237) );
  AOI211X1 U552 ( .A0(n411), .A1(n73), .B0(n256), .C0(n255), .Y(n257) );
  AOI211X1 U553 ( .A0(n141), .A1(n73), .B0(n216), .C0(n215), .Y(n217) );
  AOI211X1 U554 ( .A0(n211), .A1(n73), .B0(n157), .C0(n156), .Y(n158) );
  INVX3 U555 ( .A(ALUinB[2]), .Y(n85) );
  INVX3 U556 ( .A(ALUinB[1]), .Y(n83) );
  INVX3 U557 ( .A(ALUinB[4]), .Y(n89) );
  INVX3 U558 ( .A(ALUinB[5]), .Y(n91) );
  NAND4X1 U559 ( .A(funct_regD[3]), .B(funct_regD[0]), .C(n517), .D(n516), .Y(
        n444) );
  NAND2X1 U560 ( .A(n36), .B(funct_regD[5]), .Y(n102) );
  NAND3BX1 U561 ( .AN(funct_regD[1]), .B(n516), .C(n36), .Y(n96) );
  NAND3BX1 U562 ( .AN(n516), .B(funct_regD[1]), .C(n36), .Y(n132) );
  CLKINVX1 U563 ( .A(funct_regD[2]), .Y(n517) );
  NOR2BX1 U564 ( .AN(n37), .B(funct_regD[0]), .Y(n36) );
  NOR2BX1 U565 ( .AN(n517), .B(funct_regD[3]), .Y(n37) );
  NOR2X1 U566 ( .A(funct_regD[3]), .B(n517), .Y(n442) );
  NAND3BX1 U567 ( .AN(funct_regD[5]), .B(funct_regD[1]), .C(n37), .Y(n101) );
  NAND4X1 U568 ( .A(ALUOp_regD[2]), .B(ALUOp_regD[3]), .C(n515), .D(n128), .Y(
        n119) );
  NAND4X1 U569 ( .A(ALUOp_regD[3]), .B(ALUOp_regD[2]), .C(n427), .D(
        ALUOp_regD[1]), .Y(n123) );
  NOR2X1 U570 ( .A(ALUOp_regD[5]), .B(ALUOp_regD[0]), .Y(n427) );
  NAND4X1 U571 ( .A(n447), .B(ALUOp_regD[3]), .C(ALUOp_regD[0]), .D(
        ALUOp_regD[2]), .Y(n120) );
  NOR2X1 U572 ( .A(ALUOp_regD[5]), .B(ALUOp_regD[1]), .Y(n447) );
  CLKINVX1 U573 ( .A(funct_regD[5]), .Y(n516) );
  CLKINVX1 U574 ( .A(funct_regD[1]), .Y(n518) );
  NAND4X1 U575 ( .A(n445), .B(funct_regD[5]), .C(funct_regD[2]), .D(
        funct_regD[1]), .Y(n133) );
  NOR2X1 U576 ( .A(funct_regD[3]), .B(funct_regD[0]), .Y(n445) );
  NAND3BX1 U577 ( .AN(ALUOp_regD[3]), .B(n515), .C(n92), .Y(n560) );
  CLKINVX1 U578 ( .A(ALUOp_regD[0]), .Y(n92) );
  CLKINVX1 U579 ( .A(ALUOp_regD[5]), .Y(n515) );
  CLKINVX1 U580 ( .A(ALUOp_regD[1]), .Y(n128) );
  NAND4X1 U581 ( .A(funct_regD[5]), .B(funct_regD[2]), .C(n518), .D(n559), .Y(
        n111) );
  CLKINVX1 U582 ( .A(ALUOp_regD[2]), .Y(n115) );
  CLKINVX1 U583 ( .A(funct_regD[3]), .Y(n559) );
  NAND2X1 U584 ( .A(ALUOp_regD[3]), .B(n515), .Y(n429) );
  NAND3BX1 U585 ( .AN(funct_regD[3]), .B(n518), .C(n93), .Y(n112) );
  AND3X2 U586 ( .A(funct_regD[2]), .B(funct_regD[5]), .C(funct_regD[0]), .Y(
        n93) );
  NAND2X1 U587 ( .A(ALUOp_regD[2]), .B(n116), .Y(n121) );
  AND3X2 U588 ( .A(n39), .B(n138), .C(n115), .Y(n38) );
  MXI2X1 U589 ( .A(n114), .B(n113), .S0(ALUOp_regD[0]), .Y(n39) );
  NAND3BX1 U590 ( .AN(funct_regD[4]), .B(n115), .C(n107), .Y(n512) );
  AND3X2 U591 ( .A(n116), .B(n128), .C(n138), .Y(n107) );
  NAND2X1 U592 ( .A(n421), .B(n418), .Y(n431) );
  INVXL U593 ( .A(ALUinA[25]), .Y(n421) );
  CLKINVX3 U594 ( .A(n101), .Y(n501) );
endmodule


module MIPS_Pipeline_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n47;
  wire   [31:1] carry;

  ADDFHX4 U1_4 ( .A(A[4]), .B(1'b0), .CI(n21), .CO(carry[5]), .S(SUM[4]) );
  NAND3X2 U1 ( .A(n17), .B(1'b1), .C(1'b1), .Y(carry[6]) );
  XOR3XL U2 ( .A(carry[5]), .B(1'b0), .C(A[5]), .Y(SUM[5]) );
  AND2X4 U4 ( .A(A[15]), .B(n36), .Y(n37) );
  CLKAND2X3 U5 ( .A(A[14]), .B(n35), .Y(n36) );
  XNOR2X2 U6 ( .A(A[31]), .B(n47), .Y(SUM[31]) );
  NAND2X1 U7 ( .A(A[27]), .B(n10), .Y(n11) );
  NAND2X2 U8 ( .A(A[30]), .B(n30), .Y(n47) );
  NAND2X1 U9 ( .A(n3), .B(n30), .Y(n6) );
  CLKAND2X8 U10 ( .A(A[29]), .B(n7), .Y(n30) );
  NAND2X4 U11 ( .A(n15), .B(n16), .Y(SUM[28]) );
  NAND2X4 U12 ( .A(A[28]), .B(n14), .Y(n15) );
  AND2X1 U13 ( .A(A[27]), .B(n40), .Y(n8) );
  CLKAND2X12 U14 ( .A(A[26]), .B(n22), .Y(n40) );
  NAND2X2 U15 ( .A(n11), .B(n12), .Y(SUM[27]) );
  CLKINVX2 U16 ( .A(n30), .Y(n4) );
  NAND2X2 U17 ( .A(A[30]), .B(n4), .Y(n5) );
  CLKXOR2X1 U18 ( .A(A[21]), .B(n43), .Y(SUM[21]) );
  CLKAND2X12 U19 ( .A(A[21]), .B(n43), .Y(n27) );
  CLKAND2X12 U20 ( .A(A[20]), .B(n26), .Y(n43) );
  CLKXOR2X1 U21 ( .A(A[7]), .B(n44), .Y(SUM[7]) );
  AND2X4 U22 ( .A(A[7]), .B(n44), .Y(n23) );
  CLKAND2X2 U23 ( .A(A[6]), .B(carry[6]), .Y(n44) );
  AND2X8 U24 ( .A(A[22]), .B(n27), .Y(n28) );
  NAND2X2 U25 ( .A(n19), .B(n20), .Y(SUM[29]) );
  AND2X2 U26 ( .A(A[18]), .B(n25), .Y(n39) );
  CLKAND2X8 U27 ( .A(A[24]), .B(n29), .Y(n42) );
  CLKAND2X6 U28 ( .A(A[19]), .B(n39), .Y(n26) );
  AND2X4 U29 ( .A(A[25]), .B(n42), .Y(n22) );
  CLKAND2X8 U30 ( .A(A[27]), .B(n40), .Y(n41) );
  AND2X6 U31 ( .A(A[8]), .B(n23), .Y(n24) );
  AND2X6 U32 ( .A(A[13]), .B(n33), .Y(n35) );
  AND2X4 U33 ( .A(A[10]), .B(n31), .Y(n32) );
  NAND2X1 U34 ( .A(A[28]), .B(n41), .Y(n2) );
  XOR2X1 U35 ( .A(A[13]), .B(n33), .Y(SUM[13]) );
  AND2X2 U36 ( .A(A[12]), .B(n34), .Y(n33) );
  AND2X4 U37 ( .A(A[16]), .B(n37), .Y(n38) );
  XOR2XL U38 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  AND2X2 U39 ( .A(A[9]), .B(n24), .Y(n31) );
  NAND2X2 U40 ( .A(n5), .B(n6), .Y(SUM[30]) );
  AND2X4 U41 ( .A(A[11]), .B(n32), .Y(n34) );
  AND2X6 U42 ( .A(A[23]), .B(n28), .Y(n29) );
  XOR2X1 U43 ( .A(A[11]), .B(n32), .Y(SUM[11]) );
  AND2X2 U44 ( .A(A[28]), .B(n41), .Y(n7) );
  INVXL U45 ( .A(A[30]), .Y(n3) );
  XOR2X1 U46 ( .A(A[22]), .B(n27), .Y(SUM[22]) );
  AND2X4 U47 ( .A(A[17]), .B(n38), .Y(n25) );
  NAND2XL U48 ( .A(A[5]), .B(carry[5]), .Y(n17) );
  XOR2X1 U49 ( .A(A[24]), .B(n29), .Y(SUM[24]) );
  AND2X6 U50 ( .A(A[3]), .B(A[2]), .Y(n21) );
  XOR2X1 U51 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  NAND2X1 U52 ( .A(n9), .B(n40), .Y(n12) );
  INVXL U53 ( .A(A[27]), .Y(n9) );
  CLKINVX1 U54 ( .A(n40), .Y(n10) );
  NAND2XL U55 ( .A(A[29]), .B(n2), .Y(n19) );
  NAND2X1 U56 ( .A(n18), .B(n7), .Y(n20) );
  INVXL U57 ( .A(A[29]), .Y(n18) );
  NAND2X1 U58 ( .A(n13), .B(n8), .Y(n16) );
  CLKINVX1 U59 ( .A(n8), .Y(n14) );
  INVXL U60 ( .A(A[28]), .Y(n13) );
  INVXL U61 ( .A(A[2]), .Y(SUM[2]) );
  XOR2X1 U62 ( .A(A[26]), .B(n22), .Y(SUM[26]) );
  XOR2X1 U63 ( .A(A[25]), .B(n42), .Y(SUM[25]) );
  XOR2X1 U64 ( .A(A[23]), .B(n28), .Y(SUM[23]) );
  XOR2X1 U65 ( .A(A[20]), .B(n26), .Y(SUM[20]) );
  XOR2X1 U66 ( .A(A[10]), .B(n31), .Y(SUM[10]) );
  XOR2X1 U67 ( .A(A[19]), .B(n39), .Y(SUM[19]) );
  XOR2X1 U68 ( .A(A[18]), .B(n25), .Y(SUM[18]) );
  XOR2X1 U69 ( .A(A[17]), .B(n38), .Y(SUM[17]) );
  XOR2X1 U70 ( .A(A[16]), .B(n37), .Y(SUM[16]) );
  XOR2X1 U71 ( .A(A[15]), .B(n36), .Y(SUM[15]) );
  XOR2X1 U72 ( .A(A[14]), .B(n35), .Y(SUM[14]) );
  XOR2X1 U73 ( .A(A[12]), .B(n34), .Y(SUM[12]) );
  XOR2X1 U74 ( .A(A[9]), .B(n24), .Y(SUM[9]) );
  XOR2X1 U75 ( .A(A[8]), .B(n23), .Y(SUM[8]) );
  CLKBUFX3 U76 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U77 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, flush,
         stallcache, stall_lw_use, JumpReg_m, MemRead_m, MemWrite_m, ALUsrc,
         RegWrite_m, Branch_DEC_m, MemRead_regD, MemWrite_regD, ALUsrc_regD,
         RegWrite_regD, JumpReg_regD, Branch_regD, RegWrite_regE,
         RegWrite_regM, Branch_DEC, MemRead, MemWrite, RegWrite, JumpReg,
         ExtOp, branchpred_his, pred_cond, predict, Jump_IF, Branch_IF, N22,
         n9, n52, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n94, n96, n97, n98, n102, n103, n105, n106, n110, n111, n115,
         n117, n120, n121, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186;
  wire   [31:0] PCplus4;
  wire   [15:0] branchOffset_D;
  wire   [5:0] opcode;
  wire   [4:0] Rs;
  wire   [4:0] Rt;
  wire   [4:0] Rd;
  wire   [4:0] shamt;
  wire   [5:0] funct;
  wire   [15:0] immediate;
  wire   [31:0] PCplus4_regI;
  wire   [1:0] MemtoReg;
  wire   [5:0] ALUOp;
  wire   [31:0] A_f;
  wire   [31:0] B_f;
  wire   [31:0] ExtOut;
  wire   [4:0] wsel;
  wire   [1:0] MemtoReg_regD;
  wire   [5:0] ALUOp_regD;
  wire   [5:0] funct_regD;
  wire   [31:0] A_regD;
  wire   [31:0] B_regD;
  wire   [31:0] ExtOut_regD;
  wire   [4:0] Rs_regD;
  wire   [4:0] Rt_regD;
  wire   [4:0] wsel_regD;
  wire   [31:0] PCplus4_regD;
  wire   [15:0] branchOffset_regD;
  wire   [31:0] tempALUinB;
  wire   [31:0] ALUout;
  wire   [1:0] MemtoReg_regE;
  wire   [4:0] wsel_regE;
  wire   [1:0] ALUout_regE;
  wire   [1:0] MemtoReg_regM;
  wire   [31:0] ALUout_regM;
  wire   [4:0] wsel_regM;
  wire   [31:0] dataOut_regM;
  wire   [1:0] RegDst;
  wire   [31:0] WriteData;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [1:0] FU_Asel;
  wire   [31:0] ALUinA;
  wire   [1:0] FU_Bsel;
  wire   [1:0] PCcur;
  wire   [2:0] PCsrc;
  wire   [31:0] PCnext;
  wire   [31:0] ALUinB;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;

  DFFRX4 \PCreg_reg[2]  ( .D(PCnext[2]), .CK(clk), .RN(n147), .Q(n189), .QN(
        n94) );
  DFFRX4 \PCreg_reg[4]  ( .D(PCnext[4]), .CK(clk), .RN(n147), .Q(n188), .QN(
        n92) );
  DFFRX4 \PCreg_reg[6]  ( .D(PCnext[6]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[4]) );
  IF_DEC_regFile i_IF_DEC_regFile ( .clk(clk), .rst_n(ICACHE_ren), .flush(
        flush), .stallcache(stallcache), .stall_lw_use(stall_lw_use), 
        .instruction_next({n91, n89, ICACHE_rdata[29:0]}), .PCplus4({n39, 
        PCplus4[30:28], n38, PCplus4[26:7], n51, PCplus4[5:0]}), 
        .branchOffset(branchOffset_D), .opcode(opcode), .Rs(Rs), .Rt(Rt), .Rd(
        Rd), .shamt(shamt), .funct(funct), .immediate(immediate), 
        .PCplus4_regI(PCplus4_regI) );
  DEC_EX_regFile i_DEC_EX_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(stallcache), .MemtoReg(MemtoReg), .ALUOp(ALUOp), .JumpReg(
        JumpReg_m), .MemRead(MemRead_m), .MemWrite(MemWrite_m), .ALUsrc(ALUsrc), .RegWrite(RegWrite_m), .Branch(Branch_DEC_m), .PCplus4_regI(PCplus4_regI), 
        .funct(funct), .branchOffset_D(branchOffset_D), .A(A_f), .B(B_f), 
        .ExtOut(ExtOut), .Rs({n142, n141, n140, n139, n138}), .Rt({n137, n136, 
        n135, n134, n133}), .wsel(wsel), .MemtoReg_regD(MemtoReg_regD), 
        .ALUOp_regD(ALUOp_regD), .MemRead_regD(MemRead_regD), .MemWrite_regD(
        MemWrite_regD), .ALUsrc_regD(ALUsrc_regD), .RegWrite_regD(
        RegWrite_regD), .funct_regD(funct_regD), .A_regD(A_regD), .B_regD(
        B_regD), .ExtOut_regD(ExtOut_regD), .Rs_regD(Rs_regD), .Rt_regD(
        Rt_regD), .wsel_regD(wsel_regD), .JumpReg_regD(JumpReg_regD), 
        .Branch_regD(Branch_regD), .PCplus4_regD(PCplus4_regD), 
        .branchOffset_regD(branchOffset_regD) );
  EX_MEM_regFile i_EX_MEM_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(stallcache), .MemtoReg_regD(MemtoReg_regD), .MemRead_regD(
        MemRead_regD), .MemWrite_regD(MemWrite_regD), .RegWrite_regD(
        RegWrite_regD), .B_regD({tempALUinB[31:23], n36, tempALUinB[21:12], 
        n37, tempALUinB[10:0]}), .wsel_regD(wsel_regD), .ALUout(ALUout), 
        .MemtoReg_regE(MemtoReg_regE), .MemRead_regE(DCACHE_ren), 
        .MemWrite_regE(DCACHE_wen), .RegWrite_regE(RegWrite_regE), .B_regE(
        DCACHE_wdata), .wsel_regE(wsel_regE), .ALUout_regE({n190, n191, n192, 
        n193, n194, DCACHE_addr[24:20], n195, n196, n197, DCACHE_addr[16:15], 
        n198, DCACHE_addr[13:12], n199, n200, n201, DCACHE_addr[8], n202, 
        DCACHE_addr[6], n203, n204, n205, n206, DCACHE_addr[1], n207, 
        ALUout_regE}) );
  MEM_WB_regFile i_MEM_WB_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(stallcache), .MemtoReg_regE(MemtoReg_regE), 
        .RegWrite_regE(RegWrite_regE), .ALUout_regE({DCACHE_addr, ALUout_regE}), .wsel_regE(wsel_regE), .dataOut(DCACHE_rdata), .MemtoReg_regM(MemtoReg_regM), 
        .RegWrite_regM(RegWrite_regM), .ALUout_regM(ALUout_regM), .wsel_regM(
        wsel_regM), .dataOut_regM(dataOut_regM) );
  maincontrol i_maincontrol ( .opcode(opcode), .funct(funct), .RegDst(RegDst), 
        .MemtoReg(MemtoReg), .ALUOp(ALUOp), .Branch(Branch_DEC), .MemRead(
        MemRead), .MemWrite(MemWrite), .ALUsrc(ALUsrc), .RegWrite(RegWrite), 
        .JumpReg(JumpReg), .ExtOp(ExtOp) );
  registerFile i_registrefFile ( .clk(clk), .rst_n(ICACHE_ren), .rsel1({n142, 
        n141, n140, n139, n138}), .rsel2({n137, n136, n135, n134, n133}), 
        .wsel(wsel_regM), .wen(RegWrite_regM), .wdata({WriteData[31:12], n47, 
        WriteData[10:0]}), .rdata1(A), .rdata2(B) );
  extender i_extender ( .shamt_i(shamt), .immed_i(immediate), .ExtOp_i(ExtOp), 
        .ExtOut_o(ExtOut) );
  MUX_5_3to1 MUX_wsel ( .data0_i({n137, n136, n135, n134, n133}), .data1_i(Rd), 
        .data2_i({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .select_i(RegDst), .data_o(
        wsel) );
  MUX_32_3to1_0 MUX_WriteData ( .data0_i(dataOut_regM), .data1_i(ALUout_regM), 
        .data2_i(ALUout_regM), .select_i(MemtoReg_regM), .data_o(WriteData) );
  MUX_32_3to1_2 MUX_ALUinA ( .data0_i(A_regD), .data1_i({WriteData[31:12], n47, 
        WriteData[10:0]}), .data2_i({DCACHE_addr, ALUout_regE}), .select_i(
        FU_Asel), .data_o(ALUinA) );
  MUX_32_3to1_1 MUX_ALUinB ( .data0_i(B_regD), .data1_i({WriteData[31:12], n47, 
        WriteData[10:0]}), .data2_i({DCACHE_addr, ALUout_regE}), .select_i(
        FU_Bsel), .data_o(tempALUinB) );
  forwarding i_forwarding ( .Rs_regD(Rs_regD), .Rt_regD({Rt_regD[4:2], n88, 
        n87}), .RegWrite_regE(RegWrite_regE), .wsel_regE(wsel_regE), 
        .RegWrite_regM(RegWrite_regM), .wsel_regM(wsel_regM), .FU_Asel(FU_Asel), .FU_Bsel(FU_Bsel) );
  hazard_detection i_hazard_detection ( .Branch_EX(Branch_regD), .equal(N22), 
        .branchpred_his(branchpred_his), .JumpReg_regD(JumpReg_regD), 
        .MemRead_regD(MemRead_regD), .Rt_regD({Rt_regD[4:2], n88, n87}), .Rs({
        n142, n141, n140, n139, n138}), .Rt({n137, n136, n135, n134, n133}), 
        .ICACHE_stall(ICACHE_stall), .DCACHE_stall(DCACHE_stall), 
        .stall_lw_use(stall_lw_use), .stallcache(stallcache), .flush(flush), 
        .pred_cond(pred_cond) );
  branch_prediction i_branch_prediction ( .clk(clk), .rst_n(n147), .branch(
        Branch_regD), .equal(N22), .predict(predict), .branchpred_his(
        branchpred_his) );
  precontrolDec i_precontrolDec ( .instruction_next({n91, n89, 
        ICACHE_rdata[29:0]}), .Jump_IF(Jump_IF), .Branch_IF(Branch_IF) );
  nextPCcalculator i_nextPCcalculator ( .PCcur({ICACHE_addr[29:17], n187, 
        ICACHE_addr[15:0], PCcur}), .PCplus4({n39, PCplus4[30:28], n38, 
        PCplus4[26:7], n51, PCplus4[5:0]}), .PCplus4_regD(PCplus4_regD), 
        .targetAddr(ICACHE_rdata[25:0]), .branchOffset_I(ICACHE_rdata[15:0]), 
        .branchOffset_regD(branchOffset_regD), .JumpRegAddr({ALUinA[31], n106, 
        ALUinA[29:23], n117, ALUinA[21:20], n120, ALUinA[18:16], n115, 
        ALUinA[14], n103, ALUinA[12], n44, n111, n41, n45, n43, n40, n46, 
        ALUinA[4:0]}), .PCsrc(PCsrc), .PCnext(PCnext) );
  PCsrcLogic i_PCsrcLogic ( .pred_cond(pred_cond), .Branch_EX(Branch_regD), 
        .Branch_IF(Branch_IF), .equal(N22), .Jump(Jump_IF), .JumpReg(
        JumpReg_regD), .predict(predict), .stallcache(stallcache), 
        .stall_lw_use(stall_lw_use), .PCsrc(PCsrc) );
  ALU i_ALU ( .ALUOp_regD(ALUOp_regD), .funct_regD(funct_regD), .ALUinA({
        ALUinA[31], n106, ALUinA[29:23], n117, ALUinA[21:20], n120, 
        ALUinA[18:16], n115, ALUinA[14], n103, ALUinA[12], n44, n111, n41, n45, 
        n43, n40, n46, ALUinA[4:0]}), .ALUinB(ALUinB), .ALUout(ALUout) );
  MIPS_Pipeline_DW01_add_0 add_403 ( .A({ICACHE_addr[29:17], n187, 
        ICACHE_addr[15:14], n54, ICACHE_addr[12:3], n188, ICACHE_addr[1], n189, 
        PCcur}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .CI(1'b0), .SUM(PCplus4) );
  DFFRX1 \PCreg_reg[0]  ( .D(PCnext[0]), .CK(clk), .RN(n147), .Q(PCcur[0]) );
  DFFRX1 \PCreg_reg[1]  ( .D(PCnext[1]), .CK(clk), .RN(n147), .Q(PCcur[1]) );
  DFFRX1 \PCreg_reg[31]  ( .D(PCnext[31]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[29]) );
  DFFRX1 \PCreg_reg[10]  ( .D(PCnext[10]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[8]) );
  DFFRX1 \PCreg_reg[12]  ( .D(PCnext[12]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[10]) );
  DFFRX2 \PCreg_reg[24]  ( .D(PCnext[24]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[22]) );
  DFFRX2 \PCreg_reg[17]  ( .D(PCnext[17]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[15]) );
  DFFRX2 \PCreg_reg[26]  ( .D(PCnext[26]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[24]) );
  DFFRX1 \PCreg_reg[14]  ( .D(PCnext[14]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[12]) );
  DFFRX1 \PCreg_reg[15]  ( .D(PCnext[15]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[13]), .QN(n49) );
  DFFRX1 \PCreg_reg[18]  ( .D(PCnext[18]), .CK(clk), .RN(n147), .Q(n187), .QN(
        n48) );
  DFFRX4 \PCreg_reg[29]  ( .D(PCnext[29]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[27]) );
  DFFRX4 \PCreg_reg[28]  ( .D(PCnext[28]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[26]) );
  DFFRX2 \PCreg_reg[8]  ( .D(PCnext[8]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[6]) );
  DFFRX4 \PCreg_reg[3]  ( .D(PCnext[3]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[1]) );
  DFFRHQX8 \PCreg_reg[5]  ( .D(PCnext[5]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[3]) );
  DFFRX2 \PCreg_reg[30]  ( .D(PCnext[30]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[28]) );
  DFFRX4 \PCreg_reg[7]  ( .D(PCnext[7]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[5]) );
  DFFRX4 \PCreg_reg[21]  ( .D(PCnext[21]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[19]) );
  DFFRX2 \PCreg_reg[19]  ( .D(PCnext[19]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[17]) );
  DFFRX4 \PCreg_reg[9]  ( .D(PCnext[9]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[7]) );
  DFFRX2 \PCreg_reg[27]  ( .D(PCnext[27]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[25]) );
  DFFRX1 \PCreg_reg[25]  ( .D(PCnext[25]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[23]) );
  DFFRX2 \PCreg_reg[23]  ( .D(PCnext[23]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[21]) );
  DFFRX4 \PCreg_reg[20]  ( .D(PCnext[20]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[18]) );
  DFFRX2 \PCreg_reg[16]  ( .D(PCnext[16]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[14]) );
  DFFRX2 \PCreg_reg[13]  ( .D(PCnext[13]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[11]) );
  DFFRX4 \PCreg_reg[22]  ( .D(PCnext[22]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[20]) );
  DFFRX2 \PCreg_reg[11]  ( .D(PCnext[11]), .CK(clk), .RN(n147), .Q(
        ICACHE_addr[9]) );
  NOR4X6 U37 ( .A(n170), .B(n169), .C(n168), .D(n167), .Y(n186) );
  XOR2X2 U38 ( .A(tempALUinB[30]), .B(ALUinA[30]), .Y(n168) );
  BUFX8 U39 ( .A(tempALUinB[22]), .Y(n36) );
  BUFX4 U40 ( .A(tempALUinB[11]), .Y(n37) );
  MX2X1 U41 ( .A(ExtOut_regD[20]), .B(tempALUinB[20]), .S0(n132), .Y(
        ALUinB[20]) );
  XOR2X4 U42 ( .A(tempALUinB[20]), .B(ALUinA[20]), .Y(n178) );
  CLKMX2X8 U43 ( .A(ExtOut_regD[25]), .B(tempALUinB[25]), .S0(n132), .Y(
        ALUinB[25]) );
  INVX8 U44 ( .A(n102), .Y(n103) );
  BUFX8 U45 ( .A(PCplus4[27]), .Y(n38) );
  BUFX8 U46 ( .A(PCplus4[31]), .Y(n39) );
  BUFX16 U47 ( .A(n205), .Y(DCACHE_addr[3]) );
  CLKINVX2 U48 ( .A(tempALUinB[7]), .Y(n55) );
  MX2X1 U49 ( .A(ExtOut_regD[16]), .B(tempALUinB[16]), .S0(n132), .Y(
        ALUinB[16]) );
  CLKMX2X2 U50 ( .A(ExtOut_regD[27]), .B(tempALUinB[27]), .S0(ALUsrc_regD), 
        .Y(ALUinB[27]) );
  NAND2X2 U51 ( .A(tempALUinB[14]), .B(n64), .Y(n65) );
  CLKINVX4 U52 ( .A(ALUinA[18]), .Y(n76) );
  CLKINVX4 U53 ( .A(ALUinA[16]), .Y(n80) );
  CLKINVX4 U54 ( .A(ALUinA[25]), .Y(n68) );
  NOR4X4 U55 ( .A(n158), .B(n157), .C(n156), .D(n155), .Y(n164) );
  CLKMX2X4 U56 ( .A(ExtOut_regD[13]), .B(tempALUinB[13]), .S0(n132), .Y(
        ALUinB[13]) );
  CLKMX2X2 U57 ( .A(ExtOut_regD[29]), .B(tempALUinB[29]), .S0(n131), .Y(
        ALUinB[29]) );
  BUFX6 U58 ( .A(n204), .Y(DCACHE_addr[4]) );
  BUFX4 U59 ( .A(Rt_regD[1]), .Y(n88) );
  CLKBUFX3 U60 ( .A(WriteData[11]), .Y(n47) );
  INVX12 U61 ( .A(n96), .Y(N22) );
  NAND2X6 U62 ( .A(n97), .B(n98), .Y(n96) );
  BUFX6 U63 ( .A(ICACHE_rdata[30]), .Y(n89) );
  CLKINVX1 U64 ( .A(n94), .Y(ICACHE_addr[0]) );
  XOR2X2 U65 ( .A(tempALUinB[28]), .B(ALUinA[28]), .Y(n170) );
  BUFX8 U66 ( .A(ALUinA[6]), .Y(n40) );
  BUFX8 U67 ( .A(ALUinA[9]), .Y(n41) );
  INVX3 U68 ( .A(ALUinA[7]), .Y(n42) );
  INVX6 U69 ( .A(n42), .Y(n43) );
  BUFX8 U70 ( .A(ALUinA[11]), .Y(n44) );
  BUFX8 U71 ( .A(ALUinA[8]), .Y(n45) );
  XOR2X4 U72 ( .A(tempALUinB[9]), .B(n41), .Y(n154) );
  BUFX12 U73 ( .A(ALUinA[5]), .Y(n46) );
  XOR2X4 U74 ( .A(tempALUinB[21]), .B(ALUinA[21]), .Y(n177) );
  CLKXOR2X2 U75 ( .A(tempALUinB[6]), .B(n40), .Y(n156) );
  MX2X1 U76 ( .A(ExtOut_regD[2]), .B(tempALUinB[2]), .S0(n131), .Y(ALUinB[2])
         );
  CLKMX2X2 U77 ( .A(ExtOut_regD[26]), .B(tempALUinB[26]), .S0(n131), .Y(
        ALUinB[26]) );
  CLKMX2X2 U78 ( .A(ExtOut_regD[3]), .B(tempALUinB[3]), .S0(n131), .Y(
        ALUinB[3]) );
  XNOR2X4 U79 ( .A(tempALUinB[8]), .B(n45), .Y(n50) );
  CLKBUFX2 U80 ( .A(PCplus4[6]), .Y(n51) );
  CLKINVX1 U81 ( .A(n48), .Y(ICACHE_addr[16]) );
  INVXL U82 ( .A(n49), .Y(n54) );
  INVX4 U83 ( .A(n90), .Y(n91) );
  INVX4 U84 ( .A(ICACHE_rdata[31]), .Y(n90) );
  XOR2X2 U85 ( .A(tempALUinB[5]), .B(n46), .Y(n157) );
  AND4X8 U86 ( .A(n166), .B(n165), .C(n164), .D(n163), .Y(n97) );
  NOR4X4 U87 ( .A(n174), .B(n173), .C(n172), .D(n171), .Y(n185) );
  AND4X8 U88 ( .A(n186), .B(n185), .C(n184), .D(n183), .Y(n98) );
  XOR2X4 U89 ( .A(tempALUinB[4]), .B(ALUinA[4]), .Y(n158) );
  XOR2X2 U90 ( .A(tempALUinB[31]), .B(ALUinA[31]), .Y(n167) );
  XOR2X2 U91 ( .A(tempALUinB[29]), .B(ALUinA[29]), .Y(n169) );
  INVX1 U92 ( .A(tempALUinB[25]), .Y(n67) );
  NAND2X4 U93 ( .A(n85), .B(n86), .Y(n171) );
  NAND2X4 U94 ( .A(n59), .B(ALUinA[2]), .Y(n62) );
  XOR2X4 U95 ( .A(tempALUinB[24]), .B(ALUinA[24]), .Y(n174) );
  CLKMX2X6 U96 ( .A(ExtOut_regD[12]), .B(tempALUinB[12]), .S0(n131), .Y(
        ALUinB[12]) );
  INVX1 U97 ( .A(tempALUinB[14]), .Y(n63) );
  MX2X2 U98 ( .A(ExtOut_regD[11]), .B(n37), .S0(n131), .Y(ALUinB[11]) );
  NOR4X6 U99 ( .A(n151), .B(n148), .C(n149), .D(n150), .Y(n166) );
  CLKMX2X6 U100 ( .A(ExtOut_regD[21]), .B(tempALUinB[21]), .S0(n132), .Y(
        ALUinB[21]) );
  NAND2X4 U101 ( .A(n61), .B(n62), .Y(n160) );
  CLKXOR2X2 U102 ( .A(tempALUinB[0]), .B(ALUinA[0]), .Y(n162) );
  CLKMX2X6 U103 ( .A(ExtOut_regD[19]), .B(tempALUinB[19]), .S0(n132), .Y(
        ALUinB[19]) );
  CLKMX2X3 U104 ( .A(ExtOut_regD[0]), .B(tempALUinB[0]), .S0(n131), .Y(
        ALUinB[0]) );
  XOR2X2 U105 ( .A(tempALUinB[13]), .B(ALUinA[13]), .Y(n150) );
  NOR4X4 U106 ( .A(n177), .B(n178), .C(n176), .D(n175), .Y(n184) );
  XOR2X4 U107 ( .A(tempALUinB[15]), .B(n115), .Y(n148) );
  NAND2X2 U108 ( .A(tempALUinB[7]), .B(n56), .Y(n57) );
  NAND2X2 U109 ( .A(n55), .B(n43), .Y(n58) );
  NAND2X4 U110 ( .A(n57), .B(n58), .Y(n155) );
  INVX2 U111 ( .A(n43), .Y(n56) );
  NAND2X4 U112 ( .A(n67), .B(ALUinA[25]), .Y(n70) );
  NAND2X2 U113 ( .A(n83), .B(ALUinA[27]), .Y(n86) );
  INVX8 U114 ( .A(ALUinA[27]), .Y(n84) );
  NAND2X2 U115 ( .A(tempALUinB[2]), .B(n60), .Y(n61) );
  INVXL U116 ( .A(tempALUinB[2]), .Y(n59) );
  INVX2 U117 ( .A(ALUinA[2]), .Y(n60) );
  NAND2X2 U118 ( .A(n63), .B(ALUinA[14]), .Y(n66) );
  NAND2X4 U119 ( .A(n65), .B(n66), .Y(n149) );
  INVX2 U120 ( .A(ALUinA[14]), .Y(n64) );
  NAND2X2 U121 ( .A(tempALUinB[25]), .B(n68), .Y(n69) );
  NAND2X2 U122 ( .A(n69), .B(n70), .Y(n173) );
  XOR2X4 U123 ( .A(tempALUinB[17]), .B(ALUinA[17]), .Y(n181) );
  NAND2X2 U124 ( .A(tempALUinB[3]), .B(n72), .Y(n73) );
  NAND2X2 U125 ( .A(n71), .B(ALUinA[3]), .Y(n74) );
  NAND2X2 U126 ( .A(n73), .B(n74), .Y(n159) );
  INVXL U127 ( .A(tempALUinB[3]), .Y(n71) );
  INVX2 U128 ( .A(ALUinA[3]), .Y(n72) );
  NAND2X2 U129 ( .A(tempALUinB[18]), .B(n76), .Y(n77) );
  NAND2X2 U130 ( .A(n75), .B(ALUinA[18]), .Y(n78) );
  NAND2X4 U131 ( .A(n77), .B(n78), .Y(n180) );
  CLKINVX2 U132 ( .A(tempALUinB[18]), .Y(n75) );
  MX2X8 U133 ( .A(ExtOut_regD[23]), .B(tempALUinB[23]), .S0(n132), .Y(
        ALUinB[23]) );
  NAND2X2 U134 ( .A(tempALUinB[16]), .B(n80), .Y(n81) );
  NAND2X2 U135 ( .A(n79), .B(ALUinA[16]), .Y(n82) );
  NAND2X2 U136 ( .A(n81), .B(n82), .Y(n182) );
  CLKINVX1 U137 ( .A(tempALUinB[16]), .Y(n79) );
  NAND2X2 U138 ( .A(tempALUinB[27]), .B(n84), .Y(n85) );
  INVX1 U139 ( .A(tempALUinB[27]), .Y(n83) );
  BUFX20 U140 ( .A(ALUinA[19]), .Y(n120) );
  XOR2X4 U141 ( .A(tempALUinB[23]), .B(ALUinA[23]), .Y(n175) );
  XOR2X4 U142 ( .A(tempALUinB[19]), .B(n120), .Y(n179) );
  BUFX8 U143 ( .A(Rt_regD[0]), .Y(n87) );
  BUFX12 U144 ( .A(n206), .Y(DCACHE_addr[2]) );
  INVX6 U145 ( .A(n92), .Y(ICACHE_addr[2]) );
  XOR2X4 U146 ( .A(tempALUinB[10]), .B(n111), .Y(n153) );
  INVX4 U147 ( .A(n105), .Y(n106) );
  AND2XL U148 ( .A(MemWrite), .B(n9), .Y(MemWrite_m) );
  NOR4BX4 U149 ( .AN(n50), .B(n154), .C(n153), .D(n152), .Y(n165) );
  XOR2X2 U150 ( .A(n36), .B(n117), .Y(n176) );
  CLKINVX6 U151 ( .A(ALUinA[10]), .Y(n110) );
  BUFX12 U152 ( .A(ALUinA[15]), .Y(n115) );
  AND2XL U153 ( .A(MemRead), .B(n9), .Y(MemRead_m) );
  AND2XL U154 ( .A(JumpReg), .B(n9), .Y(JumpReg_m) );
  AND2XL U155 ( .A(Branch_DEC), .B(n9), .Y(Branch_DEC_m) );
  INVX3 U156 ( .A(n129), .Y(n126) );
  INVX3 U157 ( .A(n130), .Y(n127) );
  INVX3 U158 ( .A(n130), .Y(n125) );
  CLKBUFX3 U159 ( .A(n130), .Y(n128) );
  CLKBUFX3 U160 ( .A(n130), .Y(n129) );
  CLKINVX1 U161 ( .A(n52), .Y(n130) );
  XOR2X1 U162 ( .A(tempALUinB[12]), .B(ALUinA[12]), .Y(n151) );
  XOR2X2 U163 ( .A(n37), .B(n44), .Y(n152) );
  NOR4X4 U164 ( .A(n162), .B(n161), .C(n160), .D(n159), .Y(n163) );
  XOR2X1 U165 ( .A(tempALUinB[1]), .B(ALUinA[1]), .Y(n161) );
  NOR4X4 U166 ( .A(n182), .B(n181), .C(n180), .D(n179), .Y(n183) );
  XOR2X1 U167 ( .A(tempALUinB[26]), .B(ALUinA[26]), .Y(n172) );
  NOR2X1 U168 ( .A(stall_lw_use), .B(flush), .Y(n9) );
  CLKBUFX3 U169 ( .A(rst_n), .Y(ICACHE_ren) );
  CLKBUFX3 U170 ( .A(ALUsrc_regD), .Y(n132) );
  CLKBUFX3 U171 ( .A(ALUsrc_regD), .Y(n131) );
  NAND2BX1 U172 ( .AN(MemtoReg[0]), .B(MemtoReg[1]), .Y(n52) );
  CLKBUFX8 U173 ( .A(rst_n), .Y(n147) );
  CLKMX2X2 U174 ( .A(ExtOut_regD[28]), .B(tempALUinB[28]), .S0(n131), .Y(
        ALUinB[28]) );
  CLKMX2X2 U175 ( .A(ExtOut_regD[30]), .B(tempALUinB[30]), .S0(n132), .Y(
        ALUinB[30]) );
  INVX8 U176 ( .A(n110), .Y(n111) );
  BUFX12 U177 ( .A(ALUinA[22]), .Y(n117) );
  CLKMX2X2 U178 ( .A(ExtOut_regD[6]), .B(tempALUinB[6]), .S0(n131), .Y(
        ALUinB[6]) );
  CLKMX2X2 U179 ( .A(ExtOut_regD[15]), .B(tempALUinB[15]), .S0(n132), .Y(
        ALUinB[15]) );
  CLKMX2X2 U180 ( .A(ExtOut_regD[7]), .B(tempALUinB[7]), .S0(n131), .Y(
        ALUinB[7]) );
  CLKMX2X2 U181 ( .A(ExtOut_regD[8]), .B(tempALUinB[8]), .S0(n131), .Y(
        ALUinB[8]) );
  CLKMX2X2 U182 ( .A(ExtOut_regD[9]), .B(tempALUinB[9]), .S0(n131), .Y(
        ALUinB[9]) );
  CLKMX2X2 U183 ( .A(ExtOut_regD[10]), .B(tempALUinB[10]), .S0(n131), .Y(
        ALUinB[10]) );
  CLKMX2X2 U184 ( .A(ExtOut_regD[22]), .B(n36), .S0(n132), .Y(ALUinB[22]) );
  CLKMX2X2 U185 ( .A(ExtOut_regD[18]), .B(tempALUinB[18]), .S0(n132), .Y(
        ALUinB[18]) );
  CLKMX2X2 U186 ( .A(ExtOut_regD[17]), .B(tempALUinB[17]), .S0(n132), .Y(
        ALUinB[17]) );
  CLKMX2X2 U187 ( .A(ExtOut_regD[14]), .B(tempALUinB[14]), .S0(n132), .Y(
        ALUinB[14]) );
  CLKMX2X2 U188 ( .A(ExtOut_regD[1]), .B(tempALUinB[1]), .S0(n131), .Y(
        ALUinB[1]) );
  CLKMX2X2 U189 ( .A(ExtOut_regD[4]), .B(tempALUinB[4]), .S0(n131), .Y(
        ALUinB[4]) );
  CLKMX2X2 U190 ( .A(ExtOut_regD[5]), .B(tempALUinB[5]), .S0(n131), .Y(
        ALUinB[5]) );
  AND2X2 U191 ( .A(RegWrite), .B(n9), .Y(RegWrite_m) );
  AO22X1 U192 ( .A0(B[0]), .A1(n127), .B0(PCplus4_regI[0]), .B1(n129), .Y(
        B_f[0]) );
  AO22X1 U193 ( .A0(B[1]), .A1(n125), .B0(PCplus4_regI[1]), .B1(n128), .Y(
        B_f[1]) );
  AO22X1 U194 ( .A0(B[2]), .A1(n125), .B0(PCplus4_regI[2]), .B1(n129), .Y(
        B_f[2]) );
  AO22X1 U195 ( .A0(B[3]), .A1(n125), .B0(PCplus4_regI[3]), .B1(n128), .Y(
        B_f[3]) );
  AO22X1 U196 ( .A0(B[4]), .A1(n125), .B0(PCplus4_regI[4]), .B1(n128), .Y(
        B_f[4]) );
  AO22X1 U197 ( .A0(B[5]), .A1(n125), .B0(PCplus4_regI[5]), .B1(n129), .Y(
        B_f[5]) );
  AO22X1 U198 ( .A0(B[6]), .A1(n125), .B0(PCplus4_regI[6]), .B1(n128), .Y(
        B_f[6]) );
  AO22X1 U199 ( .A0(B[7]), .A1(n125), .B0(PCplus4_regI[7]), .B1(n128), .Y(
        B_f[7]) );
  AO22X1 U200 ( .A0(B[8]), .A1(n125), .B0(PCplus4_regI[8]), .B1(n128), .Y(
        B_f[8]) );
  AO22X1 U201 ( .A0(B[9]), .A1(n126), .B0(PCplus4_regI[9]), .B1(n129), .Y(
        B_f[9]) );
  AO22X1 U202 ( .A0(B[10]), .A1(n127), .B0(PCplus4_regI[10]), .B1(n128), .Y(
        B_f[10]) );
  AO22X1 U203 ( .A0(B[11]), .A1(n127), .B0(PCplus4_regI[11]), .B1(n129), .Y(
        B_f[11]) );
  AO22X1 U204 ( .A0(B[12]), .A1(n126), .B0(PCplus4_regI[12]), .B1(n129), .Y(
        B_f[12]) );
  AO22X1 U205 ( .A0(B[13]), .A1(n126), .B0(PCplus4_regI[13]), .B1(n128), .Y(
        B_f[13]) );
  AO22X1 U206 ( .A0(B[14]), .A1(n127), .B0(PCplus4_regI[14]), .B1(n129), .Y(
        B_f[14]) );
  AO22X1 U207 ( .A0(B[15]), .A1(n127), .B0(PCplus4_regI[15]), .B1(n128), .Y(
        B_f[15]) );
  AO22X1 U208 ( .A0(B[16]), .A1(n126), .B0(PCplus4_regI[16]), .B1(n128), .Y(
        B_f[16]) );
  AO22X1 U209 ( .A0(B[17]), .A1(n125), .B0(PCplus4_regI[17]), .B1(n128), .Y(
        B_f[17]) );
  AO22X1 U210 ( .A0(B[18]), .A1(n125), .B0(PCplus4_regI[18]), .B1(n128), .Y(
        B_f[18]) );
  AO22X1 U211 ( .A0(B[19]), .A1(n125), .B0(PCplus4_regI[19]), .B1(n128), .Y(
        B_f[19]) );
  AO22X1 U212 ( .A0(B[20]), .A1(n125), .B0(PCplus4_regI[20]), .B1(n129), .Y(
        B_f[20]) );
  AO22X1 U213 ( .A0(B[21]), .A1(n125), .B0(PCplus4_regI[21]), .B1(n129), .Y(
        B_f[21]) );
  AO22X1 U214 ( .A0(B[22]), .A1(n125), .B0(PCplus4_regI[22]), .B1(n129), .Y(
        B_f[22]) );
  AO22X1 U215 ( .A0(B[23]), .A1(n125), .B0(PCplus4_regI[23]), .B1(n129), .Y(
        B_f[23]) );
  AO22X1 U216 ( .A0(B[24]), .A1(n125), .B0(PCplus4_regI[24]), .B1(n129), .Y(
        B_f[24]) );
  AO22X1 U217 ( .A0(B[25]), .A1(n125), .B0(PCplus4_regI[25]), .B1(n129), .Y(
        B_f[25]) );
  AO22X1 U218 ( .A0(B[26]), .A1(n125), .B0(PCplus4_regI[26]), .B1(n130), .Y(
        B_f[26]) );
  AO22X1 U219 ( .A0(B[27]), .A1(n125), .B0(PCplus4_regI[27]), .B1(n128), .Y(
        B_f[27]) );
  AO22X1 U220 ( .A0(B[28]), .A1(n125), .B0(PCplus4_regI[28]), .B1(n130), .Y(
        B_f[28]) );
  AO22X1 U221 ( .A0(B[29]), .A1(n125), .B0(PCplus4_regI[29]), .B1(n128), .Y(
        B_f[29]) );
  AO22X1 U222 ( .A0(B[30]), .A1(n125), .B0(PCplus4_regI[30]), .B1(n128), .Y(
        B_f[30]) );
  AO22X1 U223 ( .A0(B[31]), .A1(n126), .B0(PCplus4_regI[31]), .B1(n128), .Y(
        B_f[31]) );
  AND2X2 U224 ( .A(A[0]), .B(n127), .Y(A_f[0]) );
  AND2X2 U225 ( .A(A[1]), .B(n127), .Y(A_f[1]) );
  AND2X2 U226 ( .A(A[2]), .B(n126), .Y(A_f[2]) );
  AND2X2 U227 ( .A(A[3]), .B(n126), .Y(A_f[3]) );
  AND2X2 U228 ( .A(A[4]), .B(n126), .Y(A_f[4]) );
  AND2X2 U229 ( .A(A[5]), .B(n126), .Y(A_f[5]) );
  AND2X2 U230 ( .A(A[6]), .B(n127), .Y(A_f[6]) );
  AND2X2 U231 ( .A(A[7]), .B(n126), .Y(A_f[7]) );
  AND2X2 U232 ( .A(A[8]), .B(n52), .Y(A_f[8]) );
  AND2X2 U233 ( .A(A[9]), .B(n52), .Y(A_f[9]) );
  AND2X2 U234 ( .A(A[10]), .B(n127), .Y(A_f[10]) );
  AND2X2 U235 ( .A(A[11]), .B(n127), .Y(A_f[11]) );
  AND2X2 U236 ( .A(A[12]), .B(n127), .Y(A_f[12]) );
  AND2X2 U237 ( .A(A[13]), .B(n127), .Y(A_f[13]) );
  AND2X2 U238 ( .A(A[14]), .B(n127), .Y(A_f[14]) );
  AND2X2 U239 ( .A(A[15]), .B(n127), .Y(A_f[15]) );
  AND2X2 U240 ( .A(A[16]), .B(n127), .Y(A_f[16]) );
  AND2X2 U241 ( .A(A[17]), .B(n127), .Y(A_f[17]) );
  AND2X2 U242 ( .A(A[18]), .B(n127), .Y(A_f[18]) );
  AND2X2 U243 ( .A(A[19]), .B(n127), .Y(A_f[19]) );
  AND2X2 U244 ( .A(A[20]), .B(n127), .Y(A_f[20]) );
  AND2X2 U245 ( .A(A[21]), .B(n127), .Y(A_f[21]) );
  AND2X2 U246 ( .A(A[22]), .B(n126), .Y(A_f[22]) );
  AND2X2 U247 ( .A(A[23]), .B(n126), .Y(A_f[23]) );
  AND2X2 U248 ( .A(A[24]), .B(n126), .Y(A_f[24]) );
  AND2X2 U249 ( .A(A[25]), .B(n126), .Y(A_f[25]) );
  AND2X2 U250 ( .A(A[26]), .B(n126), .Y(A_f[26]) );
  AND2X2 U251 ( .A(A[27]), .B(n126), .Y(A_f[27]) );
  AND2X2 U252 ( .A(A[28]), .B(n126), .Y(A_f[28]) );
  AND2X2 U253 ( .A(A[29]), .B(n126), .Y(A_f[29]) );
  AND2X2 U254 ( .A(A[30]), .B(n126), .Y(A_f[30]) );
  AND2X2 U255 ( .A(A[31]), .B(n126), .Y(A_f[31]) );
  CLKBUFX3 U256 ( .A(Rt[2]), .Y(n135) );
  CLKBUFX3 U257 ( .A(Rt[3]), .Y(n136) );
  CLKBUFX3 U258 ( .A(Rt[0]), .Y(n133) );
  CLKBUFX3 U259 ( .A(Rt[1]), .Y(n134) );
  CLKBUFX3 U260 ( .A(Rt[4]), .Y(n137) );
  CLKBUFX3 U261 ( .A(Rs[3]), .Y(n141) );
  CLKBUFX3 U262 ( .A(Rs[2]), .Y(n140) );
  CLKBUFX3 U263 ( .A(Rs[1]), .Y(n139) );
  CLKBUFX3 U264 ( .A(Rs[0]), .Y(n138) );
  CLKBUFX3 U265 ( .A(Rs[4]), .Y(n142) );
  BUFX16 U266 ( .A(n193), .Y(DCACHE_addr[26]) );
  BUFX16 U267 ( .A(n202), .Y(DCACHE_addr[7]) );
  CLKINVX1 U268 ( .A(ALUinA[13]), .Y(n102) );
  BUFX16 U269 ( .A(n199), .Y(DCACHE_addr[11]) );
  CLKINVX1 U270 ( .A(ALUinA[30]), .Y(n105) );
  BUFX16 U271 ( .A(n191), .Y(DCACHE_addr[28]) );
  BUFX16 U272 ( .A(n198), .Y(DCACHE_addr[14]) );
  BUFX16 U273 ( .A(n201), .Y(DCACHE_addr[9]) );
  BUFX16 U274 ( .A(n207), .Y(DCACHE_addr[0]) );
  BUFX16 U275 ( .A(n196), .Y(DCACHE_addr[18]) );
  BUFX16 U276 ( .A(n203), .Y(DCACHE_addr[5]) );
  BUFX16 U277 ( .A(n195), .Y(DCACHE_addr[19]) );
  BUFX16 U278 ( .A(n200), .Y(DCACHE_addr[10]) );
  BUFX16 U279 ( .A(n192), .Y(DCACHE_addr[27]) );
  CLKINVX1 U280 ( .A(n197), .Y(n121) );
  INVX16 U281 ( .A(n121), .Y(DCACHE_addr[17]) );
  BUFX16 U282 ( .A(n190), .Y(DCACHE_addr[29]) );
  BUFX16 U283 ( .A(n194), .Y(DCACHE_addr[25]) );
  CLKMX2X4 U284 ( .A(ExtOut_regD[24]), .B(tempALUinB[24]), .S0(n132), .Y(
        ALUinB[24]) );
  CLKMX2X4 U285 ( .A(ExtOut_regD[31]), .B(tempALUinB[31]), .S0(ALUsrc_regD), 
        .Y(ALUinB[31]) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1226, n1227, n1228, n1229, n1230, \blocktag[7][24] ,
         \blocktag[7][23] , \blocktag[7][22] , \blocktag[7][18] ,
         \blocktag[7][17] , \blocktag[7][14] , \blocktag[7][12] ,
         \blocktag[7][10] , \blocktag[7][6] , \blocktag[7][5] ,
         \blocktag[7][3] , \blocktag[7][2] , \blocktag[7][0] ,
         \blocktag[6][24] , \blocktag[6][23] , \blocktag[6][22] ,
         \blocktag[6][18] , \blocktag[6][17] , \blocktag[6][14] ,
         \blocktag[6][12] , \blocktag[6][10] , \blocktag[6][6] ,
         \blocktag[6][5] , \blocktag[6][3] , \blocktag[6][2] ,
         \blocktag[6][0] , \blocktag[5][24] , \blocktag[5][23] ,
         \blocktag[5][22] , \blocktag[5][18] , \blocktag[5][17] ,
         \blocktag[5][14] , \blocktag[5][12] , \blocktag[5][10] ,
         \blocktag[5][6] , \blocktag[5][5] , \blocktag[5][3] ,
         \blocktag[5][2] , \blocktag[5][0] , \blocktag[4][24] ,
         \blocktag[4][23] , \blocktag[4][22] , \blocktag[4][18] ,
         \blocktag[4][17] , \blocktag[4][14] , \blocktag[4][12] ,
         \blocktag[4][10] , \blocktag[4][6] , \blocktag[4][5] ,
         \blocktag[4][3] , \blocktag[4][2] , \blocktag[4][0] ,
         \blocktag[3][24] , \blocktag[3][23] , \blocktag[3][22] ,
         \blocktag[3][18] , \blocktag[3][17] , \blocktag[3][14] ,
         \blocktag[3][12] , \blocktag[3][10] , \blocktag[3][5] ,
         \blocktag[3][3] , \blocktag[3][2] , \blocktag[3][0] ,
         \blocktag[2][24] , \blocktag[2][23] , \blocktag[2][22] ,
         \blocktag[2][18] , \blocktag[2][17] , \blocktag[2][14] ,
         \blocktag[2][12] , \blocktag[2][10] , \blocktag[2][5] ,
         \blocktag[2][3] , \blocktag[2][2] , \blocktag[2][0] ,
         \blocktag[1][24] , \blocktag[1][23] , \blocktag[1][22] ,
         \blocktag[1][18] , \blocktag[1][17] , \blocktag[1][14] ,
         \blocktag[1][12] , \blocktag[1][10] , \blocktag[1][5] ,
         \blocktag[1][3] , \blocktag[1][2] , \blocktag[1][0] ,
         \blocktag[0][24] , \blocktag[0][23] , \blocktag[0][22] ,
         \blocktag[0][18] , \blocktag[0][17] , \blocktag[0][14] ,
         \blocktag[0][12] , \blocktag[0][10] , \blocktag[0][5] ,
         \blocktag[0][3] , \blocktag[0][2] , \blocktag[0][0] , valid, dirty,
         \block[7][127] , \block[7][126] , \block[7][125] , \block[7][124] ,
         \block[7][123] , \block[7][122] , \block[7][121] , \block[7][120] ,
         \block[7][119] , \block[7][118] , \block[7][117] , \block[7][116] ,
         \block[7][115] , \block[7][114] , \block[7][113] , \block[7][112] ,
         \block[7][111] , \block[7][110] , \block[7][109] , \block[7][108] ,
         \block[7][107] , \block[7][106] , \block[7][105] , \block[7][104] ,
         \block[7][103] , \block[7][102] , \block[7][101] , \block[7][100] ,
         \block[7][99] , \block[7][98] , \block[7][97] , \block[7][96] ,
         \block[7][95] , \block[7][94] , \block[7][93] , \block[7][92] ,
         \block[7][91] , \block[7][90] , \block[7][89] , \block[7][88] ,
         \block[7][87] , \block[7][86] , \block[7][85] , \block[7][84] ,
         \block[7][83] , \block[7][82] , \block[7][81] , \block[7][80] ,
         \block[7][79] , \block[7][78] , \block[7][77] , \block[7][76] ,
         \block[7][75] , \block[7][74] , \block[7][73] , \block[7][72] ,
         \block[7][71] , \block[7][70] , \block[7][69] , \block[7][68] ,
         \block[7][67] , \block[7][66] , \block[7][65] , \block[7][64] ,
         \block[7][63] , \block[7][62] , \block[7][61] , \block[7][60] ,
         \block[7][59] , \block[7][58] , \block[7][57] , \block[7][56] ,
         \block[7][55] , \block[7][54] , \block[7][53] , \block[7][52] ,
         \block[7][51] , \block[7][50] , \block[7][49] , \block[7][48] ,
         \block[7][47] , \block[7][46] , \block[7][45] , \block[7][44] ,
         \block[7][43] , \block[7][42] , \block[7][41] , \block[7][40] ,
         \block[7][39] , \block[7][38] , \block[7][37] , \block[7][36] ,
         \block[7][35] , \block[7][34] , \block[7][33] , \block[7][32] ,
         \block[7][31] , \block[7][30] , \block[7][29] , \block[7][28] ,
         \block[7][27] , \block[7][26] , \block[7][25] , \block[7][24] ,
         \block[7][23] , \block[7][22] , \block[7][21] , \block[7][20] ,
         \block[7][19] , \block[7][18] , \block[7][17] , \block[7][16] ,
         \block[7][15] , \block[7][14] , \block[7][13] , \block[7][12] ,
         \block[7][11] , \block[7][10] , \block[7][9] , \block[7][8] ,
         \block[7][7] , \block[7][6] , \block[7][5] , \block[7][4] ,
         \block[7][3] , \block[7][2] , \block[7][1] , \block[7][0] ,
         \block[6][127] , \block[6][126] , \block[6][125] , \block[6][124] ,
         \block[6][123] , \block[6][122] , \block[6][121] , \block[6][120] ,
         \block[6][119] , \block[6][118] , \block[6][117] , \block[6][116] ,
         \block[6][115] , \block[6][114] , \block[6][113] , \block[6][112] ,
         \block[6][111] , \block[6][110] , \block[6][109] , \block[6][108] ,
         \block[6][107] , \block[6][106] , \block[6][105] , \block[6][104] ,
         \block[6][103] , \block[6][102] , \block[6][101] , \block[6][100] ,
         \block[6][99] , \block[6][98] , \block[6][97] , \block[6][96] ,
         \block[6][95] , \block[6][94] , \block[6][93] , \block[6][92] ,
         \block[6][91] , \block[6][90] , \block[6][89] , \block[6][88] ,
         \block[6][87] , \block[6][86] , \block[6][85] , \block[6][84] ,
         \block[6][83] , \block[6][82] , \block[6][81] , \block[6][80] ,
         \block[6][79] , \block[6][78] , \block[6][77] , \block[6][76] ,
         \block[6][75] , \block[6][74] , \block[6][73] , \block[6][72] ,
         \block[6][71] , \block[6][70] , \block[6][69] , \block[6][68] ,
         \block[6][67] , \block[6][66] , \block[6][65] , \block[6][64] ,
         \block[6][63] , \block[6][62] , \block[6][61] , \block[6][60] ,
         \block[6][59] , \block[6][58] , \block[6][57] , \block[6][56] ,
         \block[6][55] , \block[6][54] , \block[6][53] , \block[6][52] ,
         \block[6][51] , \block[6][50] , \block[6][49] , \block[6][48] ,
         \block[6][47] , \block[6][46] , \block[6][45] , \block[6][44] ,
         \block[6][43] , \block[6][42] , \block[6][41] , \block[6][40] ,
         \block[6][39] , \block[6][38] , \block[6][37] , \block[6][36] ,
         \block[6][35] , \block[6][34] , \block[6][33] , \block[6][32] ,
         \block[6][31] , \block[6][30] , \block[6][29] , \block[6][28] ,
         \block[6][27] , \block[6][26] , \block[6][25] , \block[6][24] ,
         \block[6][23] , \block[6][22] , \block[6][21] , \block[6][20] ,
         \block[6][19] , \block[6][18] , \block[6][17] , \block[6][16] ,
         \block[6][15] , \block[6][14] , \block[6][13] , \block[6][12] ,
         \block[6][11] , \block[6][10] , \block[6][9] , \block[6][8] ,
         \block[6][7] , \block[6][6] , \block[6][5] , \block[6][4] ,
         \block[6][3] , \block[6][2] , \block[6][1] , \block[6][0] ,
         \block[5][127] , \block[5][126] , \block[5][125] , \block[5][124] ,
         \block[5][123] , \block[5][122] , \block[5][121] , \block[5][120] ,
         \block[5][119] , \block[5][118] , \block[5][117] , \block[5][116] ,
         \block[5][115] , \block[5][114] , \block[5][113] , \block[5][112] ,
         \block[5][111] , \block[5][110] , \block[5][109] , \block[5][108] ,
         \block[5][107] , \block[5][106] , \block[5][105] , \block[5][104] ,
         \block[5][103] , \block[5][102] , \block[5][101] , \block[5][100] ,
         \block[5][99] , \block[5][98] , \block[5][97] , \block[5][96] ,
         \block[5][95] , \block[5][94] , \block[5][93] , \block[5][92] ,
         \block[5][91] , \block[5][90] , \block[5][89] , \block[5][88] ,
         \block[5][87] , \block[5][86] , \block[5][85] , \block[5][84] ,
         \block[5][83] , \block[5][82] , \block[5][81] , \block[5][80] ,
         \block[5][79] , \block[5][78] , \block[5][77] , \block[5][76] ,
         \block[5][75] , \block[5][74] , \block[5][73] , \block[5][72] ,
         \block[5][71] , \block[5][70] , \block[5][69] , \block[5][68] ,
         \block[5][67] , \block[5][66] , \block[5][65] , \block[5][64] ,
         \block[5][63] , \block[5][62] , \block[5][61] , \block[5][60] ,
         \block[5][59] , \block[5][58] , \block[5][57] , \block[5][56] ,
         \block[5][55] , \block[5][54] , \block[5][53] , \block[5][52] ,
         \block[5][51] , \block[5][50] , \block[5][49] , \block[5][48] ,
         \block[5][47] , \block[5][46] , \block[5][45] , \block[5][44] ,
         \block[5][43] , \block[5][42] , \block[5][41] , \block[5][40] ,
         \block[5][39] , \block[5][38] , \block[5][37] , \block[5][36] ,
         \block[5][35] , \block[5][34] , \block[5][33] , \block[5][32] ,
         \block[5][31] , \block[5][30] , \block[5][29] , \block[5][28] ,
         \block[5][27] , \block[5][26] , \block[5][25] , \block[5][24] ,
         \block[5][23] , \block[5][22] , \block[5][21] , \block[5][20] ,
         \block[5][19] , \block[5][18] , \block[5][17] , \block[5][16] ,
         \block[5][15] , \block[5][14] , \block[5][13] , \block[5][12] ,
         \block[5][11] , \block[5][10] , \block[5][9] , \block[5][8] ,
         \block[5][7] , \block[5][6] , \block[5][5] , \block[5][4] ,
         \block[5][3] , \block[5][2] , \block[5][1] , \block[5][0] ,
         \block[4][127] , \block[4][126] , \block[4][125] , \block[4][124] ,
         \block[4][123] , \block[4][122] , \block[4][121] , \block[4][120] ,
         \block[4][119] , \block[4][118] , \block[4][117] , \block[4][116] ,
         \block[4][115] , \block[4][114] , \block[4][113] , \block[4][112] ,
         \block[4][111] , \block[4][110] , \block[4][109] , \block[4][108] ,
         \block[4][107] , \block[4][106] , \block[4][105] , \block[4][104] ,
         \block[4][103] , \block[4][102] , \block[4][101] , \block[4][100] ,
         \block[4][99] , \block[4][98] , \block[4][97] , \block[4][96] ,
         \block[4][95] , \block[4][94] , \block[4][93] , \block[4][92] ,
         \block[4][91] , \block[4][90] , \block[4][89] , \block[4][88] ,
         \block[4][87] , \block[4][86] , \block[4][85] , \block[4][84] ,
         \block[4][83] , \block[4][82] , \block[4][81] , \block[4][80] ,
         \block[4][79] , \block[4][78] , \block[4][77] , \block[4][76] ,
         \block[4][75] , \block[4][74] , \block[4][73] , \block[4][72] ,
         \block[4][71] , \block[4][70] , \block[4][69] , \block[4][68] ,
         \block[4][67] , \block[4][66] , \block[4][65] , \block[4][64] ,
         \block[4][63] , \block[4][62] , \block[4][61] , \block[4][60] ,
         \block[4][59] , \block[4][58] , \block[4][57] , \block[4][56] ,
         \block[4][55] , \block[4][54] , \block[4][53] , \block[4][52] ,
         \block[4][51] , \block[4][50] , \block[4][49] , \block[4][48] ,
         \block[4][47] , \block[4][46] , \block[4][45] , \block[4][44] ,
         \block[4][43] , \block[4][42] , \block[4][41] , \block[4][40] ,
         \block[4][39] , \block[4][38] , \block[4][37] , \block[4][36] ,
         \block[4][35] , \block[4][34] , \block[4][33] , \block[4][32] ,
         \block[4][31] , \block[4][30] , \block[4][29] , \block[4][28] ,
         \block[4][27] , \block[4][26] , \block[4][25] , \block[4][24] ,
         \block[4][23] , \block[4][22] , \block[4][21] , \block[4][20] ,
         \block[4][19] , \block[4][18] , \block[4][17] , \block[4][16] ,
         \block[4][15] , \block[4][14] , \block[4][13] , \block[4][12] ,
         \block[4][11] , \block[4][10] , \block[4][9] , \block[4][8] ,
         \block[4][7] , \block[4][6] , \block[4][5] , \block[4][4] ,
         \block[4][3] , \block[4][2] , \block[4][1] , \block[4][0] ,
         \block[3][127] , \block[3][126] , \block[3][125] , \block[3][124] ,
         \block[3][123] , \block[3][122] , \block[3][121] , \block[3][120] ,
         \block[3][119] , \block[3][118] , \block[3][117] , \block[3][116] ,
         \block[3][115] , \block[3][114] , \block[3][113] , \block[3][112] ,
         \block[3][111] , \block[3][110] , \block[3][109] , \block[3][108] ,
         \block[3][107] , \block[3][106] , \block[3][105] , \block[3][104] ,
         \block[3][103] , \block[3][102] , \block[3][101] , \block[3][100] ,
         \block[3][99] , \block[3][98] , \block[3][97] , \block[3][96] ,
         \block[3][95] , \block[3][94] , \block[3][93] , \block[3][92] ,
         \block[3][91] , \block[3][90] , \block[3][89] , \block[3][88] ,
         \block[3][87] , \block[3][86] , \block[3][85] , \block[3][84] ,
         \block[3][83] , \block[3][82] , \block[3][81] , \block[3][80] ,
         \block[3][79] , \block[3][78] , \block[3][77] , \block[3][76] ,
         \block[3][75] , \block[3][74] , \block[3][73] , \block[3][72] ,
         \block[3][71] , \block[3][70] , \block[3][69] , \block[3][68] ,
         \block[3][67] , \block[3][66] , \block[3][65] , \block[3][64] ,
         \block[3][63] , \block[3][62] , \block[3][61] , \block[3][60] ,
         \block[3][59] , \block[3][58] , \block[3][57] , \block[3][56] ,
         \block[3][55] , \block[3][54] , \block[3][53] , \block[3][52] ,
         \block[3][51] , \block[3][50] , \block[3][49] , \block[3][48] ,
         \block[3][47] , \block[3][46] , \block[3][45] , \block[3][44] ,
         \block[3][43] , \block[3][42] , \block[3][41] , \block[3][40] ,
         \block[3][39] , \block[3][38] , \block[3][37] , \block[3][36] ,
         \block[3][35] , \block[3][34] , \block[3][33] , \block[3][32] ,
         \block[3][31] , \block[3][30] , \block[3][29] , \block[3][28] ,
         \block[3][27] , \block[3][26] , \block[3][25] , \block[3][24] ,
         \block[3][23] , \block[3][22] , \block[3][21] , \block[3][20] ,
         \block[3][19] , \block[3][18] , \block[3][17] , \block[3][16] ,
         \block[3][15] , \block[3][14] , \block[3][13] , \block[3][12] ,
         \block[3][11] , \block[3][10] , \block[3][9] , \block[3][8] ,
         \block[3][7] , \block[3][6] , \block[3][5] , \block[3][4] ,
         \block[3][3] , \block[3][2] , \block[3][1] , \block[3][0] ,
         \block[2][127] , \block[2][126] , \block[2][125] , \block[2][124] ,
         \block[2][123] , \block[2][122] , \block[2][121] , \block[2][120] ,
         \block[2][119] , \block[2][118] , \block[2][117] , \block[2][116] ,
         \block[2][115] , \block[2][114] , \block[2][113] , \block[2][112] ,
         \block[2][111] , \block[2][110] , \block[2][109] , \block[2][108] ,
         \block[2][107] , \block[2][106] , \block[2][105] , \block[2][104] ,
         \block[2][103] , \block[2][102] , \block[2][101] , \block[2][100] ,
         \block[2][99] , \block[2][98] , \block[2][97] , \block[2][96] ,
         \block[2][95] , \block[2][94] , \block[2][93] , \block[2][92] ,
         \block[2][91] , \block[2][90] , \block[2][89] , \block[2][88] ,
         \block[2][87] , \block[2][86] , \block[2][85] , \block[2][84] ,
         \block[2][83] , \block[2][82] , \block[2][81] , \block[2][80] ,
         \block[2][79] , \block[2][78] , \block[2][77] , \block[2][76] ,
         \block[2][75] , \block[2][74] , \block[2][73] , \block[2][72] ,
         \block[2][71] , \block[2][70] , \block[2][69] , \block[2][68] ,
         \block[2][67] , \block[2][66] , \block[2][65] , \block[2][64] ,
         \block[2][63] , \block[2][62] , \block[2][61] , \block[2][60] ,
         \block[2][59] , \block[2][58] , \block[2][57] , \block[2][56] ,
         \block[2][55] , \block[2][54] , \block[2][53] , \block[2][52] ,
         \block[2][51] , \block[2][50] , \block[2][49] , \block[2][48] ,
         \block[2][47] , \block[2][46] , \block[2][45] , \block[2][44] ,
         \block[2][43] , \block[2][42] , \block[2][41] , \block[2][40] ,
         \block[2][39] , \block[2][38] , \block[2][37] , \block[2][36] ,
         \block[2][35] , \block[2][34] , \block[2][33] , \block[2][32] ,
         \block[2][31] , \block[2][30] , \block[2][29] , \block[2][28] ,
         \block[2][27] , \block[2][26] , \block[2][25] , \block[2][24] ,
         \block[2][23] , \block[2][22] , \block[2][21] , \block[2][20] ,
         \block[2][19] , \block[2][18] , \block[2][17] , \block[2][16] ,
         \block[2][15] , \block[2][14] , \block[2][13] , \block[2][12] ,
         \block[2][11] , \block[2][10] , \block[2][9] , \block[2][8] ,
         \block[2][7] , \block[2][6] , \block[2][5] , \block[2][4] ,
         \block[2][3] , \block[2][2] , \block[2][1] , \block[2][0] ,
         \block[1][127] , \block[1][126] , \block[1][125] , \block[1][124] ,
         \block[1][123] , \block[1][122] , \block[1][121] , \block[1][120] ,
         \block[1][119] , \block[1][118] , \block[1][117] , \block[1][116] ,
         \block[1][115] , \block[1][114] , \block[1][113] , \block[1][112] ,
         \block[1][111] , \block[1][110] , \block[1][109] , \block[1][108] ,
         \block[1][107] , \block[1][106] , \block[1][105] , \block[1][104] ,
         \block[1][103] , \block[1][102] , \block[1][101] , \block[1][100] ,
         \block[1][99] , \block[1][98] , \block[1][97] , \block[1][96] ,
         \block[1][95] , \block[1][94] , \block[1][93] , \block[1][92] ,
         \block[1][91] , \block[1][90] , \block[1][89] , \block[1][88] ,
         \block[1][87] , \block[1][86] , \block[1][85] , \block[1][84] ,
         \block[1][83] , \block[1][82] , \block[1][81] , \block[1][80] ,
         \block[1][79] , \block[1][78] , \block[1][77] , \block[1][76] ,
         \block[1][75] , \block[1][74] , \block[1][73] , \block[1][72] ,
         \block[1][71] , \block[1][70] , \block[1][69] , \block[1][68] ,
         \block[1][67] , \block[1][66] , \block[1][65] , \block[1][64] ,
         \block[1][63] , \block[1][62] , \block[1][61] , \block[1][60] ,
         \block[1][59] , \block[1][58] , \block[1][57] , \block[1][56] ,
         \block[1][55] , \block[1][54] , \block[1][53] , \block[1][52] ,
         \block[1][51] , \block[1][50] , \block[1][49] , \block[1][48] ,
         \block[1][47] , \block[1][46] , \block[1][45] , \block[1][44] ,
         \block[1][43] , \block[1][42] , \block[1][41] , \block[1][40] ,
         \block[1][39] , \block[1][38] , \block[1][37] , \block[1][36] ,
         \block[1][35] , \block[1][34] , \block[1][33] , \block[1][32] ,
         \block[1][31] , \block[1][30] , \block[1][29] , \block[1][28] ,
         \block[1][27] , \block[1][26] , \block[1][25] , \block[1][24] ,
         \block[1][23] , \block[1][22] , \block[1][21] , \block[1][20] ,
         \block[1][19] , \block[1][18] , \block[1][17] , \block[1][16] ,
         \block[1][15] , \block[1][14] , \block[1][13] , \block[1][12] ,
         \block[1][11] , \block[1][10] , \block[1][9] , \block[1][8] ,
         \block[1][7] , \block[1][6] , \block[1][5] , \block[1][4] ,
         \block[1][3] , \block[1][2] , \block[1][1] , \block[1][0] ,
         \block[0][127] , \block[0][126] , \block[0][125] , \block[0][124] ,
         \block[0][123] , \block[0][122] , \block[0][121] , \block[0][120] ,
         \block[0][119] , \block[0][118] , \block[0][117] , \block[0][116] ,
         \block[0][115] , \block[0][114] , \block[0][113] , \block[0][112] ,
         \block[0][111] , \block[0][110] , \block[0][109] , \block[0][108] ,
         \block[0][107] , \block[0][106] , \block[0][105] , \block[0][104] ,
         \block[0][103] , \block[0][102] , \block[0][101] , \block[0][100] ,
         \block[0][99] , \block[0][98] , \block[0][97] , \block[0][96] ,
         \block[0][95] , \block[0][94] , \block[0][93] , \block[0][92] ,
         \block[0][91] , \block[0][90] , \block[0][89] , \block[0][88] ,
         \block[0][87] , \block[0][86] , \block[0][85] , \block[0][84] ,
         \block[0][83] , \block[0][82] , \block[0][81] , \block[0][80] ,
         \block[0][79] , \block[0][78] , \block[0][77] , \block[0][76] ,
         \block[0][75] , \block[0][74] , \block[0][73] , \block[0][72] ,
         \block[0][71] , \block[0][70] , \block[0][69] , \block[0][68] ,
         \block[0][67] , \block[0][66] , \block[0][65] , \block[0][64] ,
         \block[0][63] , \block[0][62] , \block[0][61] , \block[0][60] ,
         \block[0][59] , \block[0][58] , \block[0][57] , \block[0][56] ,
         \block[0][55] , \block[0][54] , \block[0][53] , \block[0][52] ,
         \block[0][51] , \block[0][50] , \block[0][49] , \block[0][48] ,
         \block[0][47] , \block[0][46] , \block[0][45] , \block[0][44] ,
         \block[0][43] , \block[0][42] , \block[0][41] , \block[0][40] ,
         \block[0][39] , \block[0][38] , \block[0][37] , \block[0][36] ,
         \block[0][35] , \block[0][34] , \block[0][33] , \block[0][32] ,
         \block[0][31] , \block[0][30] , \block[0][29] , \block[0][28] ,
         \block[0][27] , \block[0][26] , \block[0][25] , \block[0][24] ,
         \block[0][23] , \block[0][22] , \block[0][21] , \block[0][20] ,
         \block[0][19] , \block[0][18] , \block[0][17] , \block[0][16] ,
         \block[0][15] , \block[0][14] , \block[0][13] , \block[0][12] ,
         \block[0][11] , \block[0][10] , \block[0][9] , \block[0][8] ,
         \block[0][7] , \block[0][6] , \block[0][5] , \block[0][4] ,
         \block[0][3] , \block[0][2] , \block[0][1] , \block[0][0] , n140,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n503, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n128, n129, n133, n134,
         n135, n136, n137, n138, n139, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n502, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n800, n801, n802, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  EDFFX1 \block_reg[7][127]  ( .D(block_next[127]), .E(n731), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFX1 \block_reg[7][126]  ( .D(block_next[126]), .E(n732), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFX1 \block_reg[7][125]  ( .D(block_next[125]), .E(n731), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFX1 \block_reg[7][124]  ( .D(block_next[124]), .E(n738), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFX1 \block_reg[7][123]  ( .D(block_next[123]), .E(n736), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFX1 \block_reg[7][122]  ( .D(block_next[122]), .E(n737), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFX1 \block_reg[7][121]  ( .D(block_next[121]), .E(n735), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFX1 \block_reg[7][120]  ( .D(block_next[120]), .E(n734), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFX1 \block_reg[7][119]  ( .D(block_next[119]), .E(n736), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFX1 \block_reg[7][118]  ( .D(block_next[118]), .E(n733), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFX1 \block_reg[7][117]  ( .D(block_next[117]), .E(n737), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFX1 \block_reg[7][116]  ( .D(block_next[116]), .E(n735), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFX1 \block_reg[7][115]  ( .D(block_next[115]), .E(n734), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFX1 \block_reg[7][114]  ( .D(block_next[114]), .E(n736), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFX1 \block_reg[7][113]  ( .D(block_next[113]), .E(n733), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFX1 \block_reg[7][112]  ( .D(block_next[112]), .E(n243), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFX1 \block_reg[7][111]  ( .D(block_next[111]), .E(n731), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFX1 \block_reg[7][110]  ( .D(block_next[110]), .E(n732), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFX1 \block_reg[7][109]  ( .D(block_next[109]), .E(n738), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFX1 \block_reg[7][108]  ( .D(block_next[108]), .E(n738), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFX1 \block_reg[7][107]  ( .D(block_next[107]), .E(n737), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFX1 \block_reg[7][106]  ( .D(block_next[106]), .E(n735), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFX1 \block_reg[7][105]  ( .D(block_next[105]), .E(n734), .CK(clk), .Q(
        \block[7][105] ) );
  EDFFX1 \block_reg[7][104]  ( .D(block_next[104]), .E(n735), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFX1 \block_reg[7][103]  ( .D(block_next[103]), .E(n734), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFX1 \block_reg[7][102]  ( .D(block_next[102]), .E(n736), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFX1 \block_reg[7][101]  ( .D(block_next[101]), .E(n733), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFX1 \block_reg[7][100]  ( .D(block_next[100]), .E(n243), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFX1 \block_reg[7][99]  ( .D(block_next[99]), .E(n731), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFX1 \block_reg[7][98]  ( .D(block_next[98]), .E(n732), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFX1 \block_reg[7][97]  ( .D(block_next[97]), .E(n738), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFX1 \block_reg[7][96]  ( .D(block_next[96]), .E(n737), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFX1 \block_reg[7][95]  ( .D(block_next[95]), .E(n735), .CK(clk), .Q(
        \block[7][95] ) );
  EDFFX1 \block_reg[7][94]  ( .D(block_next[94]), .E(n734), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFX1 \block_reg[7][93]  ( .D(block_next[93]), .E(n736), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFX1 \block_reg[7][92]  ( .D(block_next[92]), .E(n733), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFX1 \block_reg[7][91]  ( .D(block_next[91]), .E(n738), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFX1 \block_reg[7][90]  ( .D(block_next[90]), .E(n738), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFX1 \block_reg[7][89]  ( .D(block_next[89]), .E(n738), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFX1 \block_reg[7][88]  ( .D(block_next[88]), .E(n738), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFX1 \block_reg[7][87]  ( .D(block_next[87]), .E(n738), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFX1 \block_reg[7][86]  ( .D(block_next[86]), .E(n738), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFX1 \block_reg[7][85]  ( .D(block_next[85]), .E(n738), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFX1 \block_reg[7][84]  ( .D(block_next[84]), .E(n738), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFX1 \block_reg[7][83]  ( .D(block_next[83]), .E(n738), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFX1 \block_reg[7][82]  ( .D(block_next[82]), .E(n738), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFX1 \block_reg[7][81]  ( .D(block_next[81]), .E(n738), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFX1 \block_reg[7][80]  ( .D(block_next[80]), .E(n738), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFX1 \block_reg[7][79]  ( .D(block_next[79]), .E(n738), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFX1 \block_reg[7][78]  ( .D(block_next[78]), .E(n737), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFX1 \block_reg[7][77]  ( .D(block_next[77]), .E(n737), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFX1 \block_reg[7][76]  ( .D(block_next[76]), .E(n737), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFX1 \block_reg[7][75]  ( .D(block_next[75]), .E(n737), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFX1 \block_reg[7][74]  ( .D(block_next[74]), .E(n737), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFX1 \block_reg[7][73]  ( .D(block_next[73]), .E(n737), .CK(clk), .Q(
        \block[7][73] ) );
  EDFFX1 \block_reg[7][72]  ( .D(block_next[72]), .E(n737), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFX1 \block_reg[7][71]  ( .D(block_next[71]), .E(n737), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFX1 \block_reg[7][70]  ( .D(block_next[70]), .E(n737), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFX1 \block_reg[7][69]  ( .D(block_next[69]), .E(n737), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFX1 \block_reg[7][68]  ( .D(block_next[68]), .E(n737), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFX1 \block_reg[7][67]  ( .D(block_next[67]), .E(n737), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFX1 \block_reg[7][66]  ( .D(block_next[66]), .E(n737), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFX1 \block_reg[7][65]  ( .D(block_next[65]), .E(n736), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFX1 \block_reg[7][64]  ( .D(block_next[64]), .E(n736), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFX1 \block_reg[7][63]  ( .D(block_next[63]), .E(n736), .CK(clk), .Q(
        \block[7][63] ) );
  EDFFX1 \block_reg[7][62]  ( .D(block_next[62]), .E(n736), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFX1 \block_reg[7][61]  ( .D(block_next[61]), .E(n736), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFX1 \block_reg[7][60]  ( .D(block_next[60]), .E(n736), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFX1 \block_reg[7][59]  ( .D(block_next[59]), .E(n736), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFX1 \block_reg[7][58]  ( .D(block_next[58]), .E(n736), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFX1 \block_reg[7][57]  ( .D(block_next[57]), .E(n736), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFX1 \block_reg[7][56]  ( .D(block_next[56]), .E(n736), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFX1 \block_reg[7][55]  ( .D(block_next[55]), .E(n736), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFX1 \block_reg[7][54]  ( .D(block_next[54]), .E(n736), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n736), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n735), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[7][51]  ( .D(block_next[51]), .E(n735), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFX1 \block_reg[7][50]  ( .D(block_next[50]), .E(n735), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n735), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[7][48]  ( .D(block_next[48]), .E(n735), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFX1 \block_reg[7][47]  ( .D(block_next[47]), .E(n735), .CK(clk), .Q(
        \block[7][47] ) );
  EDFFX1 \block_reg[7][46]  ( .D(block_next[46]), .E(n735), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFX1 \block_reg[7][45]  ( .D(block_next[45]), .E(n735), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFX1 \block_reg[7][44]  ( .D(block_next[44]), .E(n735), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFX1 \block_reg[7][43]  ( .D(block_next[43]), .E(n735), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFX1 \block_reg[7][42]  ( .D(block_next[42]), .E(n735), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n735), .CK(clk), .Q(
        \block[7][41] ) );
  EDFFX1 \block_reg[7][40]  ( .D(block_next[40]), .E(n735), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFX1 \block_reg[7][39]  ( .D(block_next[39]), .E(n734), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n734), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n734), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n734), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n734), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n734), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFX1 \block_reg[7][33]  ( .D(block_next[33]), .E(n734), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n734), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[7][31]  ( .D(block_next[31]), .E(n734), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFX1 \block_reg[7][30]  ( .D(block_next[30]), .E(n734), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFX1 \block_reg[7][29]  ( .D(block_next[29]), .E(n734), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFX1 \block_reg[7][28]  ( .D(block_next[28]), .E(n734), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFX1 \block_reg[7][27]  ( .D(block_next[27]), .E(n734), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFX1 \block_reg[7][26]  ( .D(block_next[26]), .E(n733), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFX1 \block_reg[7][25]  ( .D(block_next[25]), .E(n733), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFX1 \block_reg[7][24]  ( .D(block_next[24]), .E(n733), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFX1 \block_reg[7][23]  ( .D(block_next[23]), .E(n733), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFX1 \block_reg[7][22]  ( .D(block_next[22]), .E(n733), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFX1 \block_reg[7][21]  ( .D(block_next[21]), .E(n733), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFX1 \block_reg[7][20]  ( .D(block_next[20]), .E(n733), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFX1 \block_reg[7][19]  ( .D(block_next[19]), .E(n733), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFX1 \block_reg[7][18]  ( .D(block_next[18]), .E(n733), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFX1 \block_reg[7][17]  ( .D(block_next[17]), .E(n733), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFX1 \block_reg[7][16]  ( .D(block_next[16]), .E(n733), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFX1 \block_reg[7][15]  ( .D(block_next[15]), .E(n733), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFX1 \block_reg[7][14]  ( .D(block_next[14]), .E(n733), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFX1 \block_reg[7][13]  ( .D(block_next[13]), .E(n732), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFX1 \block_reg[7][12]  ( .D(block_next[12]), .E(n732), .CK(clk), .Q(
        \block[7][12] ) );
  EDFFX1 \block_reg[7][11]  ( .D(block_next[11]), .E(n732), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFX1 \block_reg[7][10]  ( .D(block_next[10]), .E(n732), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFX1 \block_reg[7][9]  ( .D(block_next[9]), .E(n732), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFX1 \block_reg[7][8]  ( .D(block_next[8]), .E(n732), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFX1 \block_reg[7][7]  ( .D(block_next[7]), .E(n732), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFX1 \block_reg[7][6]  ( .D(block_next[6]), .E(n732), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFX1 \block_reg[7][5]  ( .D(block_next[5]), .E(n732), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFX1 \block_reg[7][4]  ( .D(block_next[4]), .E(n732), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFX1 \block_reg[7][3]  ( .D(block_next[3]), .E(n732), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFX1 \block_reg[7][2]  ( .D(block_next[2]), .E(n732), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFX1 \block_reg[7][1]  ( .D(block_next[1]), .E(n732), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFX1 \block_reg[7][0]  ( .D(block_next[0]), .E(n243), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFX1 \block_reg[3][127]  ( .D(block_next[127]), .E(n767), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFX1 \block_reg[3][126]  ( .D(block_next[126]), .E(n767), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFX1 \block_reg[3][125]  ( .D(block_next[125]), .E(n766), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFX1 \block_reg[3][124]  ( .D(block_next[124]), .E(n768), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFX1 \block_reg[3][123]  ( .D(block_next[123]), .E(n769), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFX1 \block_reg[3][122]  ( .D(block_next[122]), .E(n764), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFX1 \block_reg[3][121]  ( .D(block_next[121]), .E(n763), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFX1 \block_reg[3][120]  ( .D(block_next[120]), .E(n765), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFX1 \block_reg[3][119]  ( .D(block_next[119]), .E(n770), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFX1 \block_reg[3][118]  ( .D(block_next[118]), .E(n765), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFX1 \block_reg[3][117]  ( .D(block_next[117]), .E(n769), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFX1 \block_reg[3][116]  ( .D(block_next[116]), .E(n764), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFX1 \block_reg[3][115]  ( .D(block_next[115]), .E(n763), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFX1 \block_reg[3][114]  ( .D(block_next[114]), .E(n765), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFX1 \block_reg[3][113]  ( .D(block_next[113]), .E(n770), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFX1 \block_reg[3][112]  ( .D(block_next[112]), .E(n239), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFX1 \block_reg[3][111]  ( .D(block_next[111]), .E(n768), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFX1 \block_reg[3][110]  ( .D(block_next[110]), .E(n767), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFX1 \block_reg[3][109]  ( .D(block_next[109]), .E(n766), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFX1 \block_reg[3][108]  ( .D(block_next[108]), .E(n768), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFX1 \block_reg[3][107]  ( .D(block_next[107]), .E(n769), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFX1 \block_reg[3][106]  ( .D(block_next[106]), .E(n764), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFX1 \block_reg[3][105]  ( .D(block_next[105]), .E(n763), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFX1 \block_reg[3][104]  ( .D(block_next[104]), .E(n770), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFX1 \block_reg[3][103]  ( .D(block_next[103]), .E(n770), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFX1 \block_reg[3][102]  ( .D(block_next[102]), .E(n770), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFX1 \block_reg[3][101]  ( .D(block_next[101]), .E(n770), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFX1 \block_reg[3][100]  ( .D(block_next[100]), .E(n770), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFX1 \block_reg[3][99]  ( .D(block_next[99]), .E(n770), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFX1 \block_reg[3][98]  ( .D(block_next[98]), .E(n770), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFX1 \block_reg[3][97]  ( .D(block_next[97]), .E(n770), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFX1 \block_reg[3][96]  ( .D(block_next[96]), .E(n770), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFX1 \block_reg[3][95]  ( .D(block_next[95]), .E(n770), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFX1 \block_reg[3][94]  ( .D(block_next[94]), .E(n770), .CK(clk), .Q(
        \block[3][94] ) );
  EDFFX1 \block_reg[3][93]  ( .D(block_next[93]), .E(n770), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFX1 \block_reg[3][92]  ( .D(block_next[92]), .E(n770), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFX1 \block_reg[3][91]  ( .D(block_next[91]), .E(n769), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFX1 \block_reg[3][90]  ( .D(block_next[90]), .E(n769), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFX1 \block_reg[3][89]  ( .D(block_next[89]), .E(n769), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFX1 \block_reg[3][88]  ( .D(block_next[88]), .E(n769), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFX1 \block_reg[3][87]  ( .D(block_next[87]), .E(n769), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFX1 \block_reg[3][86]  ( .D(block_next[86]), .E(n769), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFX1 \block_reg[3][85]  ( .D(block_next[85]), .E(n769), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFX1 \block_reg[3][84]  ( .D(block_next[84]), .E(n769), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFX1 \block_reg[3][83]  ( .D(block_next[83]), .E(n769), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFX1 \block_reg[3][82]  ( .D(block_next[82]), .E(n769), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFX1 \block_reg[3][81]  ( .D(block_next[81]), .E(n769), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFX1 \block_reg[3][80]  ( .D(block_next[80]), .E(n769), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFX1 \block_reg[3][79]  ( .D(block_next[79]), .E(n769), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFX1 \block_reg[3][78]  ( .D(block_next[78]), .E(n764), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFX1 \block_reg[3][77]  ( .D(block_next[77]), .E(n763), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFX1 \block_reg[3][76]  ( .D(block_next[76]), .E(n765), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFX1 \block_reg[3][75]  ( .D(block_next[75]), .E(n770), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFX1 \block_reg[3][74]  ( .D(block_next[74]), .E(n239), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFX1 \block_reg[3][73]  ( .D(block_next[73]), .E(n767), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFX1 \block_reg[3][72]  ( .D(block_next[72]), .E(n766), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFX1 \block_reg[3][71]  ( .D(block_next[71]), .E(n768), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFX1 \block_reg[3][70]  ( .D(block_next[70]), .E(n769), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFX1 \block_reg[3][69]  ( .D(block_next[69]), .E(n764), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFX1 \block_reg[3][68]  ( .D(block_next[68]), .E(n763), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFX1 \block_reg[3][67]  ( .D(block_next[67]), .E(n765), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFX1 \block_reg[3][66]  ( .D(block_next[66]), .E(n770), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFX1 \block_reg[3][65]  ( .D(block_next[65]), .E(n768), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFX1 \block_reg[3][64]  ( .D(block_next[64]), .E(n768), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[3][63]  ( .D(block_next[63]), .E(n768), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFX1 \block_reg[3][62]  ( .D(block_next[62]), .E(n768), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFX1 \block_reg[3][61]  ( .D(block_next[61]), .E(n768), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFX1 \block_reg[3][60]  ( .D(block_next[60]), .E(n768), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFX1 \block_reg[3][59]  ( .D(block_next[59]), .E(n768), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFX1 \block_reg[3][58]  ( .D(block_next[58]), .E(n768), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFX1 \block_reg[3][57]  ( .D(block_next[57]), .E(n768), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFX1 \block_reg[3][56]  ( .D(block_next[56]), .E(n768), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFX1 \block_reg[3][55]  ( .D(block_next[55]), .E(n768), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFX1 \block_reg[3][54]  ( .D(block_next[54]), .E(n768), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n768), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n767), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[3][51]  ( .D(block_next[51]), .E(n767), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFX1 \block_reg[3][50]  ( .D(block_next[50]), .E(n767), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n767), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[3][48]  ( .D(block_next[48]), .E(n767), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFX1 \block_reg[3][47]  ( .D(block_next[47]), .E(n767), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFX1 \block_reg[3][46]  ( .D(block_next[46]), .E(n767), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFX1 \block_reg[3][45]  ( .D(block_next[45]), .E(n767), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFX1 \block_reg[3][44]  ( .D(block_next[44]), .E(n767), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFX1 \block_reg[3][43]  ( .D(block_next[43]), .E(n767), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFX1 \block_reg[3][42]  ( .D(block_next[42]), .E(n767), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n767), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[3][40]  ( .D(block_next[40]), .E(n767), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFX1 \block_reg[3][39]  ( .D(block_next[39]), .E(n766), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n766), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n766), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n766), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n766), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n766), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[3][33]  ( .D(block_next[33]), .E(n766), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n766), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[3][31]  ( .D(block_next[31]), .E(n766), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFX1 \block_reg[3][30]  ( .D(block_next[30]), .E(n766), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFX1 \block_reg[3][29]  ( .D(block_next[29]), .E(n766), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFX1 \block_reg[3][28]  ( .D(block_next[28]), .E(n766), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFX1 \block_reg[3][27]  ( .D(block_next[27]), .E(n766), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFX1 \block_reg[3][26]  ( .D(block_next[26]), .E(n239), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFX1 \block_reg[3][25]  ( .D(block_next[25]), .E(n239), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFX1 \block_reg[3][24]  ( .D(block_next[24]), .E(n239), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFX1 \block_reg[3][23]  ( .D(block_next[23]), .E(n766), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFX1 \block_reg[3][22]  ( .D(block_next[22]), .E(n767), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFX1 \block_reg[3][21]  ( .D(block_next[21]), .E(n766), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n768), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFX1 \block_reg[3][19]  ( .D(block_next[19]), .E(n769), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFX1 \block_reg[3][18]  ( .D(block_next[18]), .E(n764), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFX1 \block_reg[3][17]  ( .D(block_next[17]), .E(n763), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFX1 \block_reg[3][16]  ( .D(block_next[16]), .E(n765), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFX1 \block_reg[3][15]  ( .D(block_next[15]), .E(n770), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFX1 \block_reg[3][14]  ( .D(block_next[14]), .E(n770), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFX1 \block_reg[3][13]  ( .D(block_next[13]), .E(n765), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFX1 \block_reg[3][12]  ( .D(block_next[12]), .E(n765), .CK(clk), .Q(
        \block[3][12] ) );
  EDFFX1 \block_reg[3][11]  ( .D(block_next[11]), .E(n765), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFX1 \block_reg[3][10]  ( .D(block_next[10]), .E(n765), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFX1 \block_reg[3][9]  ( .D(block_next[9]), .E(n765), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFX1 \block_reg[3][8]  ( .D(block_next[8]), .E(n765), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFX1 \block_reg[3][7]  ( .D(block_next[7]), .E(n765), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFX1 \block_reg[3][6]  ( .D(block_next[6]), .E(n765), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFX1 \block_reg[3][5]  ( .D(block_next[5]), .E(n765), .CK(clk), .Q(
        \block[3][5] ) );
  EDFFX1 \block_reg[3][4]  ( .D(block_next[4]), .E(n765), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFX1 \block_reg[3][3]  ( .D(block_next[3]), .E(n765), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFX1 \block_reg[3][2]  ( .D(block_next[2]), .E(n765), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFX1 \block_reg[3][1]  ( .D(block_next[1]), .E(n765), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFX1 \block_reg[3][0]  ( .D(block_next[0]), .E(n764), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFX1 \block_reg[5][127]  ( .D(block_next[127]), .E(n751), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFX1 \block_reg[5][126]  ( .D(block_next[126]), .E(n751), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFX1 \block_reg[5][125]  ( .D(block_next[125]), .E(n750), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFX1 \block_reg[5][124]  ( .D(block_next[124]), .E(n752), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFX1 \block_reg[5][123]  ( .D(block_next[123]), .E(n753), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFX1 \block_reg[5][122]  ( .D(block_next[122]), .E(n748), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFX1 \block_reg[5][121]  ( .D(block_next[121]), .E(n747), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFX1 \block_reg[5][120]  ( .D(block_next[120]), .E(n749), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFX1 \block_reg[5][119]  ( .D(block_next[119]), .E(n754), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFX1 \block_reg[5][118]  ( .D(block_next[118]), .E(n749), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFX1 \block_reg[5][117]  ( .D(block_next[117]), .E(n753), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFX1 \block_reg[5][116]  ( .D(block_next[116]), .E(n748), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFX1 \block_reg[5][115]  ( .D(block_next[115]), .E(n747), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFX1 \block_reg[5][114]  ( .D(block_next[114]), .E(n749), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFX1 \block_reg[5][113]  ( .D(block_next[113]), .E(n754), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFX1 \block_reg[5][112]  ( .D(block_next[112]), .E(n241), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFX1 \block_reg[5][111]  ( .D(block_next[111]), .E(n752), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFX1 \block_reg[5][110]  ( .D(block_next[110]), .E(n751), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFX1 \block_reg[5][109]  ( .D(block_next[109]), .E(n750), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFX1 \block_reg[5][108]  ( .D(block_next[108]), .E(n752), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFX1 \block_reg[5][107]  ( .D(block_next[107]), .E(n753), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFX1 \block_reg[5][106]  ( .D(block_next[106]), .E(n748), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFX1 \block_reg[5][105]  ( .D(block_next[105]), .E(n747), .CK(clk), .Q(
        \block[5][105] ) );
  EDFFX1 \block_reg[5][104]  ( .D(block_next[104]), .E(n754), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFX1 \block_reg[5][103]  ( .D(block_next[103]), .E(n754), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFX1 \block_reg[5][102]  ( .D(block_next[102]), .E(n754), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFX1 \block_reg[5][101]  ( .D(block_next[101]), .E(n754), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFX1 \block_reg[5][100]  ( .D(block_next[100]), .E(n754), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFX1 \block_reg[5][99]  ( .D(block_next[99]), .E(n754), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFX1 \block_reg[5][98]  ( .D(block_next[98]), .E(n754), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFX1 \block_reg[5][97]  ( .D(block_next[97]), .E(n754), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFX1 \block_reg[5][96]  ( .D(block_next[96]), .E(n754), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFX1 \block_reg[5][95]  ( .D(block_next[95]), .E(n754), .CK(clk), .Q(
        \block[5][95] ) );
  EDFFX1 \block_reg[5][94]  ( .D(block_next[94]), .E(n754), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFX1 \block_reg[5][93]  ( .D(block_next[93]), .E(n754), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFX1 \block_reg[5][92]  ( .D(block_next[92]), .E(n754), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFX1 \block_reg[5][91]  ( .D(block_next[91]), .E(n753), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFX1 \block_reg[5][90]  ( .D(block_next[90]), .E(n753), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFX1 \block_reg[5][89]  ( .D(block_next[89]), .E(n753), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFX1 \block_reg[5][88]  ( .D(block_next[88]), .E(n753), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFX1 \block_reg[5][87]  ( .D(block_next[87]), .E(n753), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFX1 \block_reg[5][86]  ( .D(block_next[86]), .E(n753), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFX1 \block_reg[5][85]  ( .D(block_next[85]), .E(n753), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFX1 \block_reg[5][84]  ( .D(block_next[84]), .E(n753), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFX1 \block_reg[5][83]  ( .D(block_next[83]), .E(n753), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFX1 \block_reg[5][82]  ( .D(block_next[82]), .E(n753), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFX1 \block_reg[5][81]  ( .D(block_next[81]), .E(n753), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFX1 \block_reg[5][80]  ( .D(block_next[80]), .E(n753), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFX1 \block_reg[5][79]  ( .D(block_next[79]), .E(n753), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFX1 \block_reg[5][78]  ( .D(block_next[78]), .E(n748), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFX1 \block_reg[5][77]  ( .D(block_next[77]), .E(n747), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFX1 \block_reg[5][76]  ( .D(block_next[76]), .E(n749), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFX1 \block_reg[5][75]  ( .D(block_next[75]), .E(n754), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFX1 \block_reg[5][74]  ( .D(block_next[74]), .E(n241), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFX1 \block_reg[5][73]  ( .D(block_next[73]), .E(n751), .CK(clk), .Q(
        \block[5][73] ) );
  EDFFX1 \block_reg[5][72]  ( .D(block_next[72]), .E(n750), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFX1 \block_reg[5][71]  ( .D(block_next[71]), .E(n752), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFX1 \block_reg[5][70]  ( .D(block_next[70]), .E(n753), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFX1 \block_reg[5][69]  ( .D(block_next[69]), .E(n748), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFX1 \block_reg[5][68]  ( .D(block_next[68]), .E(n747), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFX1 \block_reg[5][67]  ( .D(block_next[67]), .E(n749), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFX1 \block_reg[5][66]  ( .D(block_next[66]), .E(n754), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFX1 \block_reg[5][65]  ( .D(block_next[65]), .E(n752), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFX1 \block_reg[5][64]  ( .D(block_next[64]), .E(n752), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFX1 \block_reg[5][63]  ( .D(block_next[63]), .E(n752), .CK(clk), .Q(
        \block[5][63] ) );
  EDFFX1 \block_reg[5][62]  ( .D(block_next[62]), .E(n752), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFX1 \block_reg[5][61]  ( .D(block_next[61]), .E(n752), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFX1 \block_reg[5][60]  ( .D(block_next[60]), .E(n752), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFX1 \block_reg[5][59]  ( .D(block_next[59]), .E(n752), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFX1 \block_reg[5][58]  ( .D(block_next[58]), .E(n752), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFX1 \block_reg[5][57]  ( .D(block_next[57]), .E(n752), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFX1 \block_reg[5][56]  ( .D(block_next[56]), .E(n752), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFX1 \block_reg[5][55]  ( .D(block_next[55]), .E(n752), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFX1 \block_reg[5][54]  ( .D(block_next[54]), .E(n752), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFX1 \block_reg[5][53]  ( .D(block_next[53]), .E(n752), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFX1 \block_reg[5][52]  ( .D(block_next[52]), .E(n751), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFX1 \block_reg[5][51]  ( .D(block_next[51]), .E(n751), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFX1 \block_reg[5][50]  ( .D(block_next[50]), .E(n751), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFX1 \block_reg[5][49]  ( .D(block_next[49]), .E(n751), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFX1 \block_reg[5][48]  ( .D(block_next[48]), .E(n751), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFX1 \block_reg[5][47]  ( .D(block_next[47]), .E(n751), .CK(clk), .Q(
        \block[5][47] ) );
  EDFFX1 \block_reg[5][46]  ( .D(block_next[46]), .E(n751), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFX1 \block_reg[5][45]  ( .D(block_next[45]), .E(n751), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFX1 \block_reg[5][44]  ( .D(block_next[44]), .E(n751), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFX1 \block_reg[5][43]  ( .D(block_next[43]), .E(n751), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFX1 \block_reg[5][42]  ( .D(block_next[42]), .E(n751), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n751), .CK(clk), .Q(
        \block[5][41] ) );
  EDFFX1 \block_reg[5][40]  ( .D(block_next[40]), .E(n751), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFX1 \block_reg[5][39]  ( .D(block_next[39]), .E(n750), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n750), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n750), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n750), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFX1 \block_reg[5][35]  ( .D(block_next[35]), .E(n750), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFX1 \block_reg[5][34]  ( .D(block_next[34]), .E(n750), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFX1 \block_reg[5][33]  ( .D(block_next[33]), .E(n750), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n750), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFX1 \block_reg[5][31]  ( .D(block_next[31]), .E(n750), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFX1 \block_reg[5][30]  ( .D(block_next[30]), .E(n750), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFX1 \block_reg[5][29]  ( .D(block_next[29]), .E(n750), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFX1 \block_reg[5][28]  ( .D(block_next[28]), .E(n750), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFX1 \block_reg[5][27]  ( .D(block_next[27]), .E(n750), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFX1 \block_reg[5][26]  ( .D(block_next[26]), .E(n241), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFX1 \block_reg[5][25]  ( .D(block_next[25]), .E(n241), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFX1 \block_reg[5][24]  ( .D(block_next[24]), .E(n241), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFX1 \block_reg[5][23]  ( .D(block_next[23]), .E(n750), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFX1 \block_reg[5][22]  ( .D(block_next[22]), .E(n751), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFX1 \block_reg[5][21]  ( .D(block_next[21]), .E(n750), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[5][20]  ( .D(block_next[20]), .E(n752), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFX1 \block_reg[5][19]  ( .D(block_next[19]), .E(n753), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFX1 \block_reg[5][18]  ( .D(block_next[18]), .E(n748), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFX1 \block_reg[5][17]  ( .D(block_next[17]), .E(n747), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFX1 \block_reg[5][16]  ( .D(block_next[16]), .E(n749), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFX1 \block_reg[5][15]  ( .D(block_next[15]), .E(n754), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[5][14]  ( .D(block_next[14]), .E(n754), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFX1 \block_reg[5][13]  ( .D(block_next[13]), .E(n749), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFX1 \block_reg[5][12]  ( .D(block_next[12]), .E(n749), .CK(clk), .Q(
        \block[5][12] ) );
  EDFFX1 \block_reg[5][11]  ( .D(block_next[11]), .E(n749), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFX1 \block_reg[5][10]  ( .D(block_next[10]), .E(n749), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFX1 \block_reg[5][9]  ( .D(block_next[9]), .E(n749), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFX1 \block_reg[5][8]  ( .D(block_next[8]), .E(n749), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFX1 \block_reg[5][7]  ( .D(block_next[7]), .E(n749), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFX1 \block_reg[5][6]  ( .D(block_next[6]), .E(n749), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFX1 \block_reg[5][5]  ( .D(block_next[5]), .E(n749), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFX1 \block_reg[5][4]  ( .D(block_next[4]), .E(n749), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFX1 \block_reg[5][3]  ( .D(block_next[3]), .E(n749), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFX1 \block_reg[5][2]  ( .D(block_next[2]), .E(n749), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFX1 \block_reg[5][1]  ( .D(block_next[1]), .E(n749), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFX1 \block_reg[5][0]  ( .D(block_next[0]), .E(n748), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFX1 \block_reg[1][127]  ( .D(block_next[127]), .E(n783), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFX1 \block_reg[1][126]  ( .D(block_next[126]), .E(n783), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFX1 \block_reg[1][125]  ( .D(block_next[125]), .E(n782), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFX1 \block_reg[1][124]  ( .D(block_next[124]), .E(n784), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFX1 \block_reg[1][123]  ( .D(block_next[123]), .E(n785), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFX1 \block_reg[1][122]  ( .D(block_next[122]), .E(n780), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFX1 \block_reg[1][121]  ( .D(block_next[121]), .E(n779), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFX1 \block_reg[1][120]  ( .D(block_next[120]), .E(n781), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFX1 \block_reg[1][119]  ( .D(block_next[119]), .E(n786), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFX1 \block_reg[1][118]  ( .D(block_next[118]), .E(n781), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFX1 \block_reg[1][117]  ( .D(block_next[117]), .E(n785), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFX1 \block_reg[1][116]  ( .D(block_next[116]), .E(n780), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFX1 \block_reg[1][115]  ( .D(block_next[115]), .E(n779), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFX1 \block_reg[1][114]  ( .D(block_next[114]), .E(n781), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFX1 \block_reg[1][113]  ( .D(block_next[113]), .E(n786), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFX1 \block_reg[1][112]  ( .D(block_next[112]), .E(n237), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFX1 \block_reg[1][111]  ( .D(block_next[111]), .E(n784), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFX1 \block_reg[1][110]  ( .D(block_next[110]), .E(n783), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFX1 \block_reg[1][109]  ( .D(block_next[109]), .E(n782), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFX1 \block_reg[1][108]  ( .D(block_next[108]), .E(n784), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFX1 \block_reg[1][107]  ( .D(block_next[107]), .E(n785), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFX1 \block_reg[1][106]  ( .D(block_next[106]), .E(n780), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFX1 \block_reg[1][105]  ( .D(block_next[105]), .E(n779), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFX1 \block_reg[1][104]  ( .D(block_next[104]), .E(n786), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFX1 \block_reg[1][103]  ( .D(block_next[103]), .E(n786), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFX1 \block_reg[1][102]  ( .D(block_next[102]), .E(n786), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFX1 \block_reg[1][101]  ( .D(block_next[101]), .E(n786), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFX1 \block_reg[1][100]  ( .D(block_next[100]), .E(n786), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFX1 \block_reg[1][99]  ( .D(block_next[99]), .E(n786), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFX1 \block_reg[1][98]  ( .D(block_next[98]), .E(n786), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFX1 \block_reg[1][97]  ( .D(block_next[97]), .E(n786), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFX1 \block_reg[1][96]  ( .D(block_next[96]), .E(n786), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFX1 \block_reg[1][95]  ( .D(block_next[95]), .E(n786), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFX1 \block_reg[1][94]  ( .D(block_next[94]), .E(n786), .CK(clk), .Q(
        \block[1][94] ) );
  EDFFX1 \block_reg[1][93]  ( .D(block_next[93]), .E(n786), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFX1 \block_reg[1][92]  ( .D(block_next[92]), .E(n786), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFX1 \block_reg[1][91]  ( .D(block_next[91]), .E(n785), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFX1 \block_reg[1][90]  ( .D(block_next[90]), .E(n785), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFX1 \block_reg[1][89]  ( .D(block_next[89]), .E(n785), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFX1 \block_reg[1][88]  ( .D(block_next[88]), .E(n785), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFX1 \block_reg[1][87]  ( .D(block_next[87]), .E(n785), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFX1 \block_reg[1][86]  ( .D(block_next[86]), .E(n785), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFX1 \block_reg[1][85]  ( .D(block_next[85]), .E(n785), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFX1 \block_reg[1][84]  ( .D(block_next[84]), .E(n785), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFX1 \block_reg[1][83]  ( .D(block_next[83]), .E(n785), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFX1 \block_reg[1][82]  ( .D(block_next[82]), .E(n785), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFX1 \block_reg[1][81]  ( .D(block_next[81]), .E(n785), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFX1 \block_reg[1][80]  ( .D(block_next[80]), .E(n785), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFX1 \block_reg[1][79]  ( .D(block_next[79]), .E(n785), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFX1 \block_reg[1][78]  ( .D(block_next[78]), .E(n780), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFX1 \block_reg[1][77]  ( .D(block_next[77]), .E(n779), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFX1 \block_reg[1][76]  ( .D(block_next[76]), .E(n781), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFX1 \block_reg[1][75]  ( .D(block_next[75]), .E(n786), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFX1 \block_reg[1][74]  ( .D(block_next[74]), .E(n237), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFX1 \block_reg[1][73]  ( .D(block_next[73]), .E(n783), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFX1 \block_reg[1][72]  ( .D(block_next[72]), .E(n782), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFX1 \block_reg[1][71]  ( .D(block_next[71]), .E(n784), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFX1 \block_reg[1][70]  ( .D(block_next[70]), .E(n785), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFX1 \block_reg[1][69]  ( .D(block_next[69]), .E(n780), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFX1 \block_reg[1][68]  ( .D(block_next[68]), .E(n779), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFX1 \block_reg[1][67]  ( .D(block_next[67]), .E(n781), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFX1 \block_reg[1][66]  ( .D(block_next[66]), .E(n786), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFX1 \block_reg[1][65]  ( .D(block_next[65]), .E(n784), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFX1 \block_reg[1][64]  ( .D(block_next[64]), .E(n784), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[1][63]  ( .D(block_next[63]), .E(n784), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFX1 \block_reg[1][62]  ( .D(block_next[62]), .E(n784), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFX1 \block_reg[1][61]  ( .D(block_next[61]), .E(n784), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFX1 \block_reg[1][60]  ( .D(block_next[60]), .E(n784), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFX1 \block_reg[1][59]  ( .D(block_next[59]), .E(n784), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFX1 \block_reg[1][58]  ( .D(block_next[58]), .E(n784), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFX1 \block_reg[1][57]  ( .D(block_next[57]), .E(n784), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFX1 \block_reg[1][56]  ( .D(block_next[56]), .E(n784), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFX1 \block_reg[1][55]  ( .D(block_next[55]), .E(n784), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFX1 \block_reg[1][54]  ( .D(block_next[54]), .E(n784), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n784), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n783), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[1][51]  ( .D(block_next[51]), .E(n783), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFX1 \block_reg[1][50]  ( .D(block_next[50]), .E(n783), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n783), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[1][48]  ( .D(block_next[48]), .E(n783), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFX1 \block_reg[1][47]  ( .D(block_next[47]), .E(n783), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFX1 \block_reg[1][46]  ( .D(block_next[46]), .E(n783), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFX1 \block_reg[1][45]  ( .D(block_next[45]), .E(n783), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFX1 \block_reg[1][44]  ( .D(block_next[44]), .E(n783), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFX1 \block_reg[1][43]  ( .D(block_next[43]), .E(n783), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFX1 \block_reg[1][42]  ( .D(block_next[42]), .E(n783), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFX1 \block_reg[1][41]  ( .D(block_next[41]), .E(n783), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[1][40]  ( .D(block_next[40]), .E(n783), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFX1 \block_reg[1][39]  ( .D(block_next[39]), .E(n782), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFX1 \block_reg[1][38]  ( .D(block_next[38]), .E(n782), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFX1 \block_reg[1][37]  ( .D(block_next[37]), .E(n782), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[1][36]  ( .D(block_next[36]), .E(n782), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(n782), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFX1 \block_reg[1][34]  ( .D(block_next[34]), .E(n782), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFX1 \block_reg[1][33]  ( .D(block_next[33]), .E(n782), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFX1 \block_reg[1][32]  ( .D(block_next[32]), .E(n782), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[1][31]  ( .D(block_next[31]), .E(n782), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFX1 \block_reg[1][30]  ( .D(block_next[30]), .E(n782), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFX1 \block_reg[1][29]  ( .D(block_next[29]), .E(n782), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFX1 \block_reg[1][28]  ( .D(block_next[28]), .E(n782), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFX1 \block_reg[1][27]  ( .D(block_next[27]), .E(n782), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFX1 \block_reg[1][26]  ( .D(block_next[26]), .E(n237), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFX1 \block_reg[1][25]  ( .D(block_next[25]), .E(n237), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFX1 \block_reg[1][24]  ( .D(block_next[24]), .E(n237), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFX1 \block_reg[1][23]  ( .D(block_next[23]), .E(n782), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFX1 \block_reg[1][22]  ( .D(block_next[22]), .E(n783), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFX1 \block_reg[1][21]  ( .D(block_next[21]), .E(n782), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n784), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFX1 \block_reg[1][19]  ( .D(block_next[19]), .E(n785), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFX1 \block_reg[1][18]  ( .D(block_next[18]), .E(n780), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFX1 \block_reg[1][17]  ( .D(block_next[17]), .E(n779), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFX1 \block_reg[1][16]  ( .D(block_next[16]), .E(n781), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFX1 \block_reg[1][15]  ( .D(block_next[15]), .E(n786), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFX1 \block_reg[1][14]  ( .D(block_next[14]), .E(n786), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFX1 \block_reg[1][13]  ( .D(block_next[13]), .E(n781), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFX1 \block_reg[1][12]  ( .D(block_next[12]), .E(n781), .CK(clk), .Q(
        \block[1][12] ) );
  EDFFX1 \block_reg[1][11]  ( .D(block_next[11]), .E(n781), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFX1 \block_reg[1][10]  ( .D(block_next[10]), .E(n781), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFX1 \block_reg[1][9]  ( .D(block_next[9]), .E(n781), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFX1 \block_reg[1][8]  ( .D(block_next[8]), .E(n781), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFX1 \block_reg[1][7]  ( .D(block_next[7]), .E(n781), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFX1 \block_reg[1][6]  ( .D(block_next[6]), .E(n781), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFX1 \block_reg[1][5]  ( .D(block_next[5]), .E(n781), .CK(clk), .Q(
        \block[1][5] ) );
  EDFFX1 \block_reg[1][4]  ( .D(block_next[4]), .E(n781), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFX1 \block_reg[1][3]  ( .D(block_next[3]), .E(n781), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFX1 \block_reg[1][2]  ( .D(block_next[2]), .E(n781), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFX1 \block_reg[1][1]  ( .D(block_next[1]), .E(n781), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFX1 \block_reg[1][0]  ( .D(block_next[0]), .E(n780), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFX1 \block_reg[4][127]  ( .D(block_next[127]), .E(n759), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFX1 \block_reg[4][126]  ( .D(block_next[126]), .E(n759), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFX1 \block_reg[4][125]  ( .D(block_next[125]), .E(n758), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFX1 \block_reg[4][124]  ( .D(block_next[124]), .E(n760), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFX1 \block_reg[4][123]  ( .D(block_next[123]), .E(n761), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFX1 \block_reg[4][122]  ( .D(block_next[122]), .E(n756), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFX1 \block_reg[4][121]  ( .D(block_next[121]), .E(n755), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFX1 \block_reg[4][120]  ( .D(block_next[120]), .E(n757), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFX1 \block_reg[4][119]  ( .D(block_next[119]), .E(n762), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFX1 \block_reg[4][118]  ( .D(block_next[118]), .E(n757), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFX1 \block_reg[4][117]  ( .D(block_next[117]), .E(n761), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFX1 \block_reg[4][116]  ( .D(block_next[116]), .E(n756), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFX1 \block_reg[4][115]  ( .D(block_next[115]), .E(n755), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFX1 \block_reg[4][114]  ( .D(block_next[114]), .E(n757), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFX1 \block_reg[4][113]  ( .D(block_next[113]), .E(n762), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFX1 \block_reg[4][112]  ( .D(block_next[112]), .E(n240), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFX1 \block_reg[4][111]  ( .D(block_next[111]), .E(n760), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFX1 \block_reg[4][110]  ( .D(block_next[110]), .E(n759), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFX1 \block_reg[4][109]  ( .D(block_next[109]), .E(n758), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFX1 \block_reg[4][108]  ( .D(block_next[108]), .E(n760), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFX1 \block_reg[4][107]  ( .D(block_next[107]), .E(n761), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFX1 \block_reg[4][106]  ( .D(block_next[106]), .E(n756), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFX1 \block_reg[4][105]  ( .D(block_next[105]), .E(n755), .CK(clk), .Q(
        \block[4][105] ) );
  EDFFX1 \block_reg[4][104]  ( .D(block_next[104]), .E(n762), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFX1 \block_reg[4][103]  ( .D(block_next[103]), .E(n762), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFX1 \block_reg[4][102]  ( .D(block_next[102]), .E(n762), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFX1 \block_reg[4][101]  ( .D(block_next[101]), .E(n762), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFX1 \block_reg[4][100]  ( .D(block_next[100]), .E(n762), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFX1 \block_reg[4][99]  ( .D(block_next[99]), .E(n762), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFX1 \block_reg[4][98]  ( .D(block_next[98]), .E(n762), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFX1 \block_reg[4][97]  ( .D(block_next[97]), .E(n762), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFX1 \block_reg[4][96]  ( .D(block_next[96]), .E(n762), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFX1 \block_reg[4][95]  ( .D(block_next[95]), .E(n762), .CK(clk), .Q(
        \block[4][95] ) );
  EDFFX1 \block_reg[4][94]  ( .D(block_next[94]), .E(n762), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFX1 \block_reg[4][93]  ( .D(block_next[93]), .E(n762), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFX1 \block_reg[4][92]  ( .D(block_next[92]), .E(n762), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFX1 \block_reg[4][91]  ( .D(block_next[91]), .E(n761), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFX1 \block_reg[4][90]  ( .D(block_next[90]), .E(n761), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFX1 \block_reg[4][89]  ( .D(block_next[89]), .E(n761), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFX1 \block_reg[4][88]  ( .D(block_next[88]), .E(n761), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFX1 \block_reg[4][87]  ( .D(block_next[87]), .E(n761), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFX1 \block_reg[4][86]  ( .D(block_next[86]), .E(n761), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFX1 \block_reg[4][85]  ( .D(block_next[85]), .E(n761), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFX1 \block_reg[4][84]  ( .D(block_next[84]), .E(n761), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFX1 \block_reg[4][83]  ( .D(block_next[83]), .E(n761), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFX1 \block_reg[4][82]  ( .D(block_next[82]), .E(n761), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFX1 \block_reg[4][81]  ( .D(block_next[81]), .E(n761), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFX1 \block_reg[4][80]  ( .D(block_next[80]), .E(n761), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFX1 \block_reg[4][79]  ( .D(block_next[79]), .E(n761), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFX1 \block_reg[4][78]  ( .D(block_next[78]), .E(n756), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFX1 \block_reg[4][77]  ( .D(block_next[77]), .E(n755), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFX1 \block_reg[4][76]  ( .D(block_next[76]), .E(n757), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFX1 \block_reg[4][75]  ( .D(block_next[75]), .E(n762), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFX1 \block_reg[4][74]  ( .D(block_next[74]), .E(n240), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFX1 \block_reg[4][73]  ( .D(block_next[73]), .E(n759), .CK(clk), .Q(
        \block[4][73] ) );
  EDFFX1 \block_reg[4][72]  ( .D(block_next[72]), .E(n758), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFX1 \block_reg[4][71]  ( .D(block_next[71]), .E(n760), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFX1 \block_reg[4][70]  ( .D(block_next[70]), .E(n761), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFX1 \block_reg[4][69]  ( .D(block_next[69]), .E(n756), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFX1 \block_reg[4][68]  ( .D(block_next[68]), .E(n755), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFX1 \block_reg[4][67]  ( .D(block_next[67]), .E(n757), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFX1 \block_reg[4][66]  ( .D(block_next[66]), .E(n762), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFX1 \block_reg[4][65]  ( .D(block_next[65]), .E(n760), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFX1 \block_reg[4][64]  ( .D(block_next[64]), .E(n760), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFX1 \block_reg[4][63]  ( .D(block_next[63]), .E(n760), .CK(clk), .Q(
        \block[4][63] ) );
  EDFFX1 \block_reg[4][62]  ( .D(block_next[62]), .E(n760), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFX1 \block_reg[4][61]  ( .D(block_next[61]), .E(n760), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFX1 \block_reg[4][60]  ( .D(block_next[60]), .E(n760), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFX1 \block_reg[4][59]  ( .D(block_next[59]), .E(n760), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFX1 \block_reg[4][58]  ( .D(block_next[58]), .E(n760), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFX1 \block_reg[4][57]  ( .D(block_next[57]), .E(n760), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFX1 \block_reg[4][56]  ( .D(block_next[56]), .E(n760), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFX1 \block_reg[4][55]  ( .D(block_next[55]), .E(n760), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFX1 \block_reg[4][54]  ( .D(block_next[54]), .E(n760), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n760), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n759), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[4][51]  ( .D(block_next[51]), .E(n759), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFX1 \block_reg[4][50]  ( .D(block_next[50]), .E(n759), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n759), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[4][48]  ( .D(block_next[48]), .E(n759), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFX1 \block_reg[4][47]  ( .D(block_next[47]), .E(n759), .CK(clk), .Q(
        \block[4][47] ) );
  EDFFX1 \block_reg[4][46]  ( .D(block_next[46]), .E(n759), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFX1 \block_reg[4][45]  ( .D(block_next[45]), .E(n759), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFX1 \block_reg[4][44]  ( .D(block_next[44]), .E(n759), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFX1 \block_reg[4][43]  ( .D(block_next[43]), .E(n759), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFX1 \block_reg[4][42]  ( .D(block_next[42]), .E(n759), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n759), .CK(clk), .Q(
        \block[4][41] ) );
  EDFFX1 \block_reg[4][40]  ( .D(block_next[40]), .E(n759), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFX1 \block_reg[4][39]  ( .D(block_next[39]), .E(n758), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n758), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n758), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n758), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n758), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFX1 \block_reg[4][34]  ( .D(block_next[34]), .E(n758), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFX1 \block_reg[4][33]  ( .D(block_next[33]), .E(n758), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n758), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[4][31]  ( .D(block_next[31]), .E(n758), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFX1 \block_reg[4][30]  ( .D(block_next[30]), .E(n758), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFX1 \block_reg[4][29]  ( .D(block_next[29]), .E(n758), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFX1 \block_reg[4][28]  ( .D(block_next[28]), .E(n758), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFX1 \block_reg[4][27]  ( .D(block_next[27]), .E(n758), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFX1 \block_reg[4][26]  ( .D(block_next[26]), .E(n240), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFX1 \block_reg[4][25]  ( .D(block_next[25]), .E(n240), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFX1 \block_reg[4][24]  ( .D(block_next[24]), .E(n240), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFX1 \block_reg[4][23]  ( .D(block_next[23]), .E(n758), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFX1 \block_reg[4][22]  ( .D(block_next[22]), .E(n759), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFX1 \block_reg[4][21]  ( .D(block_next[21]), .E(n758), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n760), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFX1 \block_reg[4][19]  ( .D(block_next[19]), .E(n761), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFX1 \block_reg[4][18]  ( .D(block_next[18]), .E(n756), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFX1 \block_reg[4][17]  ( .D(block_next[17]), .E(n755), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFX1 \block_reg[4][16]  ( .D(block_next[16]), .E(n757), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFX1 \block_reg[4][15]  ( .D(block_next[15]), .E(n762), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFX1 \block_reg[4][14]  ( .D(block_next[14]), .E(n762), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFX1 \block_reg[4][13]  ( .D(block_next[13]), .E(n757), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFX1 \block_reg[4][12]  ( .D(block_next[12]), .E(n757), .CK(clk), .Q(
        \block[4][12] ) );
  EDFFX1 \block_reg[4][11]  ( .D(block_next[11]), .E(n757), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFX1 \block_reg[4][10]  ( .D(block_next[10]), .E(n757), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFX1 \block_reg[4][9]  ( .D(block_next[9]), .E(n757), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFX1 \block_reg[4][8]  ( .D(block_next[8]), .E(n757), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFX1 \block_reg[4][7]  ( .D(block_next[7]), .E(n757), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFX1 \block_reg[4][6]  ( .D(block_next[6]), .E(n757), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFX1 \block_reg[4][5]  ( .D(block_next[5]), .E(n757), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFX1 \block_reg[4][4]  ( .D(block_next[4]), .E(n757), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFX1 \block_reg[4][3]  ( .D(block_next[3]), .E(n757), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFX1 \block_reg[4][2]  ( .D(block_next[2]), .E(n757), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFX1 \block_reg[4][1]  ( .D(block_next[1]), .E(n757), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFX1 \block_reg[4][0]  ( .D(block_next[0]), .E(n756), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFX1 \block_reg[0][127]  ( .D(block_next[127]), .E(n791), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFX1 \block_reg[0][126]  ( .D(block_next[126]), .E(n791), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFX1 \block_reg[0][125]  ( .D(block_next[125]), .E(n790), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFX1 \block_reg[0][124]  ( .D(block_next[124]), .E(n792), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFX1 \block_reg[0][123]  ( .D(block_next[123]), .E(n793), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFX1 \block_reg[0][122]  ( .D(block_next[122]), .E(n788), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFX1 \block_reg[0][121]  ( .D(block_next[121]), .E(n787), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFX1 \block_reg[0][120]  ( .D(block_next[120]), .E(n789), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFX1 \block_reg[0][119]  ( .D(block_next[119]), .E(n794), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFX1 \block_reg[0][118]  ( .D(block_next[118]), .E(n789), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFX1 \block_reg[0][117]  ( .D(block_next[117]), .E(n793), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFX1 \block_reg[0][116]  ( .D(block_next[116]), .E(n788), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFX1 \block_reg[0][115]  ( .D(block_next[115]), .E(n787), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFX1 \block_reg[0][114]  ( .D(block_next[114]), .E(n789), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFX1 \block_reg[0][113]  ( .D(block_next[113]), .E(n794), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFX1 \block_reg[0][112]  ( .D(block_next[112]), .E(n236), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFX1 \block_reg[0][111]  ( .D(block_next[111]), .E(n792), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFX1 \block_reg[0][110]  ( .D(block_next[110]), .E(n791), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFX1 \block_reg[0][109]  ( .D(block_next[109]), .E(n790), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFX1 \block_reg[0][108]  ( .D(block_next[108]), .E(n792), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFX1 \block_reg[0][107]  ( .D(block_next[107]), .E(n793), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFX1 \block_reg[0][106]  ( .D(block_next[106]), .E(n788), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFX1 \block_reg[0][105]  ( .D(block_next[105]), .E(n787), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFX1 \block_reg[0][104]  ( .D(block_next[104]), .E(n794), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFX1 \block_reg[0][103]  ( .D(block_next[103]), .E(n794), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFX1 \block_reg[0][102]  ( .D(block_next[102]), .E(n794), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFX1 \block_reg[0][101]  ( .D(block_next[101]), .E(n794), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFX1 \block_reg[0][100]  ( .D(block_next[100]), .E(n794), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFX1 \block_reg[0][99]  ( .D(block_next[99]), .E(n794), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFX1 \block_reg[0][98]  ( .D(block_next[98]), .E(n794), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFX1 \block_reg[0][97]  ( .D(block_next[97]), .E(n794), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFX1 \block_reg[0][96]  ( .D(block_next[96]), .E(n794), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFX1 \block_reg[0][95]  ( .D(block_next[95]), .E(n794), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFX1 \block_reg[0][94]  ( .D(block_next[94]), .E(n794), .CK(clk), .Q(
        \block[0][94] ) );
  EDFFX1 \block_reg[0][93]  ( .D(block_next[93]), .E(n794), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFX1 \block_reg[0][92]  ( .D(block_next[92]), .E(n794), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFX1 \block_reg[0][91]  ( .D(block_next[91]), .E(n793), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFX1 \block_reg[0][90]  ( .D(block_next[90]), .E(n793), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFX1 \block_reg[0][89]  ( .D(block_next[89]), .E(n793), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFX1 \block_reg[0][88]  ( .D(block_next[88]), .E(n793), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFX1 \block_reg[0][87]  ( .D(block_next[87]), .E(n793), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFX1 \block_reg[0][86]  ( .D(block_next[86]), .E(n793), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFX1 \block_reg[0][85]  ( .D(block_next[85]), .E(n793), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFX1 \block_reg[0][84]  ( .D(block_next[84]), .E(n793), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFX1 \block_reg[0][83]  ( .D(block_next[83]), .E(n793), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFX1 \block_reg[0][82]  ( .D(block_next[82]), .E(n793), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFX1 \block_reg[0][81]  ( .D(block_next[81]), .E(n793), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFX1 \block_reg[0][80]  ( .D(block_next[80]), .E(n793), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFX1 \block_reg[0][79]  ( .D(block_next[79]), .E(n793), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFX1 \block_reg[0][78]  ( .D(block_next[78]), .E(n788), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFX1 \block_reg[0][77]  ( .D(block_next[77]), .E(n787), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFX1 \block_reg[0][76]  ( .D(block_next[76]), .E(n789), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFX1 \block_reg[0][75]  ( .D(block_next[75]), .E(n794), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFX1 \block_reg[0][74]  ( .D(block_next[74]), .E(n236), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFX1 \block_reg[0][73]  ( .D(block_next[73]), .E(n791), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFX1 \block_reg[0][72]  ( .D(block_next[72]), .E(n790), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFX1 \block_reg[0][71]  ( .D(block_next[71]), .E(n792), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFX1 \block_reg[0][70]  ( .D(block_next[70]), .E(n793), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFX1 \block_reg[0][69]  ( .D(block_next[69]), .E(n788), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFX1 \block_reg[0][68]  ( .D(block_next[68]), .E(n787), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFX1 \block_reg[0][67]  ( .D(block_next[67]), .E(n789), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFX1 \block_reg[0][66]  ( .D(block_next[66]), .E(n794), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFX1 \block_reg[0][65]  ( .D(block_next[65]), .E(n792), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFX1 \block_reg[0][64]  ( .D(block_next[64]), .E(n792), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[0][63]  ( .D(block_next[63]), .E(n792), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFX1 \block_reg[0][62]  ( .D(block_next[62]), .E(n792), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFX1 \block_reg[0][61]  ( .D(block_next[61]), .E(n792), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFX1 \block_reg[0][60]  ( .D(block_next[60]), .E(n792), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFX1 \block_reg[0][59]  ( .D(block_next[59]), .E(n792), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFX1 \block_reg[0][58]  ( .D(block_next[58]), .E(n792), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFX1 \block_reg[0][57]  ( .D(block_next[57]), .E(n792), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFX1 \block_reg[0][56]  ( .D(block_next[56]), .E(n792), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFX1 \block_reg[0][55]  ( .D(block_next[55]), .E(n792), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFX1 \block_reg[0][54]  ( .D(block_next[54]), .E(n792), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n792), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n791), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[0][51]  ( .D(block_next[51]), .E(n791), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFX1 \block_reg[0][50]  ( .D(block_next[50]), .E(n791), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n791), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[0][48]  ( .D(block_next[48]), .E(n791), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFX1 \block_reg[0][47]  ( .D(block_next[47]), .E(n791), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFX1 \block_reg[0][46]  ( .D(block_next[46]), .E(n791), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFX1 \block_reg[0][45]  ( .D(block_next[45]), .E(n791), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFX1 \block_reg[0][44]  ( .D(block_next[44]), .E(n791), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFX1 \block_reg[0][43]  ( .D(block_next[43]), .E(n791), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFX1 \block_reg[0][42]  ( .D(block_next[42]), .E(n791), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n791), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[0][40]  ( .D(block_next[40]), .E(n791), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFX1 \block_reg[0][39]  ( .D(block_next[39]), .E(n790), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n790), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n790), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n790), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n790), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[0][34]  ( .D(block_next[34]), .E(n790), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFX1 \block_reg[0][33]  ( .D(block_next[33]), .E(n790), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n790), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[0][31]  ( .D(block_next[31]), .E(n790), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFX1 \block_reg[0][30]  ( .D(block_next[30]), .E(n790), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFX1 \block_reg[0][29]  ( .D(block_next[29]), .E(n790), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFX1 \block_reg[0][28]  ( .D(block_next[28]), .E(n790), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFX1 \block_reg[0][27]  ( .D(block_next[27]), .E(n790), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFX1 \block_reg[0][26]  ( .D(block_next[26]), .E(n236), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFX1 \block_reg[0][25]  ( .D(block_next[25]), .E(n236), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFX1 \block_reg[0][24]  ( .D(block_next[24]), .E(n236), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFX1 \block_reg[0][23]  ( .D(block_next[23]), .E(n790), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFX1 \block_reg[0][22]  ( .D(block_next[22]), .E(n791), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFX1 \block_reg[0][21]  ( .D(block_next[21]), .E(n790), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n792), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFX1 \block_reg[0][19]  ( .D(block_next[19]), .E(n793), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFX1 \block_reg[0][18]  ( .D(block_next[18]), .E(n788), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFX1 \block_reg[0][17]  ( .D(block_next[17]), .E(n787), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFX1 \block_reg[0][16]  ( .D(block_next[16]), .E(n789), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFX1 \block_reg[0][15]  ( .D(block_next[15]), .E(n794), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFX1 \block_reg[0][14]  ( .D(block_next[14]), .E(n794), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFX1 \block_reg[0][13]  ( .D(block_next[13]), .E(n789), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFX1 \block_reg[0][12]  ( .D(block_next[12]), .E(n789), .CK(clk), .Q(
        \block[0][12] ) );
  EDFFX1 \block_reg[0][11]  ( .D(block_next[11]), .E(n789), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFX1 \block_reg[0][10]  ( .D(block_next[10]), .E(n789), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFX1 \block_reg[0][9]  ( .D(block_next[9]), .E(n789), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFX1 \block_reg[0][8]  ( .D(block_next[8]), .E(n789), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFX1 \block_reg[0][7]  ( .D(block_next[7]), .E(n789), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFX1 \block_reg[0][6]  ( .D(block_next[6]), .E(n789), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFX1 \block_reg[0][5]  ( .D(block_next[5]), .E(n789), .CK(clk), .Q(
        \block[0][5] ) );
  EDFFX1 \block_reg[0][4]  ( .D(block_next[4]), .E(n789), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFX1 \block_reg[0][3]  ( .D(block_next[3]), .E(n789), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFX1 \block_reg[0][2]  ( .D(block_next[2]), .E(n789), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFX1 \block_reg[0][1]  ( .D(block_next[1]), .E(n789), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFX1 \block_reg[0][0]  ( .D(block_next[0]), .E(n788), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFX1 \block_reg[6][127]  ( .D(block_next[127]), .E(n739), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFX1 \block_reg[6][126]  ( .D(block_next[126]), .E(n740), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFX1 \block_reg[6][125]  ( .D(block_next[125]), .E(n739), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFX1 \block_reg[6][124]  ( .D(block_next[124]), .E(n746), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFX1 \block_reg[6][123]  ( .D(block_next[123]), .E(n744), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFX1 \block_reg[6][122]  ( .D(block_next[122]), .E(n745), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFX1 \block_reg[6][121]  ( .D(block_next[121]), .E(n743), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFX1 \block_reg[6][120]  ( .D(block_next[120]), .E(n742), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFX1 \block_reg[6][119]  ( .D(block_next[119]), .E(n744), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFX1 \block_reg[6][118]  ( .D(block_next[118]), .E(n741), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFX1 \block_reg[6][117]  ( .D(block_next[117]), .E(n745), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFX1 \block_reg[6][116]  ( .D(block_next[116]), .E(n743), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFX1 \block_reg[6][115]  ( .D(block_next[115]), .E(n742), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFX1 \block_reg[6][114]  ( .D(block_next[114]), .E(n744), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFX1 \block_reg[6][113]  ( .D(block_next[113]), .E(n741), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFX1 \block_reg[6][112]  ( .D(block_next[112]), .E(n242), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFX1 \block_reg[6][111]  ( .D(block_next[111]), .E(n739), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFX1 \block_reg[6][110]  ( .D(block_next[110]), .E(n740), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFX1 \block_reg[6][109]  ( .D(block_next[109]), .E(n746), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFX1 \block_reg[6][108]  ( .D(block_next[108]), .E(n746), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFX1 \block_reg[6][107]  ( .D(block_next[107]), .E(n745), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFX1 \block_reg[6][106]  ( .D(block_next[106]), .E(n743), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFX1 \block_reg[6][105]  ( .D(block_next[105]), .E(n742), .CK(clk), .Q(
        \block[6][105] ) );
  EDFFX1 \block_reg[6][104]  ( .D(block_next[104]), .E(n743), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFX1 \block_reg[6][103]  ( .D(block_next[103]), .E(n742), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFX1 \block_reg[6][102]  ( .D(block_next[102]), .E(n744), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFX1 \block_reg[6][101]  ( .D(block_next[101]), .E(n741), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFX1 \block_reg[6][100]  ( .D(block_next[100]), .E(n242), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFX1 \block_reg[6][99]  ( .D(block_next[99]), .E(n739), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFX1 \block_reg[6][98]  ( .D(block_next[98]), .E(n740), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFX1 \block_reg[6][97]  ( .D(block_next[97]), .E(n746), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFX1 \block_reg[6][96]  ( .D(block_next[96]), .E(n745), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFX1 \block_reg[6][95]  ( .D(block_next[95]), .E(n743), .CK(clk), .Q(
        \block[6][95] ) );
  EDFFX1 \block_reg[6][94]  ( .D(block_next[94]), .E(n742), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFX1 \block_reg[6][93]  ( .D(block_next[93]), .E(n744), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFX1 \block_reg[6][92]  ( .D(block_next[92]), .E(n741), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFX1 \block_reg[6][91]  ( .D(block_next[91]), .E(n746), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFX1 \block_reg[6][90]  ( .D(block_next[90]), .E(n746), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFX1 \block_reg[6][89]  ( .D(block_next[89]), .E(n746), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFX1 \block_reg[6][88]  ( .D(block_next[88]), .E(n746), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFX1 \block_reg[6][87]  ( .D(block_next[87]), .E(n746), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFX1 \block_reg[6][86]  ( .D(block_next[86]), .E(n746), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFX1 \block_reg[6][85]  ( .D(block_next[85]), .E(n746), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFX1 \block_reg[6][84]  ( .D(block_next[84]), .E(n746), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFX1 \block_reg[6][83]  ( .D(block_next[83]), .E(n746), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFX1 \block_reg[6][82]  ( .D(block_next[82]), .E(n746), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFX1 \block_reg[6][81]  ( .D(block_next[81]), .E(n746), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFX1 \block_reg[6][80]  ( .D(block_next[80]), .E(n746), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFX1 \block_reg[6][79]  ( .D(block_next[79]), .E(n746), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFX1 \block_reg[6][78]  ( .D(block_next[78]), .E(n745), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFX1 \block_reg[6][77]  ( .D(block_next[77]), .E(n745), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFX1 \block_reg[6][76]  ( .D(block_next[76]), .E(n745), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFX1 \block_reg[6][75]  ( .D(block_next[75]), .E(n745), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFX1 \block_reg[6][74]  ( .D(block_next[74]), .E(n745), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFX1 \block_reg[6][73]  ( .D(block_next[73]), .E(n745), .CK(clk), .Q(
        \block[6][73] ) );
  EDFFX1 \block_reg[6][72]  ( .D(block_next[72]), .E(n745), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFX1 \block_reg[6][71]  ( .D(block_next[71]), .E(n745), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFX1 \block_reg[6][70]  ( .D(block_next[70]), .E(n745), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFX1 \block_reg[6][69]  ( .D(block_next[69]), .E(n745), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFX1 \block_reg[6][68]  ( .D(block_next[68]), .E(n745), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFX1 \block_reg[6][67]  ( .D(block_next[67]), .E(n745), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFX1 \block_reg[6][66]  ( .D(block_next[66]), .E(n745), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFX1 \block_reg[6][65]  ( .D(block_next[65]), .E(n744), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFX1 \block_reg[6][64]  ( .D(block_next[64]), .E(n744), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFX1 \block_reg[6][63]  ( .D(block_next[63]), .E(n744), .CK(clk), .Q(
        \block[6][63] ) );
  EDFFX1 \block_reg[6][62]  ( .D(block_next[62]), .E(n744), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFX1 \block_reg[6][61]  ( .D(block_next[61]), .E(n744), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFX1 \block_reg[6][60]  ( .D(block_next[60]), .E(n744), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFX1 \block_reg[6][59]  ( .D(block_next[59]), .E(n744), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFX1 \block_reg[6][58]  ( .D(block_next[58]), .E(n744), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFX1 \block_reg[6][57]  ( .D(block_next[57]), .E(n744), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFX1 \block_reg[6][56]  ( .D(block_next[56]), .E(n744), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFX1 \block_reg[6][55]  ( .D(block_next[55]), .E(n744), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFX1 \block_reg[6][54]  ( .D(block_next[54]), .E(n744), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n744), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n743), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[6][51]  ( .D(block_next[51]), .E(n743), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFX1 \block_reg[6][50]  ( .D(block_next[50]), .E(n743), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFX1 \block_reg[6][49]  ( .D(block_next[49]), .E(n743), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFX1 \block_reg[6][48]  ( .D(block_next[48]), .E(n743), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFX1 \block_reg[6][47]  ( .D(block_next[47]), .E(n743), .CK(clk), .Q(
        \block[6][47] ) );
  EDFFX1 \block_reg[6][46]  ( .D(block_next[46]), .E(n743), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFX1 \block_reg[6][45]  ( .D(block_next[45]), .E(n743), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFX1 \block_reg[6][44]  ( .D(block_next[44]), .E(n743), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFX1 \block_reg[6][43]  ( .D(block_next[43]), .E(n743), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFX1 \block_reg[6][42]  ( .D(block_next[42]), .E(n743), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n743), .CK(clk), .Q(
        \block[6][41] ) );
  EDFFX1 \block_reg[6][40]  ( .D(block_next[40]), .E(n743), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFX1 \block_reg[6][39]  ( .D(block_next[39]), .E(n742), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n742), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n742), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n742), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n742), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFX1 \block_reg[6][34]  ( .D(block_next[34]), .E(n742), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFX1 \block_reg[6][33]  ( .D(block_next[33]), .E(n742), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n742), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[6][31]  ( .D(block_next[31]), .E(n742), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFX1 \block_reg[6][30]  ( .D(block_next[30]), .E(n742), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFX1 \block_reg[6][29]  ( .D(block_next[29]), .E(n742), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFX1 \block_reg[6][28]  ( .D(block_next[28]), .E(n742), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFX1 \block_reg[6][27]  ( .D(block_next[27]), .E(n742), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFX1 \block_reg[6][26]  ( .D(block_next[26]), .E(n741), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFX1 \block_reg[6][25]  ( .D(block_next[25]), .E(n741), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFX1 \block_reg[6][24]  ( .D(block_next[24]), .E(n741), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFX1 \block_reg[6][23]  ( .D(block_next[23]), .E(n741), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFX1 \block_reg[6][22]  ( .D(block_next[22]), .E(n741), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFX1 \block_reg[6][21]  ( .D(block_next[21]), .E(n741), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n741), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFX1 \block_reg[6][19]  ( .D(block_next[19]), .E(n741), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFX1 \block_reg[6][18]  ( .D(block_next[18]), .E(n741), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFX1 \block_reg[6][17]  ( .D(block_next[17]), .E(n741), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFX1 \block_reg[6][16]  ( .D(block_next[16]), .E(n741), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFX1 \block_reg[6][15]  ( .D(block_next[15]), .E(n741), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFX1 \block_reg[6][14]  ( .D(block_next[14]), .E(n741), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFX1 \block_reg[6][13]  ( .D(block_next[13]), .E(n740), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFX1 \block_reg[6][12]  ( .D(block_next[12]), .E(n740), .CK(clk), .Q(
        \block[6][12] ) );
  EDFFX1 \block_reg[6][11]  ( .D(block_next[11]), .E(n740), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFX1 \block_reg[6][10]  ( .D(block_next[10]), .E(n740), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFX1 \block_reg[6][9]  ( .D(block_next[9]), .E(n740), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFX1 \block_reg[6][8]  ( .D(block_next[8]), .E(n740), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFX1 \block_reg[6][7]  ( .D(block_next[7]), .E(n740), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFX1 \block_reg[6][6]  ( .D(block_next[6]), .E(n740), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFX1 \block_reg[6][5]  ( .D(block_next[5]), .E(n740), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFX1 \block_reg[6][4]  ( .D(block_next[4]), .E(n740), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFX1 \block_reg[6][3]  ( .D(block_next[3]), .E(n740), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFX1 \block_reg[6][2]  ( .D(block_next[2]), .E(n740), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFX1 \block_reg[6][1]  ( .D(block_next[1]), .E(n740), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFX1 \block_reg[6][0]  ( .D(block_next[0]), .E(n242), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFX1 \block_reg[2][127]  ( .D(block_next[127]), .E(n775), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFX1 \block_reg[2][126]  ( .D(block_next[126]), .E(n775), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFX1 \block_reg[2][125]  ( .D(block_next[125]), .E(n774), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFX1 \block_reg[2][124]  ( .D(block_next[124]), .E(n776), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFX1 \block_reg[2][123]  ( .D(block_next[123]), .E(n777), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFX1 \block_reg[2][122]  ( .D(block_next[122]), .E(n772), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFX1 \block_reg[2][121]  ( .D(block_next[121]), .E(n771), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFX1 \block_reg[2][120]  ( .D(block_next[120]), .E(n773), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFX1 \block_reg[2][119]  ( .D(block_next[119]), .E(n778), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFX1 \block_reg[2][118]  ( .D(block_next[118]), .E(n773), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFX1 \block_reg[2][117]  ( .D(block_next[117]), .E(n777), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFX1 \block_reg[2][116]  ( .D(block_next[116]), .E(n772), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFX1 \block_reg[2][115]  ( .D(block_next[115]), .E(n771), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFX1 \block_reg[2][114]  ( .D(block_next[114]), .E(n773), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFX1 \block_reg[2][113]  ( .D(block_next[113]), .E(n778), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFX1 \block_reg[2][112]  ( .D(block_next[112]), .E(n238), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFX1 \block_reg[2][111]  ( .D(block_next[111]), .E(n776), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFX1 \block_reg[2][110]  ( .D(block_next[110]), .E(n775), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFX1 \block_reg[2][109]  ( .D(block_next[109]), .E(n774), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFX1 \block_reg[2][108]  ( .D(block_next[108]), .E(n776), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFX1 \block_reg[2][107]  ( .D(block_next[107]), .E(n777), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFX1 \block_reg[2][106]  ( .D(block_next[106]), .E(n772), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFX1 \block_reg[2][105]  ( .D(block_next[105]), .E(n771), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFX1 \block_reg[2][104]  ( .D(block_next[104]), .E(n778), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFX1 \block_reg[2][103]  ( .D(block_next[103]), .E(n778), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFX1 \block_reg[2][102]  ( .D(block_next[102]), .E(n778), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFX1 \block_reg[2][101]  ( .D(block_next[101]), .E(n778), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFX1 \block_reg[2][100]  ( .D(block_next[100]), .E(n778), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFX1 \block_reg[2][99]  ( .D(block_next[99]), .E(n778), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFX1 \block_reg[2][98]  ( .D(block_next[98]), .E(n778), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFX1 \block_reg[2][97]  ( .D(block_next[97]), .E(n778), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFX1 \block_reg[2][96]  ( .D(block_next[96]), .E(n778), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFX1 \block_reg[2][95]  ( .D(block_next[95]), .E(n778), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFX1 \block_reg[2][94]  ( .D(block_next[94]), .E(n778), .CK(clk), .Q(
        \block[2][94] ) );
  EDFFX1 \block_reg[2][93]  ( .D(block_next[93]), .E(n778), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFX1 \block_reg[2][92]  ( .D(block_next[92]), .E(n778), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFX1 \block_reg[2][91]  ( .D(block_next[91]), .E(n777), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFX1 \block_reg[2][90]  ( .D(block_next[90]), .E(n777), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFX1 \block_reg[2][89]  ( .D(block_next[89]), .E(n777), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFX1 \block_reg[2][88]  ( .D(block_next[88]), .E(n777), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFX1 \block_reg[2][87]  ( .D(block_next[87]), .E(n777), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFX1 \block_reg[2][86]  ( .D(block_next[86]), .E(n777), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFX1 \block_reg[2][85]  ( .D(block_next[85]), .E(n777), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFX1 \block_reg[2][84]  ( .D(block_next[84]), .E(n777), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFX1 \block_reg[2][83]  ( .D(block_next[83]), .E(n777), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFX1 \block_reg[2][82]  ( .D(block_next[82]), .E(n777), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFX1 \block_reg[2][81]  ( .D(block_next[81]), .E(n777), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFX1 \block_reg[2][80]  ( .D(block_next[80]), .E(n777), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFX1 \block_reg[2][79]  ( .D(block_next[79]), .E(n777), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFX1 \block_reg[2][78]  ( .D(block_next[78]), .E(n772), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFX1 \block_reg[2][77]  ( .D(block_next[77]), .E(n771), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFX1 \block_reg[2][76]  ( .D(block_next[76]), .E(n773), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFX1 \block_reg[2][75]  ( .D(block_next[75]), .E(n778), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFX1 \block_reg[2][74]  ( .D(block_next[74]), .E(n238), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFX1 \block_reg[2][73]  ( .D(block_next[73]), .E(n775), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFX1 \block_reg[2][72]  ( .D(block_next[72]), .E(n774), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFX1 \block_reg[2][71]  ( .D(block_next[71]), .E(n776), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFX1 \block_reg[2][70]  ( .D(block_next[70]), .E(n777), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFX1 \block_reg[2][69]  ( .D(block_next[69]), .E(n772), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFX1 \block_reg[2][68]  ( .D(block_next[68]), .E(n771), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFX1 \block_reg[2][67]  ( .D(block_next[67]), .E(n773), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFX1 \block_reg[2][66]  ( .D(block_next[66]), .E(n778), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFX1 \block_reg[2][65]  ( .D(block_next[65]), .E(n776), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFX1 \block_reg[2][64]  ( .D(block_next[64]), .E(n776), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFX1 \block_reg[2][63]  ( .D(block_next[63]), .E(n776), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFX1 \block_reg[2][62]  ( .D(block_next[62]), .E(n776), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFX1 \block_reg[2][61]  ( .D(block_next[61]), .E(n776), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFX1 \block_reg[2][60]  ( .D(block_next[60]), .E(n776), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFX1 \block_reg[2][59]  ( .D(block_next[59]), .E(n776), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFX1 \block_reg[2][58]  ( .D(block_next[58]), .E(n776), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFX1 \block_reg[2][57]  ( .D(block_next[57]), .E(n776), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFX1 \block_reg[2][56]  ( .D(block_next[56]), .E(n776), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFX1 \block_reg[2][55]  ( .D(block_next[55]), .E(n776), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFX1 \block_reg[2][54]  ( .D(block_next[54]), .E(n776), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFX1 \block_reg[2][53]  ( .D(block_next[53]), .E(n776), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFX1 \block_reg[2][52]  ( .D(block_next[52]), .E(n775), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFX1 \block_reg[2][51]  ( .D(block_next[51]), .E(n775), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFX1 \block_reg[2][50]  ( .D(block_next[50]), .E(n775), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFX1 \block_reg[2][49]  ( .D(block_next[49]), .E(n775), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFX1 \block_reg[2][48]  ( .D(block_next[48]), .E(n775), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFX1 \block_reg[2][47]  ( .D(block_next[47]), .E(n775), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFX1 \block_reg[2][46]  ( .D(block_next[46]), .E(n775), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFX1 \block_reg[2][45]  ( .D(block_next[45]), .E(n775), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFX1 \block_reg[2][44]  ( .D(block_next[44]), .E(n775), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFX1 \block_reg[2][43]  ( .D(block_next[43]), .E(n775), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFX1 \block_reg[2][42]  ( .D(block_next[42]), .E(n775), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFX1 \block_reg[2][41]  ( .D(block_next[41]), .E(n775), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFX1 \block_reg[2][40]  ( .D(block_next[40]), .E(n775), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFX1 \block_reg[2][39]  ( .D(block_next[39]), .E(n774), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFX1 \block_reg[2][38]  ( .D(block_next[38]), .E(n774), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFX1 \block_reg[2][37]  ( .D(block_next[37]), .E(n774), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFX1 \block_reg[2][36]  ( .D(block_next[36]), .E(n774), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFX1 \block_reg[2][35]  ( .D(block_next[35]), .E(n774), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFX1 \block_reg[2][34]  ( .D(block_next[34]), .E(n774), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFX1 \block_reg[2][33]  ( .D(block_next[33]), .E(n774), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFX1 \block_reg[2][32]  ( .D(block_next[32]), .E(n774), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFX1 \block_reg[2][31]  ( .D(block_next[31]), .E(n774), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFX1 \block_reg[2][30]  ( .D(block_next[30]), .E(n774), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFX1 \block_reg[2][29]  ( .D(block_next[29]), .E(n774), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFX1 \block_reg[2][28]  ( .D(block_next[28]), .E(n774), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFX1 \block_reg[2][27]  ( .D(block_next[27]), .E(n774), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFX1 \block_reg[2][26]  ( .D(block_next[26]), .E(n238), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFX1 \block_reg[2][25]  ( .D(block_next[25]), .E(n238), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFX1 \block_reg[2][24]  ( .D(block_next[24]), .E(n238), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFX1 \block_reg[2][23]  ( .D(block_next[23]), .E(n774), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFX1 \block_reg[2][22]  ( .D(block_next[22]), .E(n775), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFX1 \block_reg[2][21]  ( .D(block_next[21]), .E(n774), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFX1 \block_reg[2][20]  ( .D(block_next[20]), .E(n776), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFX1 \block_reg[2][19]  ( .D(block_next[19]), .E(n777), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFX1 \block_reg[2][18]  ( .D(block_next[18]), .E(n772), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFX1 \block_reg[2][17]  ( .D(block_next[17]), .E(n771), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFX1 \block_reg[2][16]  ( .D(block_next[16]), .E(n773), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFX1 \block_reg[2][15]  ( .D(block_next[15]), .E(n778), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFX1 \block_reg[2][14]  ( .D(block_next[14]), .E(n778), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFX1 \block_reg[2][13]  ( .D(block_next[13]), .E(n773), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFX1 \block_reg[2][12]  ( .D(block_next[12]), .E(n773), .CK(clk), .Q(
        \block[2][12] ) );
  EDFFX1 \block_reg[2][11]  ( .D(block_next[11]), .E(n773), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFX1 \block_reg[2][10]  ( .D(block_next[10]), .E(n773), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFX1 \block_reg[2][9]  ( .D(block_next[9]), .E(n773), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFX1 \block_reg[2][8]  ( .D(block_next[8]), .E(n773), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFX1 \block_reg[2][7]  ( .D(block_next[7]), .E(n773), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFX1 \block_reg[2][6]  ( .D(block_next[6]), .E(n773), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFX1 \block_reg[2][5]  ( .D(block_next[5]), .E(n773), .CK(clk), .Q(
        \block[2][5] ) );
  EDFFX1 \block_reg[2][4]  ( .D(block_next[4]), .E(n773), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFX1 \block_reg[2][3]  ( .D(block_next[3]), .E(n773), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFX1 \block_reg[2][2]  ( .D(block_next[2]), .E(n773), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFX1 \block_reg[2][1]  ( .D(block_next[1]), .E(n773), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFX1 \block_reg[2][0]  ( .D(block_next[0]), .E(n772), .CK(clk), .Q(
        \block[2][0] ) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n494), .CK(clk), .RN(n805), .Q(blockdirty[7]), .QN(n478) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n490), .CK(clk), .RN(n804), .Q(blockdirty[3]), .QN(n474) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n493), .CK(clk), .RN(n805), .Q(blockdirty[6]), .QN(n477) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n489), .CK(clk), .RN(n804), .Q(blockdirty[2]), .QN(n473) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(n72), .E(n736), .CK(clk), .Q(
        \blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(n71), .E(n734), .CK(clk), .Q(
        \blocktag[7][23] ) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(n70), .E(n735), .CK(clk), .Q(
        \blocktag[7][22] ) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(n69), .E(n738), .CK(clk), .QN(n219) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(n68), .E(n732), .CK(clk), .QN(n227) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(n67), .E(n732), .CK(clk), .QN(n235) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(n73), .E(n733), .CK(clk), .Q(
        \blocktag[7][18] ) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(n66), .E(n737), .CK(clk), .Q(
        \blocktag[7][17] ) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(n65), .E(n731), .CK(clk), .QN(n171) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(n64), .E(n243), .CK(clk), .QN(n179) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(n63), .E(n733), .CK(clk), .Q(
        \blocktag[7][14] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(n62), .E(n243), .CK(clk), .QN(n163) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(n61), .E(n731), .CK(clk), .Q(
        \blocktag[7][12] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(n60), .E(n731), .CK(clk), .QN(n195) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(n59), .E(n731), .CK(clk), .Q(
        \blocktag[7][10] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(n58), .E(n731), .CK(clk), .QN(n187) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(n57), .E(n731), .CK(clk), .QN(n211) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(n56), .E(n731), .CK(clk), .QN(n203) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(n55), .E(n731), .CK(clk), .Q(
        \blocktag[7][6] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(n269), .E(n731), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(n54), .E(n731), .CK(clk), .QN(n143) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(n74), .E(n731), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(n268), .E(n731), .CK(clk), .Q(
        \blocktag[7][2] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(n53), .E(n731), .CK(clk), .QN(n155) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(n52), .E(n731), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(n72), .E(n764), .CK(clk), .Q(
        \blocktag[3][24] ) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(n71), .E(n764), .CK(clk), .Q(
        \blocktag[3][23] ) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(n70), .E(n764), .CK(clk), .Q(
        \blocktag[3][22] ) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(n69), .E(n764), .CK(clk), .QN(n215) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(n68), .E(n764), .CK(clk), .QN(n223) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(n67), .E(n764), .CK(clk), .QN(n231) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(n73), .E(n764), .CK(clk), .Q(
        \blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(n66), .E(n764), .CK(clk), .Q(
        \blocktag[3][17] ) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(n65), .E(n764), .CK(clk), .QN(n167) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(n64), .E(n764), .CK(clk), .QN(n175) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(n63), .E(n764), .CK(clk), .Q(
        \blocktag[3][14] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(n62), .E(n764), .CK(clk), .QN(n159) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(n61), .E(n763), .CK(clk), .Q(
        \blocktag[3][12] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(n60), .E(n763), .CK(clk), .QN(n191) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(n59), .E(n763), .CK(clk), .Q(
        \blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[3][9]  ( .D(n58), .E(n763), .CK(clk), .QN(n183) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(n57), .E(n763), .CK(clk), .QN(n207) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(n56), .E(n763), .CK(clk), .QN(n199) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(n55), .E(n763), .CK(clk), .QN(n147) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(n269), .E(n763), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(n54), .E(n763), .CK(clk), .QN(n138) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(n74), .E(n763), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(n268), .E(n763), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(n53), .E(n763), .CK(clk), .QN(n151) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(n52), .E(n763), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(n72), .E(n748), .CK(clk), .Q(
        \blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(n71), .E(n748), .CK(clk), .Q(
        \blocktag[5][23] ) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(n70), .E(n748), .CK(clk), .Q(
        \blocktag[5][22] ) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(n69), .E(n748), .CK(clk), .QN(n217) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(n68), .E(n748), .CK(clk), .QN(n225) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(n67), .E(n748), .CK(clk), .QN(n233) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(n73), .E(n748), .CK(clk), .Q(
        \blocktag[5][18] ) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(n66), .E(n748), .CK(clk), .Q(
        \blocktag[5][17] ) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(n65), .E(n748), .CK(clk), .QN(n169) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(n64), .E(n748), .CK(clk), .QN(n177) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(n63), .E(n748), .CK(clk), .Q(
        \blocktag[5][14] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(n62), .E(n748), .CK(clk), .QN(n161) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(n61), .E(n747), .CK(clk), .Q(
        \blocktag[5][12] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(n60), .E(n747), .CK(clk), .QN(n193) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(n59), .E(n747), .CK(clk), .Q(
        \blocktag[5][10] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(n58), .E(n747), .CK(clk), .QN(n185) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(n57), .E(n747), .CK(clk), .QN(n209) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(n56), .E(n747), .CK(clk), .QN(n201) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(n55), .E(n747), .CK(clk), .Q(
        \blocktag[5][6] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(n269), .E(n747), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(n54), .E(n747), .CK(clk), .QN(n141) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(n74), .E(n747), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(n268), .E(n747), .CK(clk), .Q(
        \blocktag[5][2] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(n53), .E(n747), .CK(clk), .QN(n153) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(n52), .E(n747), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(n72), .E(n780), .CK(clk), .Q(
        \blocktag[1][24] ) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(n71), .E(n780), .CK(clk), .Q(
        \blocktag[1][23] ) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(n70), .E(n780), .CK(clk), .Q(
        \blocktag[1][22] ) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(n69), .E(n780), .CK(clk), .QN(n213) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(n68), .E(n780), .CK(clk), .QN(n221) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(n67), .E(n780), .CK(clk), .QN(n229) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(n73), .E(n780), .CK(clk), .Q(
        \blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(n66), .E(n780), .CK(clk), .Q(
        \blocktag[1][17] ) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(n65), .E(n780), .CK(clk), .QN(n165) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(n64), .E(n780), .CK(clk), .QN(n173) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(n63), .E(n780), .CK(clk), .Q(
        \blocktag[1][14] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(n62), .E(n780), .CK(clk), .QN(n157) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(n61), .E(n779), .CK(clk), .Q(
        \blocktag[1][12] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(n60), .E(n779), .CK(clk), .QN(n189) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(n59), .E(n779), .CK(clk), .Q(
        \blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[1][9]  ( .D(n58), .E(n779), .CK(clk), .QN(n181) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(n57), .E(n779), .CK(clk), .QN(n205) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(n56), .E(n779), .CK(clk), .QN(n197) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(n55), .E(n779), .CK(clk), .QN(n145) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(n269), .E(n779), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(n54), .E(n779), .CK(clk), .QN(n136) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(n74), .E(n779), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(n268), .E(n779), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(n53), .E(n779), .CK(clk), .QN(n149) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(n52), .E(n779), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(n72), .E(n756), .CK(clk), .Q(
        \blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(n71), .E(n756), .CK(clk), .Q(
        \blocktag[4][23] ) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(n70), .E(n756), .CK(clk), .Q(
        \blocktag[4][22] ) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(n69), .E(n756), .CK(clk), .QN(n216) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(n68), .E(n756), .CK(clk), .QN(n224) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(n67), .E(n756), .CK(clk), .QN(n232) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(n73), .E(n756), .CK(clk), .Q(
        \blocktag[4][18] ) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(n66), .E(n756), .CK(clk), .Q(
        \blocktag[4][17] ) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(n65), .E(n756), .CK(clk), .QN(n168) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(n64), .E(n756), .CK(clk), .QN(n176) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(n63), .E(n756), .CK(clk), .Q(
        \blocktag[4][14] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(n62), .E(n756), .CK(clk), .QN(n160) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(n61), .E(n755), .CK(clk), .Q(
        \blocktag[4][12] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(n60), .E(n755), .CK(clk), .QN(n192) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(n59), .E(n755), .CK(clk), .Q(
        \blocktag[4][10] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(n58), .E(n755), .CK(clk), .QN(n184) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(n57), .E(n755), .CK(clk), .QN(n208) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(n56), .E(n755), .CK(clk), .QN(n200) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(n55), .E(n755), .CK(clk), .Q(
        \blocktag[4][6] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(n269), .E(n755), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(n54), .E(n755), .CK(clk), .QN(n139) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(n74), .E(n755), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(n268), .E(n755), .CK(clk), .Q(
        \blocktag[4][2] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(n53), .E(n755), .CK(clk), .QN(n152) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(n52), .E(n755), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(n72), .E(n788), .CK(clk), .Q(
        \blocktag[0][24] ) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(n71), .E(n788), .CK(clk), .Q(
        \blocktag[0][23] ) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(n70), .E(n788), .CK(clk), .Q(
        \blocktag[0][22] ) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(n69), .E(n788), .CK(clk), .QN(n212) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(n68), .E(n788), .CK(clk), .QN(n220) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(n67), .E(n788), .CK(clk), .QN(n228) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(n73), .E(n788), .CK(clk), .Q(
        \blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(n66), .E(n788), .CK(clk), .Q(
        \blocktag[0][17] ) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(n65), .E(n788), .CK(clk), .QN(n164) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(n64), .E(n788), .CK(clk), .QN(n172) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(n63), .E(n788), .CK(clk), .Q(
        \blocktag[0][14] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(n62), .E(n788), .CK(clk), .QN(n156) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(n61), .E(n787), .CK(clk), .Q(
        \blocktag[0][12] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(n60), .E(n787), .CK(clk), .QN(n188) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(n59), .E(n787), .CK(clk), .Q(
        \blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[0][9]  ( .D(n58), .E(n787), .CK(clk), .QN(n180) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(n57), .E(n787), .CK(clk), .QN(n204) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(n56), .E(n787), .CK(clk), .QN(n196) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(n55), .E(n787), .CK(clk), .QN(n144) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(n269), .E(n787), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(n54), .E(n787), .CK(clk), .QN(n135) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(n74), .E(n787), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(n268), .E(n787), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(n53), .E(n787), .CK(clk), .QN(n148) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(n52), .E(n787), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(n72), .E(n744), .CK(clk), .Q(
        \blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(n71), .E(n742), .CK(clk), .Q(
        \blocktag[6][23] ) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(n70), .E(n743), .CK(clk), .Q(
        \blocktag[6][22] ) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(n69), .E(n746), .CK(clk), .QN(n218) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(n68), .E(n740), .CK(clk), .QN(n226) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(n67), .E(n740), .CK(clk), .QN(n234) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(n73), .E(n741), .CK(clk), .Q(
        \blocktag[6][18] ) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(n66), .E(n745), .CK(clk), .Q(
        \blocktag[6][17] ) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(n65), .E(n739), .CK(clk), .QN(n170) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(n64), .E(n242), .CK(clk), .QN(n178) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(n63), .E(n741), .CK(clk), .Q(
        \blocktag[6][14] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(n62), .E(n242), .CK(clk), .QN(n162) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(n61), .E(n739), .CK(clk), .Q(
        \blocktag[6][12] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(n60), .E(n739), .CK(clk), .QN(n194) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(n59), .E(n739), .CK(clk), .Q(
        \blocktag[6][10] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(n58), .E(n739), .CK(clk), .QN(n186) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(n57), .E(n739), .CK(clk), .QN(n210) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(n56), .E(n739), .CK(clk), .QN(n202) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(n55), .E(n739), .CK(clk), .Q(
        \blocktag[6][6] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(n269), .E(n739), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(n54), .E(n739), .CK(clk), .QN(n142) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(n74), .E(n739), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(n268), .E(n739), .CK(clk), .Q(
        \blocktag[6][2] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(n53), .E(n739), .CK(clk), .QN(n154) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(n52), .E(n739), .CK(clk), .Q(
        \blocktag[6][0] ) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(n72), .E(n772), .CK(clk), .Q(
        \blocktag[2][24] ) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(n71), .E(n772), .CK(clk), .Q(
        \blocktag[2][23] ) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(n70), .E(n772), .CK(clk), .Q(
        \blocktag[2][22] ) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(n69), .E(n772), .CK(clk), .QN(n214) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(n68), .E(n772), .CK(clk), .QN(n222) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(n67), .E(n772), .CK(clk), .QN(n230) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(n73), .E(n772), .CK(clk), .Q(
        \blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(n66), .E(n772), .CK(clk), .Q(
        \blocktag[2][17] ) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(n65), .E(n772), .CK(clk), .QN(n166) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(n64), .E(n772), .CK(clk), .QN(n174) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(n63), .E(n772), .CK(clk), .Q(
        \blocktag[2][14] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(n62), .E(n772), .CK(clk), .QN(n158) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(n61), .E(n771), .CK(clk), .Q(
        \blocktag[2][12] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(n60), .E(n771), .CK(clk), .QN(n190) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(n59), .E(n771), .CK(clk), .Q(
        \blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[2][9]  ( .D(n58), .E(n771), .CK(clk), .QN(n182) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(n57), .E(n771), .CK(clk), .QN(n206) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(n56), .E(n771), .CK(clk), .QN(n198) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(n55), .E(n771), .CK(clk), .QN(n146) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(n269), .E(n771), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(n54), .E(n771), .CK(clk), .QN(n137) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(n74), .E(n771), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(n268), .E(n771), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(n53), .E(n771), .CK(clk), .QN(n150) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(n52), .E(n771), .CK(clk), .Q(
        \blocktag[2][0] ) );
  DFFRX1 \blockvalid_reg[7]  ( .D(n503), .CK(clk), .RN(n805), .Q(blockvalid[7]), .QN(n486) );
  DFFRX1 \blockvalid_reg[3]  ( .D(n498), .CK(clk), .RN(n804), .Q(blockvalid[3]), .QN(n482) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n500), .CK(clk), .RN(n804), .Q(blockvalid[5]), .QN(n484) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n496), .CK(clk), .RN(n804), .Q(blockvalid[1]), .QN(n480) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n492), .CK(clk), .RN(n804), .Q(blockdirty[5]), .QN(n476) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n488), .CK(clk), .RN(n804), .Q(blockdirty[1]), .QN(n472) );
  DFFRX1 \blockvalid_reg[4]  ( .D(n499), .CK(clk), .RN(n804), .Q(blockvalid[4]), .QN(n483) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n495), .CK(clk), .RN(n804), .Q(blockvalid[0]), .QN(n479) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n491), .CK(clk), .RN(n804), .Q(blockdirty[4]), .QN(n475) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n487), .CK(clk), .RN(n804), .Q(blockdirty[0]), .QN(n471) );
  DFFRX1 \blockvalid_reg[6]  ( .D(n501), .CK(clk), .RN(n805), .Q(blockvalid[6]), .QN(n485) );
  DFFRX1 \blockvalid_reg[2]  ( .D(n497), .CK(clk), .RN(n804), .Q(blockvalid[2]), .QN(n481) );
  BUFX4 U3 ( .A(n904), .Y(n693) );
  BUFX4 U4 ( .A(n696), .Y(n698) );
  BUFX4 U5 ( .A(n248), .Y(n706) );
  BUFX4 U6 ( .A(n868), .Y(n687) );
  CLKBUFX4 U7 ( .A(n248), .Y(n708) );
  OAI221X4 U8 ( .A0(n710), .A1(n959), .B0(n706), .B1(n1169), .C0(n958), .Y(
        block_next[21]) );
  CLKBUFX4 U9 ( .A(n868), .Y(n688) );
  OAI221X4 U10 ( .A0(n687), .A1(n1188), .B0(n951), .B1(n691), .C0(n842), .Y(
        block_next[121]) );
  CLKBUFX3 U11 ( .A(n868), .Y(n689) );
  BUFX4 U12 ( .A(N33), .Y(n627) );
  MXI2X2 U13 ( .A(n610), .B(n611), .S0(N33), .Y(tag[7]) );
  MXI2X2 U14 ( .A(n608), .B(n609), .S0(N33), .Y(tag[8]) );
  AOI2BB1XL U15 ( .A0N(n829), .A1N(n283), .B0(n282), .Y(n830) );
  CLKAND2X2 U16 ( .A(n282), .B(n1059), .Y(n271) );
  BUFX4 U17 ( .A(n249), .Y(n700) );
  CLKBUFX4 U18 ( .A(n904), .Y(n695) );
  BUFX20 U19 ( .A(n665), .Y(n682) );
  CLKBUFX3 U20 ( .A(n663), .Y(n665) );
  OAI221X4 U21 ( .A0(n699), .A1(n1160), .B0(n961), .B1(n703), .C0(n917), .Y(
        block_next[52]) );
  CLKBUFX4 U22 ( .A(n249), .Y(n699) );
  OAI221X4 U23 ( .A0(n700), .A1(n1100), .B0(n985), .B1(n702), .C0(n929), .Y(
        block_next[40]) );
  NAND4X2 U24 ( .A(n810), .B(n809), .C(n808), .D(n807), .Y(n828) );
  CLKXOR2X4 U25 ( .A(n1039), .B(proc_addr[13]), .Y(n809) );
  OAI221X4 U26 ( .A0(n709), .A1(n983), .B0(n707), .B1(n1109), .C0(n982), .Y(
        block_next[9]) );
  BUFX8 U27 ( .A(n248), .Y(n707) );
  OAI221X4 U28 ( .A0(n694), .A1(n1116), .B0(n979), .B1(n697), .C0(n892), .Y(
        block_next[75]) );
  CLKBUFX4 U29 ( .A(n904), .Y(n694) );
  OAI221X4 U30 ( .A0(n710), .A1(n961), .B0(n706), .B1(n1164), .C0(n960), .Y(
        block_next[20]) );
  OAI221X4 U31 ( .A0(n709), .A1(n985), .B0(n707), .B1(n1104), .C0(n984), .Y(
        block_next[8]) );
  CLKBUFX8 U32 ( .A(n664), .Y(n684) );
  BUFX8 U33 ( .A(n663), .Y(n664) );
  INVXL U34 ( .A(N32), .Y(n797) );
  INVX12 U35 ( .A(n1003), .Y(proc_stall) );
  NAND2X8 U36 ( .A(n1054), .B(n835), .Y(n1003) );
  INVX6 U37 ( .A(tag[12]), .Y(n1031) );
  MXI2X2 U38 ( .A(n600), .B(n601), .S0(n628), .Y(tag[12]) );
  NOR3X2 U39 ( .A(n265), .B(n266), .C(n267), .Y(n819) );
  XNOR2X2 U40 ( .A(n1007), .B(proc_addr[29]), .Y(n265) );
  CLKINVX8 U41 ( .A(tag[6]), .Y(n1043) );
  MXI2X4 U42 ( .A(n612), .B(n613), .S0(N33), .Y(tag[6]) );
  INVX4 U43 ( .A(tag[14]), .Y(n1027) );
  BUFX4 U44 ( .A(n616), .Y(n1) );
  MX4X1 U45 ( .A(n148), .B(n149), .C(n150), .D(n151), .S0(n684), .S1(n129), 
        .Y(n616) );
  INVX16 U46 ( .A(n128), .Y(n129) );
  CLKINVX8 U47 ( .A(tag[1]), .Y(n1049) );
  MXI2X4 U48 ( .A(n1), .B(n617), .S0(N33), .Y(tag[1]) );
  CLKINVX8 U49 ( .A(tag[23]), .Y(n1009) );
  MXI2X4 U50 ( .A(n580), .B(n581), .S0(n628), .Y(tag[23]) );
  INVX4 U51 ( .A(tag[19]), .Y(n1017) );
  INVX4 U52 ( .A(tag[20]), .Y(n1015) );
  INVX4 U53 ( .A(tag[21]), .Y(n1013) );
  CLKINVX8 U54 ( .A(tag[9]), .Y(n1037) );
  MXI2X4 U55 ( .A(n606), .B(n607), .S0(N33), .Y(tag[9]) );
  CLKINVX8 U56 ( .A(tag[22]), .Y(n1011) );
  MXI2X4 U57 ( .A(n582), .B(n583), .S0(n628), .Y(tag[22]) );
  MXI2X4 U58 ( .A(n618), .B(n619), .S0(N33), .Y(tag[0]) );
  MXI4X2 U59 ( .A(\blocktag[4][0] ), .B(\blocktag[5][0] ), .C(\blocktag[6][0] ), .D(\blocktag[7][0] ), .S0(n684), .S1(n129), .Y(n619) );
  MXI4X2 U60 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(\blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n684), .S1(n129), .Y(n618) );
  MXI2X4 U61 ( .A(n578), .B(n579), .S0(n627), .Y(tag[24]) );
  MXI4X4 U62 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n682), .S1(n654), .Y(
        n579) );
  MXI4X4 U63 ( .A(\blocktag[0][24] ), .B(\blocktag[1][24] ), .C(
        \blocktag[2][24] ), .D(\blocktag[3][24] ), .S0(n682), .S1(n654), .Y(
        n578) );
  NOR4X4 U64 ( .A(n814), .B(n813), .C(n812), .D(n811), .Y(n815) );
  CLKBUFX3 U65 ( .A(n657), .Y(n660) );
  BUFX4 U66 ( .A(N32), .Y(n657) );
  CLKBUFX3 U67 ( .A(n795), .Y(n686) );
  INVX12 U68 ( .A(n796), .Y(n795) );
  XNOR2X1 U69 ( .A(n1051), .B(proc_addr[5]), .Y(n266) );
  CLKBUFX3 U70 ( .A(n660), .Y(n631) );
  BUFX2 U71 ( .A(n686), .Y(n663) );
  BUFX16 U72 ( .A(n660), .Y(n632) );
  CLKINVX1 U73 ( .A(proc_read), .Y(n832) );
  AND2X2 U74 ( .A(n258), .B(n905), .Y(n254) );
  AND2X2 U75 ( .A(n870), .B(n869), .Y(n258) );
  NAND2X1 U76 ( .A(n832), .B(n1059), .Y(n1054) );
  CLKBUFX8 U77 ( .A(n1227), .Y(n802) );
  INVX6 U78 ( .A(N31), .Y(n796) );
  AND2X2 U79 ( .A(n1057), .B(n1058), .Y(n257) );
  MXI2X2 U80 ( .A(n604), .B(n605), .S0(N33), .Y(tag[10]) );
  MXI2X1 U81 ( .A(n596), .B(n597), .S0(n628), .Y(tag[14]) );
  MXI2X1 U82 ( .A(n594), .B(n595), .S0(n628), .Y(tag[15]) );
  MXI2X1 U83 ( .A(n592), .B(n593), .S0(n628), .Y(tag[16]) );
  MXI2X1 U84 ( .A(n590), .B(n591), .S0(n628), .Y(tag[17]) );
  MXI2X1 U85 ( .A(n584), .B(n585), .S0(n628), .Y(tag[21]) );
  MXI4X1 U86 ( .A(\blocktag[0][23] ), .B(\blocktag[1][23] ), .C(
        \blocktag[2][23] ), .D(\blocktag[3][23] ), .S0(n682), .S1(n655), .Y(
        n580) );
  MXI4X1 U87 ( .A(\blocktag[4][23] ), .B(\blocktag[5][23] ), .C(
        \blocktag[6][23] ), .D(\blocktag[7][23] ), .S0(n682), .S1(n655), .Y(
        n581) );
  INVX3 U88 ( .A(tag[0]), .Y(n1051) );
  CLKMX2X2 U89 ( .A(n274), .B(n275), .S0(N33), .Y(tag[3]) );
  CLKMX2X4 U90 ( .A(n278), .B(n279), .S0(n627), .Y(tag[5]) );
  CLKINVX1 U91 ( .A(tag[7]), .Y(n1041) );
  CLKINVX1 U92 ( .A(tag[8]), .Y(n1039) );
  INVX1 U93 ( .A(tag[11]), .Y(n1033) );
  CLKINVX1 U94 ( .A(tag[13]), .Y(n1029) );
  CLKINVX1 U95 ( .A(tag[15]), .Y(n1025) );
  INVX3 U96 ( .A(tag[16]), .Y(n1023) );
  CLKINVX1 U97 ( .A(tag[17]), .Y(n1021) );
  CLKMX2X2 U98 ( .A(n276), .B(n277), .S0(n628), .Y(tag[18]) );
  CLKINVX1 U99 ( .A(tag[24]), .Y(n1007) );
  BUFX4 U100 ( .A(n1002), .Y(n709) );
  MX4X1 U101 ( .A(\blocktag[4][3] ), .B(\blocktag[5][3] ), .C(\blocktag[6][3] ), .D(\blocktag[7][3] ), .S0(n684), .S1(n129), .Y(n275) );
  MX4X1 U102 ( .A(\blocktag[0][3] ), .B(\blocktag[1][3] ), .C(\blocktag[2][3] ), .D(\blocktag[3][3] ), .S0(n684), .S1(n129), .Y(n274) );
  OAI221X4 U103 ( .A0(n695), .A1(n1096), .B0(n987), .B1(n698), .C0(n896), .Y(
        block_next[71]) );
  OAI221X4 U104 ( .A0(n694), .A1(n1111), .B0(n981), .B1(n697), .C0(n893), .Y(
        block_next[74]) );
  OAI221X4 U105 ( .A0(n695), .A1(n1066), .B0(n999), .B1(n697), .C0(n902), .Y(
        block_next[65]) );
  OAI221X4 U106 ( .A0(n693), .A1(n1161), .B0(n961), .B1(n698), .C0(n883), .Y(
        block_next[84]) );
  OAI221X4 U107 ( .A0(n694), .A1(n1106), .B0(n983), .B1(n697), .C0(n894), .Y(
        block_next[73]) );
  OAI221X4 U108 ( .A0(n695), .A1(n1061), .B0(n1001), .B1(n697), .C0(n903), .Y(
        block_next[64]) );
  OAI221X4 U109 ( .A0(n693), .A1(n1186), .B0(n951), .B1(n697), .C0(n878), .Y(
        block_next[89]) );
  OAI221X4 U110 ( .A0(n694), .A1(n1101), .B0(n985), .B1(n697), .C0(n895), .Y(
        block_next[72]) );
  CLKINVX1 U111 ( .A(N33), .Y(n798) );
  BUFX4 U112 ( .A(N33), .Y(n628) );
  AND2X2 U113 ( .A(n283), .B(proc_stall), .Y(n270) );
  CLKBUFX3 U114 ( .A(n795), .Y(n685) );
  CLKBUFX2 U115 ( .A(n658), .Y(n629) );
  CLKBUFX3 U116 ( .A(n1218), .Y(n724) );
  CLKBUFX2 U117 ( .A(n630), .Y(n637) );
  AND2X1 U118 ( .A(n834), .B(n76), .Y(n255) );
  CLKBUFX2 U119 ( .A(n627), .Y(n620) );
  NAND2X1 U120 ( .A(mem_write), .B(blockdata[0]), .Y(n2) );
  NAND2X1 U121 ( .A(n802), .B(blockdata[8]), .Y(n3) );
  NAND2X1 U122 ( .A(n802), .B(blockdata[9]), .Y(n4) );
  NAND2X1 U123 ( .A(n802), .B(blockdata[16]), .Y(n5) );
  NAND2X1 U124 ( .A(n802), .B(blockdata[17]), .Y(n6) );
  NAND2X1 U125 ( .A(n802), .B(blockdata[18]), .Y(n7) );
  NAND2X1 U126 ( .A(n802), .B(blockdata[19]), .Y(n8) );
  NAND2X1 U127 ( .A(n802), .B(blockdata[20]), .Y(n9) );
  NAND2X1 U128 ( .A(n802), .B(blockdata[21]), .Y(n10) );
  NAND2X1 U129 ( .A(n802), .B(blockdata[22]), .Y(n11) );
  NAND2X1 U130 ( .A(n802), .B(blockdata[23]), .Y(n12) );
  NAND2X1 U131 ( .A(n802), .B(blockdata[26]), .Y(n13) );
  NAND2X1 U132 ( .A(n802), .B(blockdata[27]), .Y(n14) );
  NAND2X1 U133 ( .A(n802), .B(blockdata[28]), .Y(n15) );
  NAND2X1 U134 ( .A(n802), .B(blockdata[29]), .Y(n16) );
  NAND2X1 U135 ( .A(n802), .B(blockdata[30]), .Y(n17) );
  NAND2X1 U136 ( .A(n802), .B(blockdata[31]), .Y(n18) );
  NAND2X1 U137 ( .A(n800), .B(blockdata[94]), .Y(n19) );
  NAND2X1 U138 ( .A(n800), .B(blockdata[95]), .Y(n20) );
  NAND2X1 U139 ( .A(n800), .B(blockdata[96]), .Y(n21) );
  NAND2X1 U140 ( .A(n800), .B(blockdata[99]), .Y(n22) );
  NAND2X1 U141 ( .A(n800), .B(blockdata[100]), .Y(n23) );
  NAND2X1 U142 ( .A(n800), .B(blockdata[101]), .Y(n24) );
  NAND2X1 U143 ( .A(n800), .B(blockdata[102]), .Y(n25) );
  NAND2X1 U144 ( .A(n800), .B(blockdata[103]), .Y(n26) );
  AOI22X1 U145 ( .A0(tag[0]), .A1(mem_write), .B0(proc_addr[5]), .B1(mem_read), 
        .Y(n27) );
  AOI22X1 U146 ( .A0(tag[1]), .A1(mem_write), .B0(proc_addr[6]), .B1(mem_read), 
        .Y(n28) );
  AOI22X1 U147 ( .A0(tag[2]), .A1(mem_write), .B0(proc_addr[7]), .B1(mem_read), 
        .Y(n29) );
  AOI22X1 U148 ( .A0(tag[3]), .A1(mem_write), .B0(proc_addr[8]), .B1(mem_read), 
        .Y(n30) );
  AOI22X1 U149 ( .A0(tag[4]), .A1(mem_write), .B0(proc_addr[9]), .B1(mem_read), 
        .Y(n31) );
  AOI22X1 U150 ( .A0(tag[5]), .A1(mem_write), .B0(proc_addr[10]), .B1(mem_read), .Y(n32) );
  AOI22X1 U151 ( .A0(tag[6]), .A1(mem_write), .B0(proc_addr[11]), .B1(mem_read), .Y(n33) );
  AOI22X1 U152 ( .A0(tag[7]), .A1(mem_write), .B0(proc_addr[12]), .B1(mem_read), .Y(n34) );
  AOI22X1 U153 ( .A0(tag[8]), .A1(mem_write), .B0(proc_addr[13]), .B1(mem_read), .Y(n35) );
  AOI22X1 U154 ( .A0(tag[9]), .A1(mem_write), .B0(proc_addr[14]), .B1(mem_read), .Y(n36) );
  AOI22X1 U155 ( .A0(tag[10]), .A1(mem_write), .B0(proc_addr[15]), .B1(
        mem_read), .Y(n37) );
  AOI22X1 U156 ( .A0(tag[11]), .A1(mem_write), .B0(proc_addr[16]), .B1(
        mem_read), .Y(n38) );
  AOI22X1 U157 ( .A0(tag[12]), .A1(mem_write), .B0(proc_addr[17]), .B1(
        mem_read), .Y(n39) );
  AOI22X1 U158 ( .A0(tag[13]), .A1(mem_write), .B0(proc_addr[18]), .B1(
        mem_read), .Y(n40) );
  AOI22X1 U159 ( .A0(tag[14]), .A1(mem_write), .B0(proc_addr[19]), .B1(
        mem_read), .Y(n41) );
  AOI22X1 U160 ( .A0(tag[15]), .A1(mem_write), .B0(proc_addr[20]), .B1(
        mem_read), .Y(n42) );
  AOI22X1 U161 ( .A0(tag[16]), .A1(mem_write), .B0(proc_addr[21]), .B1(
        mem_read), .Y(n43) );
  AOI22X1 U162 ( .A0(tag[17]), .A1(mem_write), .B0(proc_addr[22]), .B1(
        mem_read), .Y(n44) );
  AOI22X1 U163 ( .A0(tag[18]), .A1(mem_write), .B0(proc_addr[23]), .B1(
        mem_read), .Y(n45) );
  AOI22X1 U164 ( .A0(tag[19]), .A1(mem_write), .B0(proc_addr[24]), .B1(
        mem_read), .Y(n46) );
  AOI22X1 U165 ( .A0(tag[20]), .A1(mem_write), .B0(proc_addr[25]), .B1(
        mem_read), .Y(n47) );
  AOI22X1 U166 ( .A0(tag[21]), .A1(mem_write), .B0(proc_addr[26]), .B1(
        mem_read), .Y(n48) );
  AOI22X1 U167 ( .A0(tag[22]), .A1(mem_write), .B0(proc_addr[27]), .B1(
        mem_read), .Y(n49) );
  AOI22X1 U168 ( .A0(tag[23]), .A1(mem_write), .B0(proc_addr[28]), .B1(
        mem_read), .Y(n50) );
  AOI22X1 U169 ( .A0(tag[24]), .A1(mem_write), .B0(proc_addr[29]), .B1(
        mem_read), .Y(n51) );
  MXI2X2 U170 ( .A(n1051), .B(n1050), .S0(n712), .Y(n52) );
  MXI2X2 U171 ( .A(n1049), .B(n1048), .S0(n712), .Y(n53) );
  MXI2X2 U172 ( .A(n1045), .B(n1044), .S0(n712), .Y(n54) );
  MXI2X2 U173 ( .A(n1043), .B(n1042), .S0(n712), .Y(n55) );
  MXI2X2 U174 ( .A(n1041), .B(n1040), .S0(n712), .Y(n56) );
  MXI2X2 U175 ( .A(n1039), .B(n1038), .S0(n712), .Y(n57) );
  MXI2X2 U176 ( .A(n1037), .B(n1036), .S0(n712), .Y(n58) );
  MXI2X2 U177 ( .A(n1035), .B(n1034), .S0(n712), .Y(n59) );
  MXI2X2 U178 ( .A(n1033), .B(n1032), .S0(n712), .Y(n60) );
  MXI2X2 U179 ( .A(n1031), .B(n1030), .S0(n712), .Y(n61) );
  MXI2X2 U180 ( .A(n1029), .B(n1028), .S0(n713), .Y(n62) );
  MXI2X2 U181 ( .A(n1027), .B(n1026), .S0(n713), .Y(n63) );
  MXI2X2 U182 ( .A(n1025), .B(n1024), .S0(n713), .Y(n64) );
  MXI2X2 U183 ( .A(n1023), .B(n1022), .S0(n713), .Y(n65) );
  MXI2X2 U184 ( .A(n1021), .B(n1020), .S0(n713), .Y(n66) );
  MXI2X2 U185 ( .A(n1017), .B(n1016), .S0(n713), .Y(n67) );
  MXI2X2 U186 ( .A(n1015), .B(n1014), .S0(n713), .Y(n68) );
  MXI2X2 U187 ( .A(n1013), .B(n1012), .S0(n713), .Y(n69) );
  MXI2X2 U188 ( .A(n1011), .B(n1010), .S0(n713), .Y(n70) );
  MXI2X2 U189 ( .A(n1009), .B(n1008), .S0(n713), .Y(n71) );
  MXI2X2 U190 ( .A(n1007), .B(n1006), .S0(n713), .Y(n72) );
  MXI2X2 U191 ( .A(n1019), .B(n1018), .S0(n713), .Y(n73) );
  MXI2X2 U192 ( .A(n1047), .B(n1046), .S0(n712), .Y(n74) );
  CLKBUFX3 U193 ( .A(n1002), .Y(n711) );
  CLKBUFX3 U194 ( .A(n1223), .Y(n728) );
  AND2X2 U195 ( .A(proc_addr[1]), .B(n1225), .Y(n75) );
  AND2X2 U196 ( .A(proc_addr[0]), .B(n1224), .Y(n76) );
  BUFX12 U197 ( .A(n800), .Y(n801) );
  AOI21X2 U198 ( .A0(mem_ready), .A1(n1054), .B0(valid), .Y(n77) );
  CLKBUFX3 U199 ( .A(n657), .Y(n659) );
  AND2X2 U200 ( .A(n802), .B(blockdata[11]), .Y(mem_wdata[11]) );
  AND2X2 U201 ( .A(n802), .B(blockdata[12]), .Y(mem_wdata[12]) );
  AND2X2 U202 ( .A(n802), .B(blockdata[13]), .Y(mem_wdata[13]) );
  AND2X2 U203 ( .A(n802), .B(blockdata[14]), .Y(mem_wdata[14]) );
  AND2X2 U204 ( .A(n800), .B(blockdata[84]), .Y(mem_wdata[84]) );
  AND2X2 U205 ( .A(n800), .B(blockdata[85]), .Y(mem_wdata[85]) );
  AND2X2 U206 ( .A(n800), .B(blockdata[86]), .Y(mem_wdata[86]) );
  AND2X2 U207 ( .A(n800), .B(blockdata[87]), .Y(mem_wdata[87]) );
  AND2X2 U208 ( .A(n800), .B(blockdata[88]), .Y(mem_wdata[88]) );
  AND2X2 U209 ( .A(n800), .B(blockdata[89]), .Y(mem_wdata[89]) );
  AND2X2 U210 ( .A(n800), .B(blockdata[90]), .Y(mem_wdata[90]) );
  AND2X2 U211 ( .A(n800), .B(blockdata[91]), .Y(mem_wdata[91]) );
  AND2X2 U212 ( .A(n800), .B(blockdata[92]), .Y(mem_wdata[92]) );
  AND2X2 U213 ( .A(n800), .B(blockdata[93]), .Y(mem_wdata[93]) );
  NAND2X1 U214 ( .A(dirty), .B(valid), .Y(n1056) );
  MXI2X1 U215 ( .A(n576), .B(n577), .S0(n627), .Y(dirty) );
  CLKAND2X12 U216 ( .A(n802), .B(blockdata[15]), .Y(mem_wdata[15]) );
  INVX12 U217 ( .A(n5), .Y(mem_wdata[16]) );
  INVX12 U218 ( .A(n6), .Y(mem_wdata[17]) );
  INVX12 U219 ( .A(n7), .Y(mem_wdata[18]) );
  INVX12 U220 ( .A(n4), .Y(mem_wdata[9]) );
  CLKAND2X12 U221 ( .A(n802), .B(blockdata[10]), .Y(mem_wdata[10]) );
  CLKAND2X12 U222 ( .A(n801), .B(blockdata[82]), .Y(mem_wdata[82]) );
  CLKAND2X12 U223 ( .A(n801), .B(blockdata[83]), .Y(mem_wdata[83]) );
  CLKAND2X12 U224 ( .A(n801), .B(blockdata[80]), .Y(mem_wdata[80]) );
  CLKAND2X12 U225 ( .A(n801), .B(blockdata[81]), .Y(mem_wdata[81]) );
  CLKAND2X12 U226 ( .A(n801), .B(blockdata[78]), .Y(mem_wdata[78]) );
  CLKAND2X12 U227 ( .A(n801), .B(blockdata[79]), .Y(mem_wdata[79]) );
  CLKAND2X12 U228 ( .A(n801), .B(blockdata[76]), .Y(mem_wdata[76]) );
  CLKAND2X12 U229 ( .A(n801), .B(blockdata[77]), .Y(mem_wdata[77]) );
  CLKAND2X12 U230 ( .A(n801), .B(blockdata[74]), .Y(mem_wdata[74]) );
  CLKAND2X12 U231 ( .A(n801), .B(blockdata[75]), .Y(mem_wdata[75]) );
  CLKAND2X12 U232 ( .A(n801), .B(blockdata[72]), .Y(mem_wdata[72]) );
  CLKAND2X12 U233 ( .A(n801), .B(blockdata[73]), .Y(mem_wdata[73]) );
  CLKAND2X12 U234 ( .A(n801), .B(blockdata[70]), .Y(mem_wdata[70]) );
  CLKAND2X12 U235 ( .A(n801), .B(blockdata[71]), .Y(mem_wdata[71]) );
  CLKAND2X12 U236 ( .A(n801), .B(blockdata[68]), .Y(mem_wdata[68]) );
  CLKAND2X12 U237 ( .A(n801), .B(blockdata[69]), .Y(mem_wdata[69]) );
  CLKAND2X12 U238 ( .A(n801), .B(blockdata[66]), .Y(mem_wdata[66]) );
  CLKAND2X12 U239 ( .A(n801), .B(blockdata[67]), .Y(mem_wdata[67]) );
  CLKAND2X12 U240 ( .A(n801), .B(blockdata[64]), .Y(mem_wdata[64]) );
  CLKAND2X12 U241 ( .A(n801), .B(blockdata[65]), .Y(mem_wdata[65]) );
  CLKAND2X12 U242 ( .A(n801), .B(blockdata[62]), .Y(mem_wdata[62]) );
  CLKAND2X12 U243 ( .A(n801), .B(blockdata[63]), .Y(mem_wdata[63]) );
  CLKAND2X12 U244 ( .A(n801), .B(blockdata[60]), .Y(mem_wdata[60]) );
  CLKAND2X12 U245 ( .A(n801), .B(blockdata[61]), .Y(mem_wdata[61]) );
  CLKAND2X12 U246 ( .A(n801), .B(blockdata[58]), .Y(mem_wdata[58]) );
  CLKAND2X12 U247 ( .A(n801), .B(blockdata[59]), .Y(mem_wdata[59]) );
  CLKAND2X12 U248 ( .A(n801), .B(blockdata[56]), .Y(mem_wdata[56]) );
  CLKAND2X12 U249 ( .A(n801), .B(blockdata[57]), .Y(mem_wdata[57]) );
  CLKAND2X12 U250 ( .A(n801), .B(blockdata[54]), .Y(mem_wdata[54]) );
  CLKAND2X12 U251 ( .A(n801), .B(blockdata[55]), .Y(mem_wdata[55]) );
  CLKAND2X12 U252 ( .A(n801), .B(blockdata[52]), .Y(mem_wdata[52]) );
  CLKAND2X12 U253 ( .A(n801), .B(blockdata[53]), .Y(mem_wdata[53]) );
  CLKAND2X12 U254 ( .A(n801), .B(blockdata[50]), .Y(mem_wdata[50]) );
  CLKAND2X12 U255 ( .A(n801), .B(blockdata[51]), .Y(mem_wdata[51]) );
  CLKAND2X12 U256 ( .A(n801), .B(blockdata[48]), .Y(mem_wdata[48]) );
  CLKAND2X12 U257 ( .A(n801), .B(blockdata[49]), .Y(mem_wdata[49]) );
  CLKAND2X12 U258 ( .A(n801), .B(blockdata[37]), .Y(mem_wdata[37]) );
  CLKAND2X12 U259 ( .A(n801), .B(blockdata[47]), .Y(mem_wdata[47]) );
  INVX12 U260 ( .A(n8), .Y(mem_wdata[19]) );
  INVX12 U261 ( .A(n9), .Y(mem_wdata[20]) );
  INVX12 U262 ( .A(n10), .Y(mem_wdata[21]) );
  INVX12 U263 ( .A(n11), .Y(mem_wdata[22]) );
  INVX12 U264 ( .A(n12), .Y(mem_wdata[23]) );
  CLKAND2X12 U265 ( .A(n802), .B(blockdata[24]), .Y(mem_wdata[24]) );
  CLKAND2X12 U266 ( .A(n802), .B(blockdata[25]), .Y(mem_wdata[25]) );
  INVX12 U267 ( .A(n19), .Y(mem_wdata[94]) );
  INVX12 U268 ( .A(n20), .Y(mem_wdata[95]) );
  INVX12 U269 ( .A(n21), .Y(mem_wdata[96]) );
  CLKAND2X12 U270 ( .A(n800), .B(blockdata[97]), .Y(mem_wdata[97]) );
  CLKAND2X12 U271 ( .A(n800), .B(blockdata[98]), .Y(mem_wdata[98]) );
  CLKAND2X12 U272 ( .A(mem_write), .B(blockdata[122]), .Y(mem_wdata[122]) );
  CLKAND2X12 U273 ( .A(mem_write), .B(blockdata[123]), .Y(mem_wdata[123]) );
  CLKAND2X12 U274 ( .A(mem_write), .B(blockdata[124]), .Y(mem_wdata[124]) );
  CLKAND2X12 U275 ( .A(mem_write), .B(blockdata[125]), .Y(mem_wdata[125]) );
  CLKBUFX6 U276 ( .A(n1227), .Y(mem_write) );
  INVX12 U277 ( .A(n27), .Y(mem_addr[3]) );
  INVX12 U278 ( .A(n28), .Y(mem_addr[4]) );
  INVX12 U279 ( .A(n29), .Y(mem_addr[5]) );
  INVX12 U280 ( .A(n30), .Y(mem_addr[6]) );
  INVX12 U281 ( .A(n31), .Y(mem_addr[7]) );
  INVX12 U282 ( .A(n32), .Y(mem_addr[8]) );
  INVX12 U283 ( .A(n33), .Y(mem_addr[9]) );
  INVX12 U284 ( .A(n34), .Y(mem_addr[10]) );
  INVX12 U285 ( .A(n35), .Y(mem_addr[11]) );
  INVX12 U286 ( .A(n36), .Y(mem_addr[12]) );
  INVX12 U287 ( .A(n37), .Y(mem_addr[13]) );
  INVX12 U288 ( .A(n38), .Y(mem_addr[14]) );
  INVX12 U289 ( .A(n39), .Y(mem_addr[15]) );
  INVX12 U290 ( .A(n40), .Y(mem_addr[16]) );
  INVX12 U291 ( .A(n41), .Y(mem_addr[17]) );
  INVX12 U292 ( .A(n42), .Y(mem_addr[18]) );
  INVX12 U293 ( .A(n43), .Y(mem_addr[19]) );
  INVX12 U294 ( .A(n44), .Y(mem_addr[20]) );
  INVX12 U295 ( .A(n45), .Y(mem_addr[21]) );
  INVX12 U296 ( .A(n46), .Y(mem_addr[22]) );
  INVX12 U297 ( .A(n47), .Y(mem_addr[23]) );
  INVX12 U298 ( .A(n48), .Y(mem_addr[24]) );
  INVX12 U299 ( .A(n49), .Y(mem_addr[25]) );
  INVX12 U300 ( .A(n50), .Y(mem_addr[26]) );
  INVX12 U301 ( .A(n51), .Y(mem_addr[27]) );
  INVX12 U302 ( .A(n2), .Y(mem_wdata[0]) );
  INVX12 U303 ( .A(n3), .Y(mem_wdata[8]) );
  INVX12 U304 ( .A(n13), .Y(mem_wdata[26]) );
  INVX12 U305 ( .A(n14), .Y(mem_wdata[27]) );
  INVX12 U306 ( .A(n15), .Y(mem_wdata[28]) );
  INVX12 U307 ( .A(n16), .Y(mem_wdata[29]) );
  INVX12 U308 ( .A(n17), .Y(mem_wdata[30]) );
  INVX12 U309 ( .A(n18), .Y(mem_wdata[31]) );
  CLKAND2X12 U310 ( .A(n802), .B(blockdata[32]), .Y(mem_wdata[32]) );
  CLKAND2X12 U311 ( .A(n802), .B(blockdata[33]), .Y(mem_wdata[33]) );
  CLKAND2X12 U312 ( .A(n802), .B(blockdata[34]), .Y(mem_wdata[34]) );
  CLKAND2X12 U313 ( .A(n802), .B(blockdata[35]), .Y(mem_wdata[35]) );
  CLKAND2X12 U314 ( .A(n802), .B(blockdata[36]), .Y(mem_wdata[36]) );
  CLKAND2X12 U315 ( .A(n802), .B(blockdata[38]), .Y(mem_wdata[38]) );
  CLKAND2X12 U316 ( .A(n802), .B(blockdata[39]), .Y(mem_wdata[39]) );
  CLKAND2X12 U317 ( .A(n802), .B(blockdata[40]), .Y(mem_wdata[40]) );
  CLKAND2X12 U318 ( .A(n802), .B(blockdata[41]), .Y(mem_wdata[41]) );
  CLKAND2X12 U319 ( .A(n802), .B(blockdata[42]), .Y(mem_wdata[42]) );
  CLKAND2X12 U320 ( .A(n802), .B(blockdata[43]), .Y(mem_wdata[43]) );
  CLKAND2X12 U321 ( .A(n802), .B(blockdata[44]), .Y(mem_wdata[44]) );
  CLKAND2X12 U322 ( .A(n802), .B(blockdata[45]), .Y(mem_wdata[45]) );
  INVX12 U323 ( .A(n22), .Y(mem_wdata[99]) );
  INVX12 U324 ( .A(n23), .Y(mem_wdata[100]) );
  INVX12 U325 ( .A(n24), .Y(mem_wdata[101]) );
  INVX12 U326 ( .A(n25), .Y(mem_wdata[102]) );
  INVX12 U327 ( .A(n26), .Y(mem_wdata[103]) );
  CLKAND2X12 U328 ( .A(n800), .B(blockdata[104]), .Y(mem_wdata[104]) );
  CLKAND2X12 U329 ( .A(n800), .B(blockdata[105]), .Y(mem_wdata[105]) );
  CLKAND2X12 U330 ( .A(n800), .B(blockdata[106]), .Y(mem_wdata[106]) );
  CLKAND2X12 U331 ( .A(n800), .B(blockdata[107]), .Y(mem_wdata[107]) );
  CLKAND2X12 U332 ( .A(n800), .B(blockdata[108]), .Y(mem_wdata[108]) );
  CLKAND2X12 U333 ( .A(n800), .B(blockdata[109]), .Y(mem_wdata[109]) );
  CLKAND2X12 U334 ( .A(n800), .B(blockdata[110]), .Y(mem_wdata[110]) );
  CLKAND2X12 U335 ( .A(n800), .B(blockdata[111]), .Y(mem_wdata[111]) );
  CLKAND2X12 U336 ( .A(n800), .B(blockdata[112]), .Y(mem_wdata[112]) );
  CLKAND2X12 U337 ( .A(n800), .B(blockdata[113]), .Y(mem_wdata[113]) );
  CLKAND2X12 U338 ( .A(n800), .B(blockdata[114]), .Y(mem_wdata[114]) );
  CLKAND2X12 U339 ( .A(n800), .B(blockdata[115]), .Y(mem_wdata[115]) );
  CLKAND2X12 U340 ( .A(n800), .B(blockdata[116]), .Y(mem_wdata[116]) );
  CLKAND2X12 U341 ( .A(n800), .B(blockdata[117]), .Y(mem_wdata[117]) );
  CLKAND2X12 U342 ( .A(n800), .B(blockdata[118]), .Y(mem_wdata[118]) );
  CLKAND2X12 U343 ( .A(n800), .B(blockdata[119]), .Y(mem_wdata[119]) );
  CLKAND2X12 U344 ( .A(n800), .B(blockdata[120]), .Y(mem_wdata[120]) );
  CLKAND2X12 U345 ( .A(n800), .B(blockdata[121]), .Y(mem_wdata[121]) );
  CLKAND2X12 U346 ( .A(n802), .B(blockdata[46]), .Y(mem_wdata[46]) );
  NAND4X2 U347 ( .A(n818), .B(n817), .C(n816), .D(n815), .Y(n827) );
  NAND4X2 U348 ( .A(n870), .B(n905), .C(n704), .D(n709), .Y(n833) );
  OAI221X4 U349 ( .A0(n688), .A1(n1103), .B0(n985), .B1(n692), .C0(n859), .Y(
        block_next[104]) );
  OAI221X4 U350 ( .A0(n687), .A1(n1183), .B0(n953), .B1(n691), .C0(n843), .Y(
        block_next[120]) );
  CLKAND2X12 U351 ( .A(mem_write), .B(blockdata[126]), .Y(mem_wdata[126]) );
  MX4X1 U352 ( .A(n164), .B(n165), .C(n166), .D(n167), .S0(n685), .S1(n658), 
        .Y(n592) );
  CLKBUFX3 U353 ( .A(n657), .Y(n658) );
  AND2XL U354 ( .A(mem_write), .B(blockdata[127]), .Y(mem_wdata[127]) );
  AND4X4 U355 ( .A(n822), .B(n821), .C(n820), .D(n819), .Y(n133) );
  BUFX6 U356 ( .A(n660), .Y(n630) );
  XOR2X4 U357 ( .A(proc_addr[8]), .B(tag[3]), .Y(n812) );
  MXI2X2 U358 ( .A(n614), .B(n615), .S0(N33), .Y(tag[4]) );
  BUFX12 U359 ( .A(n664), .Y(n683) );
  MX4X1 U360 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n682), .S1(n655), 
        .Y(n585) );
  MX4X1 U361 ( .A(n232), .B(n233), .C(n234), .D(n235), .S0(n682), .S1(n655), 
        .Y(n589) );
  MX4X1 U362 ( .A(n224), .B(n225), .C(n226), .D(n227), .S0(n682), .S1(n655), 
        .Y(n587) );
  BUFX16 U363 ( .A(n634), .Y(n655) );
  CLKBUFX3 U364 ( .A(n632), .Y(n633) );
  CLKINVX6 U365 ( .A(n656), .Y(n128) );
  CLKBUFX2 U366 ( .A(n633), .Y(n656) );
  XOR2X4 U367 ( .A(proc_addr[23]), .B(tag[18]), .Y(n811) );
  MXI2X1 U368 ( .A(n560), .B(n561), .S0(n627), .Y(blockdata[7]) );
  MXI2X1 U369 ( .A(n562), .B(n563), .S0(n627), .Y(blockdata[6]) );
  MXI2X1 U370 ( .A(n564), .B(n565), .S0(n627), .Y(blockdata[5]) );
  CLKAND2X12 U371 ( .A(n801), .B(blockdata[7]), .Y(mem_wdata[7]) );
  MXI2X1 U372 ( .A(n566), .B(n567), .S0(n627), .Y(blockdata[4]) );
  CLKAND2X12 U373 ( .A(n801), .B(blockdata[6]), .Y(mem_wdata[6]) );
  MXI2X1 U374 ( .A(n568), .B(n569), .S0(n627), .Y(blockdata[3]) );
  CLKAND2X12 U375 ( .A(n801), .B(blockdata[5]), .Y(mem_wdata[5]) );
  MXI2X1 U376 ( .A(n570), .B(n571), .S0(n627), .Y(blockdata[2]) );
  CLKAND2X12 U377 ( .A(n801), .B(blockdata[4]), .Y(mem_wdata[4]) );
  MXI2X1 U378 ( .A(n572), .B(n573), .S0(n627), .Y(blockdata[1]) );
  BUFX12 U379 ( .A(n1228), .Y(mem_addr[2]) );
  NOR2XL U380 ( .A(n257), .B(n798), .Y(n1228) );
  CLKAND2X12 U381 ( .A(n801), .B(blockdata[3]), .Y(mem_wdata[3]) );
  BUFX12 U382 ( .A(n1229), .Y(mem_addr[1]) );
  NOR2XL U383 ( .A(n257), .B(n797), .Y(n1229) );
  OR2X1 U384 ( .A(n257), .B(n796), .Y(n1230) );
  INVX12 U385 ( .A(n1230), .Y(mem_addr[0]) );
  CLKAND2X12 U386 ( .A(n801), .B(blockdata[2]), .Y(mem_wdata[2]) );
  CLKAND2X12 U387 ( .A(n801), .B(blockdata[1]), .Y(mem_wdata[1]) );
  XOR2XL U388 ( .A(n1025), .B(proc_addr[20]), .Y(n826) );
  CLKBUFX8 U389 ( .A(n1227), .Y(n800) );
  CLKBUFX2 U390 ( .A(n270), .Y(n720) );
  NAND3BX1 U391 ( .AN(n705), .B(n258), .C(n711), .Y(n871) );
  NAND2X1 U392 ( .A(mem_rdata[0]), .B(n713), .Y(n1000) );
  AND2X2 U393 ( .A(n254), .B(n704), .Y(n248) );
  AND2X2 U394 ( .A(n254), .B(n711), .Y(n249) );
  XOR2X1 U395 ( .A(n1013), .B(proc_addr[26]), .Y(n820) );
  XOR2X1 U396 ( .A(n1049), .B(proc_addr[6]), .Y(n824) );
  XOR2X1 U397 ( .A(n1029), .B(proc_addr[18]), .Y(n825) );
  XOR2X1 U398 ( .A(n1017), .B(proc_addr[24]), .Y(n821) );
  XOR2X1 U399 ( .A(n1015), .B(proc_addr[25]), .Y(n822) );
  XOR2X1 U400 ( .A(n1041), .B(proc_addr[12]), .Y(n810) );
  XOR2X1 U401 ( .A(n1033), .B(proc_addr[16]), .Y(n808) );
  XNOR2X1 U402 ( .A(n1009), .B(proc_addr[28]), .Y(n267) );
  XNOR2X1 U403 ( .A(n1011), .B(proc_addr[27]), .Y(n261) );
  XNOR2X1 U404 ( .A(n1035), .B(proc_addr[15]), .Y(n259) );
  XOR2X4 U405 ( .A(n1043), .B(proc_addr[11]), .Y(n818) );
  XOR2X4 U406 ( .A(n1045), .B(proc_addr[9]), .Y(n817) );
  XOR2X4 U407 ( .A(n1037), .B(proc_addr[14]), .Y(n816) );
  MXI4XL U408 ( .A(\blocktag[4][6] ), .B(\blocktag[5][6] ), .C(
        \blocktag[6][6] ), .D(\blocktag[7][6] ), .S0(n683), .S1(n636), .Y(n613) );
  CLKMX2X2 U409 ( .A(n272), .B(n273), .S0(n627), .Y(valid) );
  XOR2X4 U410 ( .A(proc_addr[10]), .B(tag[5]), .Y(n813) );
  XOR2X4 U411 ( .A(proc_addr[7]), .B(tag[2]), .Y(n814) );
  BUFX12 U412 ( .A(n635), .Y(n654) );
  CLKBUFX2 U413 ( .A(n635), .Y(n653) );
  CLKBUFX2 U414 ( .A(n686), .Y(n662) );
  CLKBUFX2 U415 ( .A(n686), .Y(n661) );
  NOR2XL U416 ( .A(n628), .B(N32), .Y(n470) );
  CLKBUFX2 U417 ( .A(n869), .Y(n690) );
  CLKBUFX2 U418 ( .A(n905), .Y(n696) );
  NOR2XL U419 ( .A(n797), .B(n628), .Y(n469) );
  NOR2XL U420 ( .A(n798), .B(N32), .Y(n468) );
  INVX3 U421 ( .A(tag[4]), .Y(n1045) );
  NAND2X4 U422 ( .A(valid), .B(n829), .Y(n835) );
  NAND4BBX4 U423 ( .AN(n828), .BN(n827), .C(n133), .D(n134), .Y(n1055) );
  AND4X4 U424 ( .A(n826), .B(n825), .C(n824), .D(n823), .Y(n134) );
  CLKINVX6 U425 ( .A(n1004), .Y(n834) );
  NAND4BXL U426 ( .AN(n1056), .B(n1055), .C(n1054), .D(n1053), .Y(n1057) );
  INVXL U427 ( .A(proc_addr[5]), .Y(n1050) );
  INVXL U428 ( .A(proc_addr[9]), .Y(n1044) );
  INVXL U429 ( .A(proc_addr[14]), .Y(n1036) );
  INVXL U430 ( .A(proc_addr[15]), .Y(n1034) );
  INVXL U431 ( .A(proc_addr[16]), .Y(n1032) );
  INVXL U432 ( .A(proc_addr[17]), .Y(n1030) );
  INVXL U433 ( .A(proc_addr[18]), .Y(n1028) );
  INVXL U434 ( .A(proc_addr[19]), .Y(n1026) );
  INVXL U435 ( .A(proc_addr[21]), .Y(n1022) );
  INVXL U436 ( .A(proc_addr[22]), .Y(n1020) );
  INVXL U437 ( .A(proc_addr[24]), .Y(n1016) );
  INVXL U438 ( .A(proc_addr[25]), .Y(n1014) );
  INVXL U439 ( .A(proc_addr[27]), .Y(n1010) );
  INVXL U440 ( .A(proc_addr[28]), .Y(n1008) );
  INVXL U441 ( .A(proc_addr[29]), .Y(n1006) );
  MX4XL U442 ( .A(n135), .B(n136), .C(n137), .D(n138), .S0(n684), .S1(n129), 
        .Y(n614) );
  MX4XL U443 ( .A(n139), .B(n141), .C(n142), .D(n143), .S0(n684), .S1(n129), 
        .Y(n615) );
  MX4XL U444 ( .A(n144), .B(n145), .C(n146), .D(n147), .S0(n684), .S1(n629), 
        .Y(n612) );
  MX4XL U445 ( .A(n152), .B(n153), .C(n154), .D(n155), .S0(n684), .S1(n129), 
        .Y(n617) );
  MX4XL U446 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n661), .S1(n658), 
        .Y(n598) );
  MX4XL U447 ( .A(n160), .B(n161), .C(n162), .D(n163), .S0(n685), .S1(n630), 
        .Y(n599) );
  MX4XL U448 ( .A(n168), .B(n169), .C(n170), .D(n171), .S0(n685), .S1(n658), 
        .Y(n593) );
  MX4XL U449 ( .A(n172), .B(n173), .C(n174), .D(n175), .S0(n685), .S1(n659), 
        .Y(n594) );
  MX4XL U450 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n661), .S1(n659), 
        .Y(n595) );
  MX4XL U451 ( .A(n180), .B(n181), .C(n182), .D(n183), .S0(n683), .S1(n636), 
        .Y(n606) );
  MX4XL U452 ( .A(n184), .B(n185), .C(n186), .D(n187), .S0(n683), .S1(n636), 
        .Y(n607) );
  MX4XL U453 ( .A(n188), .B(n189), .C(n190), .D(n191), .S0(n683), .S1(n630), 
        .Y(n602) );
  MX4XL U454 ( .A(n192), .B(n193), .C(n194), .D(n195), .S0(n683), .S1(n659), 
        .Y(n603) );
  MX4XL U455 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n683), .S1(n658), 
        .Y(n610) );
  MX4XL U456 ( .A(n200), .B(n201), .C(n202), .D(n203), .S0(n683), .S1(n630), 
        .Y(n611) );
  MX4XL U457 ( .A(n204), .B(n205), .C(n206), .D(n207), .S0(n683), .S1(n630), 
        .Y(n608) );
  MX4XL U458 ( .A(n208), .B(n209), .C(n210), .D(n211), .S0(n683), .S1(n630), 
        .Y(n609) );
  MX4XL U459 ( .A(n212), .B(n213), .C(n214), .D(n215), .S0(n682), .S1(n655), 
        .Y(n584) );
  MX4XL U460 ( .A(n220), .B(n221), .C(n222), .D(n223), .S0(n682), .S1(n655), 
        .Y(n586) );
  MX4XL U461 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n666), .S1(n654), .Y(n272) );
  MX4XL U462 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n666), .S1(n654), .Y(n273) );
  MX4XL U463 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n685), .S1(n655), .Y(
        n276) );
  MX4XL U464 ( .A(\blocktag[4][18] ), .B(\blocktag[5][18] ), .C(
        \blocktag[6][18] ), .D(\blocktag[7][18] ), .S0(n685), .S1(n655), .Y(
        n277) );
  CLKMX2X4 U465 ( .A(n280), .B(n281), .S0(N33), .Y(tag[2]) );
  MX4XL U466 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(\blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n684), .S1(n129), .Y(n280) );
  MX4XL U467 ( .A(\blocktag[4][2] ), .B(\blocktag[5][2] ), .C(\blocktag[6][2] ), .D(\blocktag[7][2] ), .S0(n684), .S1(n129), .Y(n281) );
  MX4XL U468 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(\blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n684), .S1(n129), .Y(n278) );
  MX4XL U469 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(\blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n684), .S1(n129), .Y(n279) );
  MX4XL U470 ( .A(n228), .B(n229), .C(n230), .D(n231), .S0(n685), .S1(n655), 
        .Y(n588) );
  MXI4XL U471 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n682), .S1(n654), .Y(n577) );
  MXI4XL U472 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n682), .S1(n654), .Y(n576) );
  NOR2BXL U473 ( .AN(proc_read), .B(n835), .Y(n282) );
  NAND3BXL U474 ( .AN(mem_ready), .B(proc_stall), .C(n1056), .Y(n1058) );
  INVXL U475 ( .A(tag[3]), .Y(n1047) );
  INVXL U476 ( .A(tag[18]), .Y(n1019) );
  MXI2XL U477 ( .A(n574), .B(n575), .S0(n627), .Y(blockdata[0]) );
  MXI4XL U478 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n666), .S1(n654), .Y(n575) );
  MXI4XL U479 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n666), .S1(n654), .Y(n574) );
  MXI4XL U480 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n666), .S1(n654), .Y(n573) );
  MXI4XL U481 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n682), .S1(n654), .Y(n572) );
  MXI4XL U482 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n666), .S1(n654), .Y(n571) );
  MXI4XL U483 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n665), .S1(n654), .Y(n570) );
  MXI4XL U484 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n666), .S1(n653), .Y(n569) );
  MXI4XL U485 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n682), .S1(n653), .Y(n568) );
  MXI4XL U486 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n666), .S1(n653), .Y(n567) );
  MXI4XL U487 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n682), .S1(n653), .Y(n566) );
  MXI4XL U488 ( .A(\block[0][5] ), .B(\block[1][5] ), .C(\block[2][5] ), .D(
        \block[3][5] ), .S0(n682), .S1(n653), .Y(n564) );
  MXI2XL U489 ( .A(n558), .B(n559), .S0(n627), .Y(blockdata[8]) );
  AND2XL U490 ( .A(mem_ready), .B(n1056), .Y(n283) );
  CLKBUFX3 U491 ( .A(n637), .Y(n650) );
  CLKBUFX3 U492 ( .A(n637), .Y(n649) );
  CLKBUFX3 U493 ( .A(n637), .Y(n644) );
  CLKBUFX3 U494 ( .A(n637), .Y(n648) );
  CLKBUFX3 U495 ( .A(n637), .Y(n643) );
  CLKBUFX3 U496 ( .A(n637), .Y(n647) );
  CLKBUFX3 U497 ( .A(n637), .Y(n642) );
  CLKBUFX3 U498 ( .A(n637), .Y(n646) );
  CLKBUFX3 U499 ( .A(n637), .Y(n641) );
  CLKBUFX3 U500 ( .A(n637), .Y(n645) );
  CLKBUFX3 U501 ( .A(n637), .Y(n640) );
  CLKBUFX3 U502 ( .A(n653), .Y(n639) );
  CLKBUFX3 U503 ( .A(n636), .Y(n652) );
  CLKBUFX3 U504 ( .A(n636), .Y(n651) );
  CLKBUFX3 U505 ( .A(n632), .Y(n634) );
  CLKBUFX3 U506 ( .A(n631), .Y(n635) );
  CLKBUFX3 U507 ( .A(n666), .Y(n675) );
  CLKBUFX3 U508 ( .A(n666), .Y(n679) );
  CLKBUFX3 U509 ( .A(n666), .Y(n674) );
  CLKBUFX3 U510 ( .A(n666), .Y(n678) );
  CLKBUFX3 U511 ( .A(n666), .Y(n673) );
  CLKBUFX3 U512 ( .A(n666), .Y(n677) );
  CLKBUFX3 U513 ( .A(n666), .Y(n672) );
  CLKBUFX3 U514 ( .A(n684), .Y(n676) );
  CLKBUFX3 U515 ( .A(n666), .Y(n671) );
  CLKBUFX3 U516 ( .A(n684), .Y(n670) );
  CLKBUFX3 U517 ( .A(n666), .Y(n669) );
  CLKBUFX3 U518 ( .A(n684), .Y(n681) );
  CLKBUFX3 U519 ( .A(n666), .Y(n668) );
  CLKBUFX3 U520 ( .A(n684), .Y(n680) );
  CLKBUFX3 U521 ( .A(n662), .Y(n667) );
  CLKBUFX3 U522 ( .A(n620), .Y(n625) );
  CLKBUFX3 U523 ( .A(n620), .Y(n624) );
  CLKBUFX3 U524 ( .A(n620), .Y(n623) );
  CLKBUFX3 U525 ( .A(n624), .Y(n622) );
  CLKBUFX3 U526 ( .A(n623), .Y(n621) );
  CLKBUFX3 U527 ( .A(n625), .Y(n626) );
  CLKBUFX3 U528 ( .A(n631), .Y(n636) );
  CLKBUFX3 U529 ( .A(n236), .Y(n789) );
  CLKBUFX3 U530 ( .A(n236), .Y(n790) );
  CLKBUFX3 U531 ( .A(n236), .Y(n791) );
  CLKBUFX3 U532 ( .A(n236), .Y(n792) );
  CLKBUFX3 U533 ( .A(n236), .Y(n793) );
  CLKBUFX3 U534 ( .A(n236), .Y(n794) );
  CLKBUFX3 U535 ( .A(n237), .Y(n781) );
  CLKBUFX3 U536 ( .A(n237), .Y(n782) );
  CLKBUFX3 U537 ( .A(n237), .Y(n783) );
  CLKBUFX3 U538 ( .A(n237), .Y(n784) );
  CLKBUFX3 U539 ( .A(n237), .Y(n785) );
  CLKBUFX3 U540 ( .A(n237), .Y(n786) );
  CLKBUFX3 U541 ( .A(n238), .Y(n773) );
  CLKBUFX3 U542 ( .A(n238), .Y(n774) );
  CLKBUFX3 U543 ( .A(n238), .Y(n775) );
  CLKBUFX3 U544 ( .A(n238), .Y(n776) );
  CLKBUFX3 U545 ( .A(n238), .Y(n777) );
  CLKBUFX3 U546 ( .A(n238), .Y(n778) );
  CLKBUFX3 U547 ( .A(n239), .Y(n765) );
  CLKBUFX3 U548 ( .A(n239), .Y(n766) );
  CLKBUFX3 U549 ( .A(n239), .Y(n767) );
  CLKBUFX3 U550 ( .A(n239), .Y(n768) );
  CLKBUFX3 U551 ( .A(n239), .Y(n769) );
  CLKBUFX3 U552 ( .A(n239), .Y(n770) );
  CLKBUFX3 U553 ( .A(n240), .Y(n757) );
  CLKBUFX3 U554 ( .A(n240), .Y(n758) );
  CLKBUFX3 U555 ( .A(n240), .Y(n759) );
  CLKBUFX3 U556 ( .A(n240), .Y(n760) );
  CLKBUFX3 U557 ( .A(n240), .Y(n761) );
  CLKBUFX3 U558 ( .A(n240), .Y(n762) );
  CLKBUFX3 U559 ( .A(n241), .Y(n749) );
  CLKBUFX3 U560 ( .A(n241), .Y(n750) );
  CLKBUFX3 U561 ( .A(n241), .Y(n751) );
  CLKBUFX3 U562 ( .A(n241), .Y(n752) );
  CLKBUFX3 U563 ( .A(n241), .Y(n753) );
  CLKBUFX3 U564 ( .A(n241), .Y(n754) );
  CLKBUFX3 U565 ( .A(n242), .Y(n740) );
  CLKBUFX3 U566 ( .A(n242), .Y(n741) );
  CLKBUFX3 U567 ( .A(n242), .Y(n742) );
  CLKBUFX3 U568 ( .A(n242), .Y(n743) );
  CLKBUFX3 U569 ( .A(n242), .Y(n744) );
  CLKBUFX3 U570 ( .A(n242), .Y(n745) );
  CLKBUFX3 U571 ( .A(n242), .Y(n746) );
  CLKBUFX3 U572 ( .A(n243), .Y(n732) );
  CLKBUFX3 U573 ( .A(n243), .Y(n733) );
  CLKBUFX3 U574 ( .A(n243), .Y(n734) );
  CLKBUFX3 U575 ( .A(n243), .Y(n735) );
  CLKBUFX3 U576 ( .A(n243), .Y(n736) );
  CLKBUFX3 U577 ( .A(n243), .Y(n737) );
  CLKBUFX3 U578 ( .A(n243), .Y(n738) );
  CLKBUFX3 U579 ( .A(n236), .Y(n787) );
  CLKBUFX3 U580 ( .A(n236), .Y(n788) );
  CLKBUFX3 U581 ( .A(n237), .Y(n779) );
  CLKBUFX3 U582 ( .A(n237), .Y(n780) );
  CLKBUFX3 U583 ( .A(n238), .Y(n771) );
  CLKBUFX3 U584 ( .A(n238), .Y(n772) );
  CLKBUFX3 U585 ( .A(n239), .Y(n763) );
  CLKBUFX3 U586 ( .A(n239), .Y(n764) );
  CLKBUFX3 U587 ( .A(n240), .Y(n755) );
  CLKBUFX3 U588 ( .A(n240), .Y(n756) );
  CLKBUFX3 U589 ( .A(n241), .Y(n747) );
  CLKBUFX3 U590 ( .A(n241), .Y(n748) );
  CLKBUFX3 U591 ( .A(n242), .Y(n739) );
  CLKBUFX3 U592 ( .A(n243), .Y(n731) );
  CLKBUFX3 U593 ( .A(n662), .Y(n666) );
  CLKBUFX3 U594 ( .A(n637), .Y(n638) );
  CLKBUFX3 U595 ( .A(n711), .Y(n710) );
  CLKBUFX3 U596 ( .A(n696), .Y(n697) );
  CLKBUFX3 U597 ( .A(n690), .Y(n692) );
  CLKBUFX3 U598 ( .A(n690), .Y(n691) );
  CLKBUFX3 U599 ( .A(n249), .Y(n701) );
  INVX3 U600 ( .A(n255), .Y(n704) );
  CLKBUFX3 U601 ( .A(n270), .Y(n712) );
  CLKBUFX3 U602 ( .A(n270), .Y(n713) );
  CLKBUFX3 U603 ( .A(n270), .Y(n714) );
  CLKBUFX3 U604 ( .A(n270), .Y(n715) );
  CLKBUFX3 U605 ( .A(n270), .Y(n716) );
  CLKBUFX3 U606 ( .A(n270), .Y(n717) );
  CLKBUFX3 U607 ( .A(n270), .Y(n718) );
  CLKBUFX3 U608 ( .A(n270), .Y(n719) );
  CLKBUFX3 U609 ( .A(n1221), .Y(n726) );
  CLKBUFX3 U610 ( .A(n1221), .Y(n727) );
  CLKBUFX3 U611 ( .A(n728), .Y(n729) );
  CLKBUFX3 U612 ( .A(n728), .Y(n730) );
  CLKBUFX3 U613 ( .A(n1218), .Y(n725) );
  CLKBUFX3 U614 ( .A(n1216), .Y(n722) );
  CLKBUFX3 U615 ( .A(n1216), .Y(n723) );
  AND2X2 U616 ( .A(n250), .B(n805), .Y(n236) );
  AND2X2 U617 ( .A(n244), .B(n805), .Y(n237) );
  AND2X2 U618 ( .A(n251), .B(n805), .Y(n238) );
  AND2X2 U619 ( .A(n245), .B(n805), .Y(n239) );
  AND2X2 U620 ( .A(n253), .B(n805), .Y(n240) );
  AND2X2 U621 ( .A(n247), .B(n805), .Y(n241) );
  AND2X2 U622 ( .A(n252), .B(n805), .Y(n242) );
  AND2X2 U623 ( .A(n246), .B(n805), .Y(n243) );
  AND2X2 U624 ( .A(n470), .B(n795), .Y(n244) );
  AND2X2 U625 ( .A(n469), .B(n795), .Y(n245) );
  AND2X2 U626 ( .A(n467), .B(n795), .Y(n246) );
  AND2X2 U627 ( .A(n468), .B(n795), .Y(n247) );
  INVX3 U628 ( .A(n705), .Y(n702) );
  CLKBUFX3 U629 ( .A(n255), .Y(n705) );
  INVX3 U630 ( .A(n705), .Y(n703) );
  CLKBUFX3 U631 ( .A(n1216), .Y(n721) );
  AND2X2 U632 ( .A(n470), .B(n796), .Y(n250) );
  AND2X2 U633 ( .A(n469), .B(n796), .Y(n251) );
  AND2X2 U634 ( .A(n467), .B(n796), .Y(n252) );
  NOR2X1 U635 ( .A(n798), .B(n797), .Y(n467) );
  AND2X2 U636 ( .A(n468), .B(n796), .Y(n253) );
  CLKBUFX3 U637 ( .A(n806), .Y(n805) );
  CLKBUFX3 U638 ( .A(n806), .Y(n804) );
  NAND2X1 U639 ( .A(n834), .B(n140), .Y(n869) );
  NAND2X1 U640 ( .A(n834), .B(n75), .Y(n905) );
  NAND2X1 U641 ( .A(n834), .B(n256), .Y(n1002) );
  CLKINVX1 U642 ( .A(n1055), .Y(n829) );
  CLKINVX1 U643 ( .A(n1057), .Y(n1227) );
  NAND2X1 U644 ( .A(n76), .B(n271), .Y(n1216) );
  NAND2X1 U645 ( .A(n75), .B(n271), .Y(n1218) );
  NAND2X1 U646 ( .A(n140), .B(n271), .Y(n1221) );
  NAND2X1 U647 ( .A(n256), .B(n271), .Y(n1223) );
  NOR2X1 U648 ( .A(n1224), .B(n1225), .Y(n140) );
  AND2X2 U649 ( .A(n1224), .B(n1225), .Y(n256) );
  CLKINVX1 U650 ( .A(proc_reset), .Y(n806) );
  CLKBUFX6 U651 ( .A(n1226), .Y(mem_read) );
  CLKINVX1 U652 ( .A(n1058), .Y(n1226) );
  CLKINVX1 U653 ( .A(tag[10]), .Y(n1035) );
  NOR3X1 U654 ( .A(n259), .B(n260), .C(n261), .Y(n823) );
  XNOR2X1 U655 ( .A(n1021), .B(proc_addr[22]), .Y(n260) );
  NOR3X1 U656 ( .A(n262), .B(n263), .C(n264), .Y(n807) );
  XNOR2X1 U657 ( .A(n1023), .B(proc_addr[21]), .Y(n262) );
  XNOR2X1 U658 ( .A(n1031), .B(proc_addr[17]), .Y(n263) );
  XNOR2X1 U659 ( .A(n1027), .B(proc_addr[19]), .Y(n264) );
  CLKMX2X2 U660 ( .A(tag[2]), .B(proc_addr[7]), .S0(n712), .Y(n268) );
  CLKMX2X2 U661 ( .A(tag[5]), .B(proc_addr[10]), .S0(n712), .Y(n269) );
  AND2X2 U662 ( .A(n1005), .B(n1004), .Y(n1052) );
  CLKINVX1 U663 ( .A(blockdata[0]), .Y(n1064) );
  CLKINVX1 U664 ( .A(blockdata[96]), .Y(n1063) );
  CLKINVX1 U665 ( .A(blockdata[1]), .Y(n1069) );
  CLKINVX1 U666 ( .A(blockdata[97]), .Y(n1068) );
  CLKINVX1 U667 ( .A(blockdata[2]), .Y(n1074) );
  CLKINVX1 U668 ( .A(blockdata[98]), .Y(n1073) );
  CLKINVX1 U669 ( .A(blockdata[3]), .Y(n1079) );
  CLKINVX1 U670 ( .A(blockdata[99]), .Y(n1078) );
  CLKINVX1 U671 ( .A(blockdata[4]), .Y(n1084) );
  CLKINVX1 U672 ( .A(blockdata[100]), .Y(n1083) );
  CLKINVX1 U673 ( .A(blockdata[5]), .Y(n1089) );
  CLKINVX1 U674 ( .A(blockdata[101]), .Y(n1088) );
  CLKINVX1 U675 ( .A(blockdata[6]), .Y(n1094) );
  CLKINVX1 U676 ( .A(blockdata[102]), .Y(n1093) );
  CLKINVX1 U677 ( .A(blockdata[7]), .Y(n1099) );
  CLKINVX1 U678 ( .A(blockdata[103]), .Y(n1098) );
  CLKINVX1 U679 ( .A(blockdata[8]), .Y(n1104) );
  CLKINVX1 U680 ( .A(blockdata[104]), .Y(n1103) );
  CLKINVX1 U681 ( .A(blockdata[9]), .Y(n1109) );
  CLKINVX1 U682 ( .A(blockdata[105]), .Y(n1108) );
  CLKINVX1 U683 ( .A(blockdata[10]), .Y(n1114) );
  CLKINVX1 U684 ( .A(blockdata[106]), .Y(n1113) );
  CLKINVX1 U685 ( .A(blockdata[11]), .Y(n1119) );
  CLKINVX1 U686 ( .A(blockdata[107]), .Y(n1118) );
  CLKINVX1 U687 ( .A(blockdata[12]), .Y(n1124) );
  CLKINVX1 U688 ( .A(blockdata[108]), .Y(n1123) );
  CLKINVX1 U689 ( .A(blockdata[13]), .Y(n1129) );
  CLKINVX1 U690 ( .A(blockdata[109]), .Y(n1128) );
  CLKINVX1 U691 ( .A(blockdata[14]), .Y(n1134) );
  CLKINVX1 U692 ( .A(blockdata[110]), .Y(n1133) );
  CLKINVX1 U693 ( .A(blockdata[15]), .Y(n1139) );
  CLKINVX1 U694 ( .A(blockdata[111]), .Y(n1138) );
  CLKINVX1 U695 ( .A(blockdata[16]), .Y(n1144) );
  CLKINVX1 U696 ( .A(blockdata[112]), .Y(n1143) );
  CLKINVX1 U697 ( .A(blockdata[17]), .Y(n1149) );
  CLKINVX1 U698 ( .A(blockdata[113]), .Y(n1148) );
  CLKINVX1 U699 ( .A(blockdata[18]), .Y(n1154) );
  CLKINVX1 U700 ( .A(blockdata[114]), .Y(n1153) );
  CLKINVX1 U701 ( .A(blockdata[19]), .Y(n1159) );
  CLKINVX1 U702 ( .A(blockdata[115]), .Y(n1158) );
  CLKINVX1 U703 ( .A(blockdata[20]), .Y(n1164) );
  CLKINVX1 U704 ( .A(blockdata[116]), .Y(n1163) );
  CLKINVX1 U705 ( .A(blockdata[21]), .Y(n1169) );
  CLKINVX1 U706 ( .A(blockdata[117]), .Y(n1168) );
  CLKINVX1 U707 ( .A(blockdata[22]), .Y(n1174) );
  CLKINVX1 U708 ( .A(blockdata[118]), .Y(n1173) );
  CLKINVX1 U709 ( .A(blockdata[23]), .Y(n1179) );
  CLKINVX1 U710 ( .A(blockdata[119]), .Y(n1178) );
  CLKINVX1 U711 ( .A(blockdata[24]), .Y(n1184) );
  CLKINVX1 U712 ( .A(blockdata[120]), .Y(n1183) );
  CLKINVX1 U713 ( .A(blockdata[25]), .Y(n1189) );
  CLKINVX1 U714 ( .A(blockdata[121]), .Y(n1188) );
  CLKINVX1 U715 ( .A(blockdata[26]), .Y(n1194) );
  CLKINVX1 U716 ( .A(blockdata[122]), .Y(n1193) );
  CLKINVX1 U717 ( .A(blockdata[27]), .Y(n1199) );
  CLKINVX1 U718 ( .A(blockdata[123]), .Y(n1198) );
  CLKINVX1 U719 ( .A(blockdata[28]), .Y(n1204) );
  CLKINVX1 U720 ( .A(blockdata[124]), .Y(n1203) );
  CLKINVX1 U721 ( .A(blockdata[29]), .Y(n1209) );
  CLKINVX1 U722 ( .A(blockdata[125]), .Y(n1208) );
  CLKINVX1 U723 ( .A(blockdata[30]), .Y(n1214) );
  CLKINVX1 U724 ( .A(blockdata[126]), .Y(n1213) );
  CLKINVX1 U725 ( .A(blockdata[31]), .Y(n1222) );
  CLKINVX1 U726 ( .A(blockdata[127]), .Y(n1220) );
  CLKINVX1 U727 ( .A(blockdata[32]), .Y(n1060) );
  CLKINVX1 U728 ( .A(blockdata[33]), .Y(n1065) );
  CLKINVX1 U729 ( .A(blockdata[34]), .Y(n1070) );
  CLKINVX1 U730 ( .A(blockdata[35]), .Y(n1075) );
  CLKINVX1 U731 ( .A(blockdata[36]), .Y(n1080) );
  CLKINVX1 U732 ( .A(blockdata[37]), .Y(n1085) );
  CLKINVX1 U733 ( .A(blockdata[38]), .Y(n1090) );
  CLKINVX1 U734 ( .A(blockdata[39]), .Y(n1095) );
  CLKINVX1 U735 ( .A(blockdata[40]), .Y(n1100) );
  CLKINVX1 U736 ( .A(blockdata[41]), .Y(n1105) );
  CLKINVX1 U737 ( .A(blockdata[42]), .Y(n1110) );
  CLKINVX1 U738 ( .A(blockdata[43]), .Y(n1115) );
  CLKINVX1 U739 ( .A(blockdata[44]), .Y(n1120) );
  CLKINVX1 U740 ( .A(blockdata[45]), .Y(n1125) );
  CLKINVX1 U741 ( .A(blockdata[46]), .Y(n1130) );
  CLKINVX1 U742 ( .A(blockdata[47]), .Y(n1135) );
  CLKINVX1 U743 ( .A(blockdata[48]), .Y(n1140) );
  CLKINVX1 U744 ( .A(blockdata[49]), .Y(n1145) );
  CLKINVX1 U745 ( .A(blockdata[50]), .Y(n1150) );
  CLKINVX1 U746 ( .A(blockdata[51]), .Y(n1155) );
  CLKINVX1 U747 ( .A(blockdata[52]), .Y(n1160) );
  CLKINVX1 U748 ( .A(blockdata[53]), .Y(n1165) );
  CLKINVX1 U749 ( .A(blockdata[54]), .Y(n1170) );
  CLKINVX1 U750 ( .A(blockdata[55]), .Y(n1175) );
  CLKINVX1 U751 ( .A(blockdata[56]), .Y(n1180) );
  CLKINVX1 U752 ( .A(blockdata[57]), .Y(n1185) );
  CLKINVX1 U753 ( .A(blockdata[58]), .Y(n1190) );
  CLKINVX1 U754 ( .A(blockdata[59]), .Y(n1195) );
  CLKINVX1 U755 ( .A(blockdata[60]), .Y(n1200) );
  CLKINVX1 U756 ( .A(blockdata[61]), .Y(n1205) );
  CLKINVX1 U757 ( .A(blockdata[62]), .Y(n1210) );
  CLKINVX1 U758 ( .A(blockdata[63]), .Y(n1215) );
  CLKINVX1 U759 ( .A(blockdata[64]), .Y(n1061) );
  CLKINVX1 U760 ( .A(blockdata[65]), .Y(n1066) );
  CLKINVX1 U761 ( .A(blockdata[66]), .Y(n1071) );
  CLKINVX1 U762 ( .A(blockdata[67]), .Y(n1076) );
  CLKINVX1 U763 ( .A(blockdata[68]), .Y(n1081) );
  CLKINVX1 U764 ( .A(blockdata[69]), .Y(n1086) );
  CLKINVX1 U765 ( .A(blockdata[70]), .Y(n1091) );
  CLKINVX1 U766 ( .A(blockdata[71]), .Y(n1096) );
  CLKINVX1 U767 ( .A(blockdata[72]), .Y(n1101) );
  CLKINVX1 U768 ( .A(blockdata[73]), .Y(n1106) );
  CLKINVX1 U769 ( .A(blockdata[74]), .Y(n1111) );
  CLKINVX1 U770 ( .A(blockdata[75]), .Y(n1116) );
  CLKINVX1 U771 ( .A(blockdata[76]), .Y(n1121) );
  CLKINVX1 U772 ( .A(blockdata[77]), .Y(n1126) );
  CLKINVX1 U773 ( .A(blockdata[78]), .Y(n1131) );
  CLKINVX1 U774 ( .A(blockdata[79]), .Y(n1136) );
  CLKINVX1 U775 ( .A(blockdata[80]), .Y(n1141) );
  CLKINVX1 U776 ( .A(blockdata[81]), .Y(n1146) );
  CLKINVX1 U777 ( .A(blockdata[82]), .Y(n1151) );
  CLKINVX1 U778 ( .A(blockdata[83]), .Y(n1156) );
  CLKINVX1 U779 ( .A(blockdata[84]), .Y(n1161) );
  CLKINVX1 U780 ( .A(blockdata[85]), .Y(n1166) );
  CLKINVX1 U781 ( .A(blockdata[86]), .Y(n1171) );
  CLKINVX1 U782 ( .A(blockdata[87]), .Y(n1176) );
  CLKINVX1 U783 ( .A(blockdata[88]), .Y(n1181) );
  CLKINVX1 U784 ( .A(blockdata[89]), .Y(n1186) );
  CLKINVX1 U785 ( .A(blockdata[90]), .Y(n1191) );
  CLKINVX1 U786 ( .A(blockdata[91]), .Y(n1196) );
  CLKINVX1 U787 ( .A(blockdata[92]), .Y(n1201) );
  CLKINVX1 U788 ( .A(blockdata[93]), .Y(n1206) );
  CLKINVX1 U789 ( .A(blockdata[94]), .Y(n1211) );
  CLKINVX1 U790 ( .A(blockdata[95]), .Y(n1217) );
  NAND2X1 U791 ( .A(mem_rdata[32]), .B(n716), .Y(n937) );
  NAND2X1 U792 ( .A(mem_rdata[33]), .B(n715), .Y(n936) );
  NAND2X1 U793 ( .A(mem_rdata[34]), .B(n719), .Y(n935) );
  NAND2X1 U794 ( .A(mem_rdata[35]), .B(n718), .Y(n934) );
  NAND2X1 U795 ( .A(mem_rdata[36]), .B(n716), .Y(n933) );
  NAND2X1 U796 ( .A(mem_rdata[37]), .B(n717), .Y(n932) );
  NAND2X1 U797 ( .A(mem_rdata[38]), .B(n714), .Y(n931) );
  NAND2X1 U798 ( .A(mem_rdata[39]), .B(n717), .Y(n930) );
  NAND2X1 U799 ( .A(mem_rdata[40]), .B(n715), .Y(n929) );
  NAND2X1 U800 ( .A(mem_rdata[41]), .B(n715), .Y(n928) );
  NAND2X1 U801 ( .A(mem_rdata[42]), .B(n715), .Y(n927) );
  NAND2X1 U802 ( .A(mem_rdata[43]), .B(n715), .Y(n926) );
  NAND2X1 U803 ( .A(mem_rdata[44]), .B(n715), .Y(n925) );
  NAND2X1 U804 ( .A(mem_rdata[45]), .B(n715), .Y(n924) );
  NAND2X1 U805 ( .A(mem_rdata[46]), .B(n715), .Y(n923) );
  NAND2X1 U806 ( .A(mem_rdata[47]), .B(n715), .Y(n922) );
  NAND2X1 U807 ( .A(mem_rdata[48]), .B(n715), .Y(n921) );
  NAND2X1 U808 ( .A(mem_rdata[49]), .B(n715), .Y(n920) );
  NAND2X1 U809 ( .A(mem_rdata[50]), .B(n715), .Y(n919) );
  NAND2X1 U810 ( .A(mem_rdata[51]), .B(n715), .Y(n918) );
  NAND2X1 U811 ( .A(mem_rdata[52]), .B(n715), .Y(n917) );
  NAND2X1 U812 ( .A(mem_rdata[53]), .B(n716), .Y(n916) );
  NAND2X1 U813 ( .A(mem_rdata[54]), .B(n716), .Y(n915) );
  NAND2X1 U814 ( .A(mem_rdata[55]), .B(n716), .Y(n914) );
  NAND2X1 U815 ( .A(mem_rdata[56]), .B(n716), .Y(n913) );
  NAND2X1 U816 ( .A(mem_rdata[57]), .B(n716), .Y(n912) );
  NAND2X1 U817 ( .A(mem_rdata[58]), .B(n716), .Y(n911) );
  NAND2X1 U818 ( .A(mem_rdata[59]), .B(n716), .Y(n910) );
  NAND2X1 U819 ( .A(mem_rdata[60]), .B(n716), .Y(n909) );
  NAND2X1 U820 ( .A(mem_rdata[61]), .B(n716), .Y(n908) );
  NAND2X1 U821 ( .A(mem_rdata[62]), .B(n716), .Y(n907) );
  NAND2X1 U822 ( .A(mem_rdata[63]), .B(n716), .Y(n906) );
  NAND2X1 U823 ( .A(mem_rdata[64]), .B(n716), .Y(n903) );
  NAND2X1 U824 ( .A(mem_rdata[65]), .B(n716), .Y(n902) );
  NAND2X1 U825 ( .A(mem_rdata[66]), .B(n717), .Y(n901) );
  NAND2X1 U826 ( .A(mem_rdata[67]), .B(n717), .Y(n900) );
  NAND2X1 U827 ( .A(mem_rdata[68]), .B(n717), .Y(n899) );
  NAND2X1 U828 ( .A(mem_rdata[69]), .B(n717), .Y(n898) );
  NAND2X1 U829 ( .A(mem_rdata[70]), .B(n717), .Y(n897) );
  NAND2X1 U830 ( .A(mem_rdata[71]), .B(n717), .Y(n896) );
  NAND2X1 U831 ( .A(mem_rdata[72]), .B(n717), .Y(n895) );
  NAND2X1 U832 ( .A(mem_rdata[73]), .B(n717), .Y(n894) );
  NAND2X1 U833 ( .A(mem_rdata[74]), .B(n717), .Y(n893) );
  NAND2X1 U834 ( .A(mem_rdata[75]), .B(n717), .Y(n892) );
  NAND2X1 U835 ( .A(mem_rdata[76]), .B(n717), .Y(n891) );
  NAND2X1 U836 ( .A(mem_rdata[77]), .B(n717), .Y(n890) );
  NAND2X1 U837 ( .A(mem_rdata[78]), .B(n717), .Y(n889) );
  NAND2X1 U838 ( .A(mem_rdata[79]), .B(n718), .Y(n888) );
  NAND2X1 U839 ( .A(mem_rdata[80]), .B(n718), .Y(n887) );
  NAND2X1 U840 ( .A(mem_rdata[81]), .B(n718), .Y(n886) );
  NAND2X1 U841 ( .A(mem_rdata[82]), .B(n718), .Y(n885) );
  NAND2X1 U842 ( .A(mem_rdata[83]), .B(n718), .Y(n884) );
  NAND2X1 U843 ( .A(mem_rdata[84]), .B(n718), .Y(n883) );
  NAND2X1 U844 ( .A(mem_rdata[85]), .B(n718), .Y(n882) );
  NAND2X1 U845 ( .A(mem_rdata[86]), .B(n718), .Y(n881) );
  NAND2X1 U846 ( .A(mem_rdata[87]), .B(n718), .Y(n880) );
  NAND2X1 U847 ( .A(mem_rdata[88]), .B(n718), .Y(n879) );
  NAND2X1 U848 ( .A(mem_rdata[89]), .B(n718), .Y(n878) );
  NAND2X1 U849 ( .A(mem_rdata[90]), .B(n718), .Y(n877) );
  NAND2X1 U850 ( .A(mem_rdata[91]), .B(n718), .Y(n876) );
  NAND2X1 U851 ( .A(mem_rdata[92]), .B(n719), .Y(n875) );
  NAND2X1 U852 ( .A(mem_rdata[93]), .B(n719), .Y(n874) );
  NAND2X1 U853 ( .A(mem_rdata[94]), .B(n719), .Y(n873) );
  NAND2X1 U854 ( .A(mem_rdata[95]), .B(n719), .Y(n872) );
  NAND2X1 U855 ( .A(mem_rdata[96]), .B(n719), .Y(n867) );
  NAND2X1 U856 ( .A(mem_rdata[97]), .B(n719), .Y(n866) );
  NAND2X1 U857 ( .A(mem_rdata[98]), .B(n719), .Y(n865) );
  NAND2X1 U858 ( .A(mem_rdata[99]), .B(n719), .Y(n864) );
  NAND2X1 U859 ( .A(mem_rdata[100]), .B(n719), .Y(n863) );
  NAND2X1 U860 ( .A(mem_rdata[101]), .B(n719), .Y(n862) );
  NAND2X1 U861 ( .A(mem_rdata[102]), .B(n719), .Y(n861) );
  NAND2X1 U862 ( .A(mem_rdata[103]), .B(n719), .Y(n860) );
  NAND2X1 U863 ( .A(mem_rdata[104]), .B(n719), .Y(n859) );
  NAND2X1 U864 ( .A(mem_rdata[105]), .B(n720), .Y(n858) );
  NAND2X1 U865 ( .A(mem_rdata[106]), .B(n720), .Y(n857) );
  NAND2X1 U866 ( .A(mem_rdata[107]), .B(n720), .Y(n856) );
  NAND2X1 U867 ( .A(mem_rdata[108]), .B(n713), .Y(n855) );
  NAND2X1 U868 ( .A(mem_rdata[109]), .B(n713), .Y(n854) );
  NAND2X1 U869 ( .A(mem_rdata[110]), .B(n716), .Y(n853) );
  NAND2X1 U870 ( .A(mem_rdata[111]), .B(n717), .Y(n852) );
  NAND2X1 U871 ( .A(mem_rdata[112]), .B(n718), .Y(n851) );
  NAND2X1 U872 ( .A(mem_rdata[113]), .B(n718), .Y(n850) );
  NAND2X1 U873 ( .A(mem_rdata[114]), .B(n714), .Y(n849) );
  NAND2X1 U874 ( .A(mem_rdata[115]), .B(n719), .Y(n848) );
  NAND2X1 U875 ( .A(mem_rdata[116]), .B(n715), .Y(n847) );
  NAND2X1 U876 ( .A(mem_rdata[117]), .B(n715), .Y(n846) );
  NAND2X1 U877 ( .A(mem_rdata[118]), .B(n720), .Y(n845) );
  NAND2X1 U878 ( .A(mem_rdata[119]), .B(n720), .Y(n844) );
  NAND2X1 U879 ( .A(mem_rdata[120]), .B(n720), .Y(n843) );
  NAND2X1 U880 ( .A(mem_rdata[121]), .B(n720), .Y(n842) );
  NAND2X1 U881 ( .A(mem_rdata[122]), .B(n720), .Y(n841) );
  NAND2X1 U882 ( .A(mem_rdata[123]), .B(n720), .Y(n840) );
  NAND2X1 U883 ( .A(mem_rdata[124]), .B(n720), .Y(n839) );
  NAND2X1 U884 ( .A(mem_rdata[125]), .B(n720), .Y(n838) );
  NAND2X1 U885 ( .A(mem_rdata[126]), .B(n720), .Y(n837) );
  NAND2X1 U886 ( .A(mem_rdata[127]), .B(n720), .Y(n836) );
  NAND2X1 U887 ( .A(mem_rdata[1]), .B(n714), .Y(n998) );
  NAND2X1 U888 ( .A(mem_rdata[2]), .B(n714), .Y(n996) );
  NAND2X1 U889 ( .A(mem_rdata[3]), .B(n714), .Y(n994) );
  NAND2X1 U890 ( .A(mem_rdata[4]), .B(n714), .Y(n992) );
  NAND2X1 U891 ( .A(mem_rdata[5]), .B(n714), .Y(n990) );
  NAND2X1 U892 ( .A(mem_rdata[6]), .B(n714), .Y(n988) );
  NAND2X1 U893 ( .A(mem_rdata[7]), .B(n714), .Y(n986) );
  NAND2X1 U894 ( .A(mem_rdata[8]), .B(n714), .Y(n984) );
  NAND2X1 U895 ( .A(mem_rdata[9]), .B(n714), .Y(n982) );
  NAND2X1 U896 ( .A(mem_rdata[10]), .B(n714), .Y(n980) );
  NAND2X1 U897 ( .A(mem_rdata[11]), .B(n714), .Y(n978) );
  NAND2X1 U898 ( .A(mem_rdata[12]), .B(n714), .Y(n976) );
  NAND2X1 U899 ( .A(mem_rdata[13]), .B(n714), .Y(n974) );
  NAND2X1 U900 ( .A(mem_rdata[14]), .B(n718), .Y(n972) );
  NAND2X1 U901 ( .A(mem_rdata[15]), .B(n716), .Y(n970) );
  NAND2X1 U902 ( .A(mem_rdata[16]), .B(n717), .Y(n968) );
  NAND2X1 U903 ( .A(mem_rdata[17]), .B(n719), .Y(n966) );
  NAND2X1 U904 ( .A(mem_rdata[18]), .B(n714), .Y(n964) );
  NAND2X1 U905 ( .A(mem_rdata[19]), .B(n715), .Y(n962) );
  NAND2X1 U906 ( .A(mem_rdata[20]), .B(n718), .Y(n960) );
  NAND2X1 U907 ( .A(mem_rdata[21]), .B(n716), .Y(n958) );
  NAND2X1 U908 ( .A(mem_rdata[22]), .B(n717), .Y(n956) );
  NAND2X1 U909 ( .A(mem_rdata[23]), .B(n719), .Y(n954) );
  NAND2X1 U910 ( .A(mem_rdata[24]), .B(n712), .Y(n952) );
  NAND2X1 U911 ( .A(mem_rdata[25]), .B(n714), .Y(n950) );
  NAND2X1 U912 ( .A(mem_rdata[26]), .B(n715), .Y(n948) );
  NAND2X1 U913 ( .A(mem_rdata[27]), .B(n719), .Y(n946) );
  NAND2X1 U914 ( .A(mem_rdata[28]), .B(n718), .Y(n944) );
  NAND2X1 U915 ( .A(mem_rdata[29]), .B(n716), .Y(n942) );
  NAND2X1 U916 ( .A(mem_rdata[30]), .B(n717), .Y(n940) );
  NAND2X1 U917 ( .A(mem_rdata[31]), .B(n714), .Y(n938) );
  INVXL U918 ( .A(proc_write), .Y(n1059) );
  MXI4X1 U919 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n683), .S1(n659), .Y(
        n604) );
  MXI4X1 U920 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n683), .S1(n659), .Y(
        n605) );
  MXI4X1 U921 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n661), .S1(n659), .Y(
        n590) );
  MXI4X1 U922 ( .A(\blocktag[4][17] ), .B(\blocktag[5][17] ), .C(
        \blocktag[6][17] ), .D(\blocktag[7][17] ), .S0(n662), .S1(n658), .Y(
        n591) );
  MXI4X1 U923 ( .A(\blocktag[0][22] ), .B(\blocktag[1][22] ), .C(
        \blocktag[2][22] ), .D(\blocktag[3][22] ), .S0(n682), .S1(n655), .Y(
        n582) );
  MXI4X1 U924 ( .A(\blocktag[4][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[7][22] ), .S0(n682), .S1(n655), .Y(
        n583) );
  MXI4X1 U925 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n685), .S1(n658), .Y(
        n596) );
  MXI4X1 U926 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n685), .S1(n658), .Y(
        n597) );
  MXI4X1 U927 ( .A(\blocktag[0][12] ), .B(\blocktag[1][12] ), .C(
        \blocktag[2][12] ), .D(\blocktag[3][12] ), .S0(n683), .S1(n659), .Y(
        n600) );
  MXI4X1 U928 ( .A(\blocktag[4][12] ), .B(\blocktag[5][12] ), .C(
        \blocktag[6][12] ), .D(\blocktag[7][12] ), .S0(n683), .S1(n659), .Y(
        n601) );
  MXI2X1 U929 ( .A(n598), .B(n599), .S0(n628), .Y(tag[13]) );
  MXI2X1 U930 ( .A(n588), .B(n589), .S0(n628), .Y(tag[19]) );
  MXI2X1 U931 ( .A(n586), .B(n587), .S0(n628), .Y(tag[20]) );
  MXI2X1 U932 ( .A(n602), .B(n603), .S0(N33), .Y(tag[11]) );
  CLKINVX1 U933 ( .A(n831), .Y(n870) );
  OAI211X1 U934 ( .A0(mem_ready), .A1(valid), .B0(n830), .C0(n1054), .Y(n831)
         );
  INVXL U935 ( .A(proc_addr[13]), .Y(n1038) );
  MXI2X1 U936 ( .A(n510), .B(n511), .S0(n625), .Y(blockdata[32]) );
  MXI4X1 U937 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n676), .S1(n650), .Y(n511) );
  MXI4X1 U938 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n672), .S1(n650), .Y(n510) );
  MXI2X1 U939 ( .A(n410), .B(n411), .S0(n625), .Y(blockdata[64]) );
  MXI4X1 U940 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n675), .S1(n645), .Y(n411) );
  MXI4X1 U941 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n675), .S1(n645), .Y(n410) );
  MXI2X1 U942 ( .A(n508), .B(n509), .S0(n624), .Y(blockdata[33]) );
  MXI4X1 U943 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n677), .S1(n649), .Y(n509) );
  MXI4X1 U944 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n674), .S1(n649), .Y(n508) );
  MXI2X1 U945 ( .A(n408), .B(n409), .S0(n625), .Y(blockdata[65]) );
  MXI4X1 U946 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n675), .S1(n645), .Y(n409) );
  MXI4X1 U947 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n675), .S1(n645), .Y(n408) );
  MXI2X1 U948 ( .A(n506), .B(n507), .S0(n624), .Y(blockdata[34]) );
  MXI4X1 U949 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n679), .S1(n649), .Y(n507) );
  MXI4X1 U950 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n671), .S1(n649), .Y(n506) );
  MXI2X1 U951 ( .A(n406), .B(n407), .S0(n625), .Y(blockdata[66]) );
  MXI4X1 U952 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n675), .S1(n645), .Y(n407) );
  MXI4X1 U953 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n675), .S1(n645), .Y(n406) );
  MXI2X1 U954 ( .A(n504), .B(n505), .S0(n624), .Y(blockdata[35]) );
  MXI4X1 U955 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n678), .S1(n649), .Y(n505) );
  MXI4X1 U956 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n669), .S1(n649), .Y(n504) );
  MXI2X1 U957 ( .A(n404), .B(n405), .S0(n623), .Y(blockdata[67]) );
  MXI4X1 U958 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n675), .S1(n645), .Y(n405) );
  MXI4X1 U959 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n675), .S1(n645), .Y(n404) );
  MXI2X1 U960 ( .A(n466), .B(n502), .S0(n624), .Y(blockdata[36]) );
  MXI4X1 U961 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n675), .S1(n649), .Y(n502) );
  MXI4X1 U962 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n668), .S1(n649), .Y(n466) );
  MXI2X1 U963 ( .A(n402), .B(n403), .S0(n625), .Y(blockdata[68]) );
  MXI4X1 U964 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n675), .S1(n645), .Y(n403) );
  MXI4X1 U965 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n675), .S1(n645), .Y(n402) );
  MXI2X1 U966 ( .A(n464), .B(n465), .S0(n624), .Y(blockdata[37]) );
  MXI4X1 U967 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n673), .S1(n649), .Y(n465) );
  MXI4X1 U968 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n684), .S1(n649), .Y(n464) );
  MXI2X1 U969 ( .A(n400), .B(n401), .S0(n626), .Y(blockdata[69]) );
  MXI4X1 U970 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n675), .S1(n644), .Y(n401) );
  MXI4X1 U971 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n675), .S1(n644), .Y(n400) );
  MXI2X1 U972 ( .A(n462), .B(n463), .S0(n624), .Y(blockdata[38]) );
  MXI4X1 U973 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n679), .S1(n649), .Y(n463) );
  MXI4X1 U974 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n679), .S1(n649), .Y(n462) );
  MXI2X1 U975 ( .A(n398), .B(n399), .S0(n626), .Y(blockdata[70]) );
  MXI4X1 U976 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n674), .S1(n644), .Y(n399) );
  MXI4X1 U977 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n675), .S1(n644), .Y(n398) );
  MXI2X1 U978 ( .A(n460), .B(n461), .S0(n624), .Y(blockdata[39]) );
  MXI4X1 U979 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n679), .S1(n648), .Y(n461) );
  MXI4X1 U980 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n679), .S1(n648), .Y(n460) );
  MXI2X1 U981 ( .A(n396), .B(n397), .S0(n622), .Y(blockdata[71]) );
  MXI4X1 U982 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n674), .S1(n644), .Y(n397) );
  MXI4X1 U983 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n674), .S1(n644), .Y(n396) );
  MXI2X1 U984 ( .A(n458), .B(n459), .S0(n624), .Y(blockdata[40]) );
  MXI4X1 U985 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n679), .S1(n648), .Y(n459) );
  MXI4X1 U986 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n679), .S1(n648), .Y(n458) );
  MXI2X1 U987 ( .A(n394), .B(n395), .S0(n621), .Y(blockdata[72]) );
  MXI4X1 U988 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n674), .S1(n644), .Y(n395) );
  MXI4X1 U989 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n674), .S1(n644), .Y(n394) );
  MXI2X1 U990 ( .A(n456), .B(n457), .S0(n624), .Y(blockdata[41]) );
  MXI4X1 U991 ( .A(\block[4][41] ), .B(\block[5][41] ), .C(\block[6][41] ), 
        .D(\block[7][41] ), .S0(n679), .S1(n648), .Y(n457) );
  MXI4X1 U992 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n679), .S1(n648), .Y(n456) );
  MXI2X1 U993 ( .A(n392), .B(n393), .S0(n622), .Y(blockdata[73]) );
  MXI4X1 U994 ( .A(\block[4][73] ), .B(\block[5][73] ), .C(\block[6][73] ), 
        .D(\block[7][73] ), .S0(n674), .S1(n644), .Y(n393) );
  MXI4X1 U995 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n674), .S1(n644), .Y(n392) );
  MXI2X1 U996 ( .A(n454), .B(n455), .S0(n624), .Y(blockdata[42]) );
  MXI4X1 U997 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n679), .S1(n648), .Y(n455) );
  MXI4X1 U998 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n679), .S1(n648), .Y(n454) );
  MXI2X1 U999 ( .A(n390), .B(n391), .S0(n627), .Y(blockdata[74]) );
  MXI4X1 U1000 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n674), .S1(n644), .Y(n391) );
  MXI4X1 U1001 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n674), .S1(n644), .Y(n390) );
  MXI2X1 U1002 ( .A(n452), .B(n453), .S0(n624), .Y(blockdata[43]) );
  MXI4X1 U1003 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n679), .S1(n648), .Y(n453) );
  MXI4X1 U1004 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n679), .S1(n648), .Y(n452) );
  MXI2X1 U1005 ( .A(n388), .B(n389), .S0(n627), .Y(blockdata[75]) );
  MXI4X1 U1006 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n674), .S1(n643), .Y(n389) );
  MXI4X1 U1007 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n674), .S1(n643), .Y(n388) );
  MXI2X1 U1008 ( .A(n450), .B(n451), .S0(n624), .Y(blockdata[44]) );
  MXI4X1 U1009 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n678), .S1(n648), .Y(n451) );
  MXI4X1 U1010 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n679), .S1(n648), .Y(n450) );
  MXI2X1 U1011 ( .A(n386), .B(n387), .S0(n627), .Y(blockdata[76]) );
  MXI4X1 U1012 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n674), .S1(n643), .Y(n387) );
  MXI4X1 U1013 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n674), .S1(n643), .Y(n386) );
  MXI2X1 U1014 ( .A(n448), .B(n449), .S0(n623), .Y(blockdata[45]) );
  MXI4X1 U1015 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n678), .S1(n647), .Y(n449) );
  MXI4X1 U1016 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n678), .S1(n647), .Y(n448) );
  MXI2X1 U1017 ( .A(n384), .B(n385), .S0(n627), .Y(blockdata[77]) );
  MXI4X1 U1018 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n673), .S1(n643), .Y(n385) );
  MXI4X1 U1019 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n673), .S1(n643), .Y(n384) );
  MXI2X1 U1020 ( .A(n446), .B(n447), .S0(n623), .Y(blockdata[46]) );
  MXI4X1 U1021 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n678), .S1(n647), .Y(n447) );
  MXI4X1 U1022 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n678), .S1(n647), .Y(n446) );
  MXI2X1 U1023 ( .A(n382), .B(n383), .S0(n627), .Y(blockdata[78]) );
  MXI4X1 U1024 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n673), .S1(n643), .Y(n383) );
  MXI4X1 U1025 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n673), .S1(n643), .Y(n382) );
  MXI2X1 U1026 ( .A(n444), .B(n445), .S0(n623), .Y(blockdata[47]) );
  MXI4X1 U1027 ( .A(\block[4][47] ), .B(\block[5][47] ), .C(\block[6][47] ), 
        .D(\block[7][47] ), .S0(n678), .S1(n647), .Y(n445) );
  MXI4X1 U1028 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n678), .S1(n647), .Y(n444) );
  MXI2X1 U1029 ( .A(n380), .B(n381), .S0(n627), .Y(blockdata[79]) );
  MXI4X1 U1030 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n673), .S1(n643), .Y(n381) );
  MXI4X1 U1031 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n673), .S1(n643), .Y(n380) );
  MXI2X1 U1032 ( .A(n442), .B(n443), .S0(n623), .Y(blockdata[48]) );
  MXI4X1 U1033 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n678), .S1(n647), .Y(n443) );
  MXI4X1 U1034 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n678), .S1(n647), .Y(n442) );
  MXI2X1 U1035 ( .A(n378), .B(n379), .S0(n627), .Y(blockdata[80]) );
  MXI4X1 U1036 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n673), .S1(n643), .Y(n379) );
  MXI4X1 U1037 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n673), .S1(n643), .Y(n378) );
  MXI2X1 U1038 ( .A(n440), .B(n441), .S0(n623), .Y(blockdata[49]) );
  MXI4X1 U1039 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n678), .S1(n647), .Y(n441) );
  MXI4X1 U1040 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n678), .S1(n647), .Y(n440) );
  MXI2X1 U1041 ( .A(n376), .B(n377), .S0(n622), .Y(blockdata[81]) );
  MXI4X1 U1042 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n673), .S1(n642), .Y(n377) );
  MXI4X1 U1043 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n673), .S1(n642), .Y(n376) );
  MXI2X1 U1044 ( .A(n438), .B(n439), .S0(n623), .Y(blockdata[50]) );
  MXI4X1 U1045 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n678), .S1(n647), .Y(n439) );
  MXI4X1 U1046 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n678), .S1(n647), .Y(n438) );
  MXI2X1 U1047 ( .A(n374), .B(n375), .S0(n622), .Y(blockdata[82]) );
  MXI4X1 U1048 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n673), .S1(n642), .Y(n375) );
  MXI4X1 U1049 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n673), .S1(n642), .Y(n374) );
  MXI2X1 U1050 ( .A(n436), .B(n437), .S0(n623), .Y(blockdata[51]) );
  MXI4X1 U1051 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n677), .S1(n646), .Y(n437) );
  MXI4X1 U1052 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n677), .S1(n646), .Y(n436) );
  MXI2X1 U1053 ( .A(n372), .B(n373), .S0(n622), .Y(blockdata[83]) );
  MXI4X1 U1054 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n672), .S1(n642), .Y(n373) );
  MXI4X1 U1055 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n673), .S1(n642), .Y(n372) );
  MXI2X1 U1056 ( .A(n434), .B(n435), .S0(n623), .Y(blockdata[52]) );
  MXI4X1 U1057 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n677), .S1(n646), .Y(n435) );
  MXI4X1 U1058 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n677), .S1(n646), .Y(n434) );
  MXI2X1 U1059 ( .A(n370), .B(n371), .S0(n622), .Y(blockdata[84]) );
  MXI4X1 U1060 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n672), .S1(n642), .Y(n371) );
  MXI4X1 U1061 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n672), .S1(n642), .Y(n370) );
  MXI2X1 U1062 ( .A(n432), .B(n433), .S0(n623), .Y(blockdata[53]) );
  MXI4X1 U1063 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n677), .S1(n646), .Y(n433) );
  MXI4X1 U1064 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n677), .S1(n646), .Y(n432) );
  MXI2X1 U1065 ( .A(n368), .B(n369), .S0(n622), .Y(blockdata[85]) );
  MXI4X1 U1066 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n672), .S1(n642), .Y(n369) );
  MXI4X1 U1067 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n672), .S1(n642), .Y(n368) );
  MXI2X1 U1068 ( .A(n430), .B(n431), .S0(n623), .Y(blockdata[54]) );
  MXI4X1 U1069 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n677), .S1(n646), .Y(n431) );
  MXI4X1 U1070 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n677), .S1(n646), .Y(n430) );
  MXI2X1 U1071 ( .A(n366), .B(n367), .S0(n622), .Y(blockdata[86]) );
  MXI4X1 U1072 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n672), .S1(n642), .Y(n367) );
  MXI4X1 U1073 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n672), .S1(n642), .Y(n366) );
  MXI2X1 U1074 ( .A(n428), .B(n429), .S0(n623), .Y(blockdata[55]) );
  MXI4X1 U1075 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n677), .S1(n646), .Y(n429) );
  MXI4X1 U1076 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n677), .S1(n646), .Y(n428) );
  MXI2X1 U1077 ( .A(n364), .B(n365), .S0(n622), .Y(blockdata[87]) );
  MXI4X1 U1078 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n672), .S1(n641), .Y(n365) );
  MXI4X1 U1079 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n672), .S1(n641), .Y(n364) );
  MXI2X1 U1080 ( .A(n426), .B(n427), .S0(n623), .Y(blockdata[56]) );
  MXI4X1 U1081 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n677), .S1(n646), .Y(n427) );
  MXI4X1 U1082 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n677), .S1(n646), .Y(n426) );
  MXI2X1 U1083 ( .A(n362), .B(n363), .S0(n622), .Y(blockdata[88]) );
  MXI4X1 U1084 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n672), .S1(n641), .Y(n363) );
  MXI4X1 U1085 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n672), .S1(n641), .Y(n362) );
  MXI2X1 U1086 ( .A(n424), .B(n425), .S0(n620), .Y(blockdata[57]) );
  MXI4X1 U1087 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n676), .S1(n647), .Y(n425) );
  MXI4X1 U1088 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n677), .S1(n645), .Y(n424) );
  MXI2X1 U1089 ( .A(n360), .B(n361), .S0(n622), .Y(blockdata[89]) );
  MXI4X1 U1090 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n672), .S1(n641), .Y(n361) );
  MXI4X1 U1091 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n672), .S1(n641), .Y(n360) );
  MXI2X1 U1092 ( .A(n422), .B(n423), .S0(n623), .Y(blockdata[58]) );
  MXI4X1 U1093 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n676), .S1(n648), .Y(n423) );
  MXI4X1 U1094 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n676), .S1(n650), .Y(n422) );
  MXI2X1 U1095 ( .A(n358), .B(n359), .S0(n622), .Y(blockdata[90]) );
  MXI4X1 U1096 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n671), .S1(n641), .Y(n359) );
  MXI4X1 U1097 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n671), .S1(n641), .Y(n358) );
  MXI2X1 U1098 ( .A(n420), .B(n421), .S0(n622), .Y(blockdata[59]) );
  MXI4X1 U1099 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n676), .S1(n646), .Y(n421) );
  MXI4X1 U1100 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n676), .S1(n647), .Y(n420) );
  MXI2X1 U1101 ( .A(n356), .B(n357), .S0(n622), .Y(blockdata[91]) );
  MXI4X1 U1102 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n671), .S1(n641), .Y(n357) );
  MXI4X1 U1103 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n671), .S1(n641), .Y(n356) );
  MXI2X1 U1104 ( .A(n418), .B(n419), .S0(n623), .Y(blockdata[60]) );
  MXI4X1 U1105 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n676), .S1(n648), .Y(n419) );
  MXI4X1 U1106 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n676), .S1(n637), .Y(n418) );
  MXI2X1 U1107 ( .A(n354), .B(n355), .S0(n622), .Y(blockdata[92]) );
  MXI4X1 U1108 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n671), .S1(n641), .Y(n355) );
  MXI4X1 U1109 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n671), .S1(n641), .Y(n354) );
  MXI2X1 U1110 ( .A(n416), .B(n417), .S0(n622), .Y(blockdata[61]) );
  MXI4X1 U1111 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n676), .S1(n649), .Y(n417) );
  MXI4X1 U1112 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n676), .S1(n646), .Y(n416) );
  MXI2X1 U1113 ( .A(n352), .B(n353), .S0(n621), .Y(blockdata[93]) );
  MXI4X1 U1114 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n671), .S1(n640), .Y(n353) );
  MXI4X1 U1115 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n671), .S1(n640), .Y(n352) );
  MXI2X1 U1116 ( .A(n414), .B(n415), .S0(n624), .Y(blockdata[62]) );
  MXI4X1 U1117 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n676), .S1(n645), .Y(n415) );
  MXI4X1 U1118 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n676), .S1(n648), .Y(n414) );
  MXI2X1 U1119 ( .A(n350), .B(n351), .S0(n621), .Y(blockdata[94]) );
  MXI4X1 U1120 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), 
        .D(\block[7][94] ), .S0(n671), .S1(n640), .Y(n351) );
  MXI4X1 U1121 ( .A(\block[0][94] ), .B(\block[1][94] ), .C(\block[2][94] ), 
        .D(\block[3][94] ), .S0(n671), .S1(n640), .Y(n350) );
  MXI2X1 U1122 ( .A(n412), .B(n413), .S0(n621), .Y(blockdata[63]) );
  MXI4X1 U1123 ( .A(\block[4][63] ), .B(\block[5][63] ), .C(\block[6][63] ), 
        .D(\block[7][63] ), .S0(n676), .S1(n645), .Y(n413) );
  MXI4X1 U1124 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n676), .S1(n645), .Y(n412) );
  MXI2X1 U1125 ( .A(n348), .B(n349), .S0(n621), .Y(blockdata[95]) );
  MXI4X1 U1126 ( .A(\block[4][95] ), .B(\block[5][95] ), .C(\block[6][95] ), 
        .D(\block[7][95] ), .S0(n671), .S1(n640), .Y(n349) );
  MXI4X1 U1127 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n671), .S1(n640), .Y(n348) );
  MXI2X1 U1128 ( .A(n346), .B(n347), .S0(n621), .Y(blockdata[96]) );
  MXI4X1 U1129 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n670), .S1(n640), .Y(n347) );
  MXI4X1 U1130 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n671), .S1(n640), .Y(n346) );
  MXI2X1 U1131 ( .A(n344), .B(n345), .S0(n621), .Y(blockdata[97]) );
  MXI4X1 U1132 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n670), .S1(n640), .Y(n345) );
  MXI4X1 U1133 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n670), .S1(n640), .Y(n344) );
  MXI2X1 U1134 ( .A(n342), .B(n343), .S0(n621), .Y(blockdata[98]) );
  MXI4X1 U1135 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n670), .S1(n640), .Y(n343) );
  MXI4X1 U1136 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n670), .S1(n640), .Y(n342) );
  MXI2X1 U1137 ( .A(n340), .B(n341), .S0(n621), .Y(blockdata[99]) );
  MXI4X1 U1138 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n670), .S1(n639), .Y(n341) );
  MXI4X1 U1139 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n670), .S1(n639), .Y(n340) );
  MXI2X1 U1140 ( .A(n338), .B(n339), .S0(n621), .Y(blockdata[100]) );
  MXI4X1 U1141 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n670), .S1(n639), .Y(n339) );
  MXI4X1 U1142 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n670), .S1(n639), .Y(n338) );
  MXI4X1 U1143 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n674), .S1(n653), .Y(n565) );
  MXI2X1 U1144 ( .A(n336), .B(n337), .S0(n621), .Y(blockdata[101]) );
  MXI4X1 U1145 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n670), .S1(n639), .Y(n337) );
  MXI4X1 U1146 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n670), .S1(n639), .Y(n336) );
  MXI4X1 U1147 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n673), .S1(n653), .Y(n563) );
  MXI4X1 U1148 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n680), .S1(n653), .Y(n562) );
  MXI2X1 U1149 ( .A(n334), .B(n335), .S0(n621), .Y(blockdata[102]) );
  MXI4X1 U1150 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n670), .S1(n639), .Y(n335) );
  MXI4X1 U1151 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n670), .S1(n639), .Y(n334) );
  MXI4X1 U1152 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n669), .S1(n653), .Y(n561) );
  MXI4X1 U1153 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n681), .S1(n653), .Y(n560) );
  MXI2X1 U1154 ( .A(n332), .B(n333), .S0(n621), .Y(blockdata[103]) );
  MXI4X1 U1155 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n669), .S1(n639), .Y(n333) );
  MXI4X1 U1156 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n669), .S1(n639), .Y(n332) );
  MXI4X1 U1157 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n667), .S1(n653), .Y(n559) );
  MXI4X1 U1158 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n667), .S1(n653), .Y(n558) );
  MXI2X1 U1159 ( .A(n330), .B(n331), .S0(n621), .Y(blockdata[104]) );
  MXI4X1 U1160 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n669), .S1(n639), .Y(n331) );
  MXI4X1 U1161 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n669), .S1(n639), .Y(n330) );
  MXI2X1 U1162 ( .A(n556), .B(n557), .S0(n626), .Y(blockdata[9]) );
  MXI4X1 U1163 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n678), .S1(n652), .Y(n557) );
  MXI4X1 U1164 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n681), .S1(n652), .Y(n556) );
  MXI2X1 U1165 ( .A(n328), .B(n329), .S0(n620), .Y(blockdata[105]) );
  MXI4X1 U1166 ( .A(\block[4][105] ), .B(\block[5][105] ), .C(\block[6][105] ), 
        .D(\block[7][105] ), .S0(n669), .S1(n641), .Y(n329) );
  MXI4X1 U1167 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n669), .S1(n649), .Y(n328) );
  MXI2X1 U1168 ( .A(n554), .B(n555), .S0(n626), .Y(blockdata[10]) );
  MXI4X1 U1169 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n676), .S1(n652), .Y(n555) );
  MXI4X1 U1170 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n675), .S1(n652), .Y(n554) );
  MXI2X1 U1171 ( .A(n326), .B(n327), .S0(n623), .Y(blockdata[106]) );
  MXI4X1 U1172 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n669), .S1(n642), .Y(n327) );
  MXI4X1 U1173 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n669), .S1(n640), .Y(n326) );
  MXI2X1 U1174 ( .A(n552), .B(n553), .S0(n626), .Y(blockdata[11]) );
  MXI4X1 U1175 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n680), .S1(n652), .Y(n553) );
  MXI4X1 U1176 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n670), .S1(n652), .Y(n552) );
  MXI2X1 U1177 ( .A(n324), .B(n325), .S0(n624), .Y(blockdata[107]) );
  MXI4X1 U1178 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n669), .S1(n644), .Y(n325) );
  MXI4X1 U1179 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n669), .S1(n643), .Y(n324) );
  MXI2X1 U1180 ( .A(n550), .B(n551), .S0(n626), .Y(blockdata[12]) );
  MXI4X1 U1181 ( .A(\block[4][12] ), .B(\block[5][12] ), .C(\block[6][12] ), 
        .D(\block[7][12] ), .S0(n681), .S1(n652), .Y(n551) );
  MXI4X1 U1182 ( .A(\block[0][12] ), .B(\block[1][12] ), .C(\block[2][12] ), 
        .D(\block[3][12] ), .S0(n681), .S1(n652), .Y(n550) );
  MXI2X1 U1183 ( .A(n322), .B(n323), .S0(n625), .Y(blockdata[108]) );
  MXI4X1 U1184 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n669), .S1(n639), .Y(n323) );
  MXI4X1 U1185 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n669), .S1(n645), .Y(n322) );
  MXI2X1 U1186 ( .A(n548), .B(n549), .S0(n626), .Y(blockdata[13]) );
  MXI4X1 U1187 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n681), .S1(n652), .Y(n549) );
  MXI4X1 U1188 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n681), .S1(n652), .Y(n548) );
  MXI2X1 U1189 ( .A(n320), .B(n321), .S0(n623), .Y(blockdata[109]) );
  MXI4X1 U1190 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n668), .S1(n642), .Y(n321) );
  MXI4X1 U1191 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n669), .S1(n647), .Y(n320) );
  MXI2X1 U1192 ( .A(n546), .B(n547), .S0(n626), .Y(blockdata[14]) );
  MXI4X1 U1193 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n681), .S1(n652), .Y(n547) );
  MXI4X1 U1194 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n681), .S1(n652), .Y(n546) );
  MXI2X1 U1195 ( .A(n318), .B(n319), .S0(n624), .Y(blockdata[110]) );
  MXI4X1 U1196 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n668), .S1(n644), .Y(n319) );
  MXI4X1 U1197 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n668), .S1(n646), .Y(n318) );
  MXI2X1 U1198 ( .A(n544), .B(n545), .S0(n626), .Y(blockdata[15]) );
  MXI4X1 U1199 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n681), .S1(n651), .Y(n545) );
  MXI4X1 U1200 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n681), .S1(n651), .Y(n544) );
  MXI2X1 U1201 ( .A(n316), .B(n317), .S0(n624), .Y(blockdata[111]) );
  MXI4X1 U1202 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n668), .S1(n641), .Y(n317) );
  MXI4X1 U1203 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n668), .S1(n643), .Y(n316) );
  MXI2X1 U1204 ( .A(n542), .B(n543), .S0(n626), .Y(blockdata[16]) );
  MXI4X1 U1205 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n681), .S1(n651), .Y(n543) );
  MXI4X1 U1206 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n681), .S1(n651), .Y(n542) );
  MXI2X1 U1207 ( .A(n314), .B(n315), .S0(n624), .Y(blockdata[112]) );
  MXI4X1 U1208 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n668), .S1(n640), .Y(n315) );
  MXI4X1 U1209 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n668), .S1(n641), .Y(n314) );
  MXI2X1 U1210 ( .A(n540), .B(n541), .S0(n626), .Y(blockdata[17]) );
  MXI4X1 U1211 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n681), .S1(n651), .Y(n541) );
  MXI4X1 U1212 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n681), .S1(n651), .Y(n540) );
  MXI2X1 U1213 ( .A(n312), .B(n313), .S0(n621), .Y(blockdata[113]) );
  MXI4X1 U1214 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n668), .S1(n641), .Y(n313) );
  MXI4X1 U1215 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n668), .S1(n642), .Y(n312) );
  MXI2X1 U1216 ( .A(n538), .B(n539), .S0(n626), .Y(blockdata[18]) );
  MXI4X1 U1217 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n680), .S1(n651), .Y(n539) );
  MXI4X1 U1218 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n681), .S1(n651), .Y(n538) );
  MXI2X1 U1219 ( .A(n310), .B(n311), .S0(n626), .Y(blockdata[114]) );
  MXI4X1 U1220 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n668), .S1(n640), .Y(n311) );
  MXI4X1 U1221 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n668), .S1(n644), .Y(n310) );
  MXI2X1 U1222 ( .A(n536), .B(n537), .S0(n626), .Y(blockdata[19]) );
  MXI4X1 U1223 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n680), .S1(n651), .Y(n537) );
  MXI4X1 U1224 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n680), .S1(n651), .Y(n536) );
  MXI2X1 U1225 ( .A(n308), .B(n309), .S0(n621), .Y(blockdata[115]) );
  MXI4X1 U1226 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n668), .S1(n641), .Y(n309) );
  MXI4X1 U1227 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n668), .S1(n640), .Y(n308) );
  MXI2X1 U1228 ( .A(n534), .B(n535), .S0(n626), .Y(blockdata[20]) );
  MXI4X1 U1229 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n680), .S1(n651), .Y(n535) );
  MXI4X1 U1230 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n680), .S1(n651), .Y(n534) );
  MXI2X1 U1231 ( .A(n306), .B(n307), .S0(n626), .Y(blockdata[116]) );
  MXI4X1 U1232 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n667), .S1(n640), .Y(n307) );
  MXI4X1 U1233 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n667), .S1(n643), .Y(n306) );
  MXI2X1 U1234 ( .A(n532), .B(n533), .S0(n625), .Y(blockdata[21]) );
  MXI4X1 U1235 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n680), .S1(n652), .Y(n533) );
  MXI4X1 U1236 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n680), .S1(n652), .Y(n532) );
  MXI2X1 U1237 ( .A(n304), .B(n305), .S0(n620), .Y(blockdata[117]) );
  MXI4X1 U1238 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n667), .S1(n638), .Y(n305) );
  MXI4X1 U1239 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n667), .S1(n638), .Y(n304) );
  MXI2X1 U1240 ( .A(n530), .B(n531), .S0(n625), .Y(blockdata[22]) );
  MXI4X1 U1241 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n680), .S1(n651), .Y(n531) );
  MXI4X1 U1242 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n680), .S1(n651), .Y(n530) );
  MXI2X1 U1243 ( .A(n302), .B(n303), .S0(n622), .Y(blockdata[118]) );
  MXI4X1 U1244 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n667), .S1(n638), .Y(n303) );
  MXI4X1 U1245 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n667), .S1(n638), .Y(n302) );
  MXI2X1 U1246 ( .A(n528), .B(n529), .S0(n625), .Y(blockdata[23]) );
  MXI4X1 U1247 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n680), .S1(n652), .Y(n529) );
  MXI4X1 U1248 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n680), .S1(n650), .Y(n528) );
  MXI2X1 U1249 ( .A(n300), .B(n301), .S0(n620), .Y(blockdata[119]) );
  MXI4X1 U1250 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n667), .S1(n638), .Y(n301) );
  MXI4X1 U1251 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n667), .S1(n638), .Y(n300) );
  MXI2X1 U1252 ( .A(n526), .B(n527), .S0(n625), .Y(blockdata[24]) );
  MXI4X1 U1253 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n680), .S1(n652), .Y(n527) );
  MXI4X1 U1254 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n680), .S1(n652), .Y(n526) );
  MXI2X1 U1255 ( .A(n298), .B(n299), .S0(n621), .Y(blockdata[120]) );
  MXI4X1 U1256 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n667), .S1(n638), .Y(n299) );
  MXI4X1 U1257 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n667), .S1(n638), .Y(n298) );
  MXI2X1 U1258 ( .A(n524), .B(n525), .S0(n625), .Y(blockdata[25]) );
  MXI4X1 U1259 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n676), .S1(n651), .Y(n525) );
  MXI4X1 U1260 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n668), .S1(n651), .Y(n524) );
  MXI2X1 U1261 ( .A(n296), .B(n297), .S0(n620), .Y(blockdata[121]) );
  MXI4X1 U1262 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n667), .S1(n638), .Y(n297) );
  MXI4X1 U1263 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n667), .S1(n638), .Y(n296) );
  MXI2X1 U1264 ( .A(n522), .B(n523), .S0(n625), .Y(blockdata[26]) );
  MXI4X1 U1265 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n671), .S1(n651), .Y(n523) );
  MXI4X1 U1266 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n679), .S1(n652), .Y(n522) );
  MXI2X1 U1267 ( .A(n294), .B(n295), .S0(n620), .Y(blockdata[122]) );
  MXI4X1 U1268 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n667), .S1(n638), .Y(n295) );
  MXI4X1 U1269 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n667), .S1(n638), .Y(n294) );
  MXI2X1 U1270 ( .A(n520), .B(n521), .S0(n625), .Y(blockdata[27]) );
  MXI4X1 U1271 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n672), .S1(n650), .Y(n521) );
  MXI4X1 U1272 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n678), .S1(n650), .Y(n520) );
  MXI2X1 U1273 ( .A(n518), .B(n519), .S0(n625), .Y(blockdata[28]) );
  MXI4X1 U1274 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n673), .S1(n650), .Y(n519) );
  MXI4X1 U1275 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n684), .S1(n650), .Y(n518) );
  MXI2X1 U1276 ( .A(n516), .B(n517), .S0(n625), .Y(blockdata[29]) );
  MXI4X1 U1277 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n675), .S1(n650), .Y(n517) );
  MXI4X1 U1278 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n684), .S1(n650), .Y(n516) );
  MXI2X1 U1279 ( .A(n514), .B(n515), .S0(n625), .Y(blockdata[30]) );
  MXI4X1 U1280 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n677), .S1(n650), .Y(n515) );
  MXI4X1 U1281 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n684), .S1(n650), .Y(n514) );
  MXI2X1 U1282 ( .A(n512), .B(n513), .S0(n625), .Y(blockdata[31]) );
  MXI4X1 U1283 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n681), .S1(n650), .Y(n513) );
  MXI4X1 U1284 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n684), .S1(n650), .Y(n512) );
  MXI2X1 U1285 ( .A(n471), .B(n1052), .S0(n250), .Y(n487) );
  MXI2X1 U1286 ( .A(n472), .B(n1052), .S0(n244), .Y(n488) );
  MXI2X1 U1287 ( .A(n473), .B(n1052), .S0(n251), .Y(n489) );
  MXI2X1 U1288 ( .A(n474), .B(n1052), .S0(n245), .Y(n490) );
  MXI2X1 U1289 ( .A(n475), .B(n1052), .S0(n253), .Y(n491) );
  MXI2X1 U1290 ( .A(n476), .B(n1052), .S0(n247), .Y(n492) );
  MXI2X1 U1291 ( .A(n477), .B(n1052), .S0(n252), .Y(n493) );
  MXI2X1 U1292 ( .A(n478), .B(n1052), .S0(n246), .Y(n494) );
  OAI221XL U1293 ( .A0(n729), .A1(n1064), .B0(n726), .B1(n1063), .C0(n1062), 
        .Y(proc_rdata[0]) );
  OA22X1 U1294 ( .A0(n725), .A1(n1061), .B0(n722), .B1(n1060), .Y(n1062) );
  OAI221XL U1295 ( .A0(n729), .A1(n1069), .B0(n726), .B1(n1068), .C0(n1067), 
        .Y(proc_rdata[1]) );
  OA22X1 U1296 ( .A0(n725), .A1(n1066), .B0(n722), .B1(n1065), .Y(n1067) );
  OAI221XL U1297 ( .A0(n729), .A1(n1074), .B0(n726), .B1(n1073), .C0(n1072), 
        .Y(proc_rdata[2]) );
  OA22X1 U1298 ( .A0(n725), .A1(n1071), .B0(n722), .B1(n1070), .Y(n1072) );
  OAI221XL U1299 ( .A0(n729), .A1(n1079), .B0(n726), .B1(n1078), .C0(n1077), 
        .Y(proc_rdata[3]) );
  OA22X1 U1300 ( .A0(n725), .A1(n1076), .B0(n722), .B1(n1075), .Y(n1077) );
  OAI221XL U1301 ( .A0(n729), .A1(n1084), .B0(n726), .B1(n1083), .C0(n1082), 
        .Y(proc_rdata[4]) );
  OA22X1 U1302 ( .A0(n725), .A1(n1081), .B0(n722), .B1(n1080), .Y(n1082) );
  OAI221XL U1303 ( .A0(n729), .A1(n1089), .B0(n726), .B1(n1088), .C0(n1087), 
        .Y(proc_rdata[5]) );
  OA22X1 U1304 ( .A0(n725), .A1(n1086), .B0(n722), .B1(n1085), .Y(n1087) );
  OAI221XL U1305 ( .A0(n729), .A1(n1094), .B0(n726), .B1(n1093), .C0(n1092), 
        .Y(proc_rdata[6]) );
  OA22X1 U1306 ( .A0(n725), .A1(n1091), .B0(n722), .B1(n1090), .Y(n1092) );
  OAI221XL U1307 ( .A0(n729), .A1(n1099), .B0(n726), .B1(n1098), .C0(n1097), 
        .Y(proc_rdata[7]) );
  OA22X1 U1308 ( .A0(n725), .A1(n1096), .B0(n722), .B1(n1095), .Y(n1097) );
  OAI221XL U1309 ( .A0(n729), .A1(n1104), .B0(n726), .B1(n1103), .C0(n1102), 
        .Y(proc_rdata[8]) );
  OA22X1 U1310 ( .A0(n725), .A1(n1101), .B0(n722), .B1(n1100), .Y(n1102) );
  OAI221XL U1311 ( .A0(n729), .A1(n1109), .B0(n726), .B1(n1108), .C0(n1107), 
        .Y(proc_rdata[9]) );
  OA22X1 U1312 ( .A0(n725), .A1(n1106), .B0(n722), .B1(n1105), .Y(n1107) );
  OAI221XL U1313 ( .A0(n729), .A1(n1114), .B0(n726), .B1(n1113), .C0(n1112), 
        .Y(proc_rdata[10]) );
  OA22X1 U1314 ( .A0(n725), .A1(n1111), .B0(n722), .B1(n1110), .Y(n1112) );
  OAI221XL U1315 ( .A0(n729), .A1(n1119), .B0(n726), .B1(n1118), .C0(n1117), 
        .Y(proc_rdata[11]) );
  OA22X1 U1316 ( .A0(n725), .A1(n1116), .B0(n722), .B1(n1115), .Y(n1117) );
  OAI221XL U1317 ( .A0(n730), .A1(n1124), .B0(n727), .B1(n1123), .C0(n1122), 
        .Y(proc_rdata[12]) );
  OA22X1 U1318 ( .A0(n724), .A1(n1121), .B0(n723), .B1(n1120), .Y(n1122) );
  OAI221XL U1319 ( .A0(n730), .A1(n1129), .B0(n727), .B1(n1128), .C0(n1127), 
        .Y(proc_rdata[13]) );
  OA22X1 U1320 ( .A0(n724), .A1(n1126), .B0(n723), .B1(n1125), .Y(n1127) );
  OAI221XL U1321 ( .A0(n730), .A1(n1134), .B0(n727), .B1(n1133), .C0(n1132), 
        .Y(proc_rdata[14]) );
  OA22X1 U1322 ( .A0(n724), .A1(n1131), .B0(n723), .B1(n1130), .Y(n1132) );
  OAI221XL U1323 ( .A0(n730), .A1(n1139), .B0(n727), .B1(n1138), .C0(n1137), 
        .Y(proc_rdata[15]) );
  OA22X1 U1324 ( .A0(n724), .A1(n1136), .B0(n723), .B1(n1135), .Y(n1137) );
  OAI221XL U1325 ( .A0(n730), .A1(n1144), .B0(n727), .B1(n1143), .C0(n1142), 
        .Y(proc_rdata[16]) );
  OA22X1 U1326 ( .A0(n724), .A1(n1141), .B0(n723), .B1(n1140), .Y(n1142) );
  OAI221XL U1327 ( .A0(n730), .A1(n1149), .B0(n727), .B1(n1148), .C0(n1147), 
        .Y(proc_rdata[17]) );
  OA22X1 U1328 ( .A0(n725), .A1(n1146), .B0(n723), .B1(n1145), .Y(n1147) );
  OAI221XL U1329 ( .A0(n730), .A1(n1154), .B0(n727), .B1(n1153), .C0(n1152), 
        .Y(proc_rdata[18]) );
  OA22X1 U1330 ( .A0(n724), .A1(n1151), .B0(n723), .B1(n1150), .Y(n1152) );
  OAI221XL U1331 ( .A0(n730), .A1(n1159), .B0(n727), .B1(n1158), .C0(n1157), 
        .Y(proc_rdata[19]) );
  OA22X1 U1332 ( .A0(n725), .A1(n1156), .B0(n723), .B1(n1155), .Y(n1157) );
  OAI221XL U1333 ( .A0(n730), .A1(n1164), .B0(n727), .B1(n1163), .C0(n1162), 
        .Y(proc_rdata[20]) );
  OA22X1 U1334 ( .A0(n1218), .A1(n1161), .B0(n723), .B1(n1160), .Y(n1162) );
  OAI221XL U1335 ( .A0(n730), .A1(n1169), .B0(n727), .B1(n1168), .C0(n1167), 
        .Y(proc_rdata[21]) );
  OA22X1 U1336 ( .A0(n1218), .A1(n1166), .B0(n723), .B1(n1165), .Y(n1167) );
  OAI221XL U1337 ( .A0(n730), .A1(n1174), .B0(n727), .B1(n1173), .C0(n1172), 
        .Y(proc_rdata[22]) );
  OA22X1 U1338 ( .A0(n1218), .A1(n1171), .B0(n723), .B1(n1170), .Y(n1172) );
  OAI221XL U1339 ( .A0(n730), .A1(n1179), .B0(n727), .B1(n1178), .C0(n1177), 
        .Y(proc_rdata[23]) );
  OA22X1 U1340 ( .A0(n1218), .A1(n1176), .B0(n723), .B1(n1175), .Y(n1177) );
  OAI221XL U1341 ( .A0(n728), .A1(n1184), .B0(n726), .B1(n1183), .C0(n1182), 
        .Y(proc_rdata[24]) );
  OA22X1 U1342 ( .A0(n724), .A1(n1181), .B0(n721), .B1(n1180), .Y(n1182) );
  OAI221XL U1343 ( .A0(n728), .A1(n1189), .B0(n727), .B1(n1188), .C0(n1187), 
        .Y(proc_rdata[25]) );
  OA22X1 U1344 ( .A0(n724), .A1(n1186), .B0(n721), .B1(n1185), .Y(n1187) );
  OAI221XL U1345 ( .A0(n728), .A1(n1194), .B0(n726), .B1(n1193), .C0(n1192), 
        .Y(proc_rdata[26]) );
  OA22X1 U1346 ( .A0(n724), .A1(n1191), .B0(n721), .B1(n1190), .Y(n1192) );
  OAI221XL U1347 ( .A0(n728), .A1(n1199), .B0(n727), .B1(n1198), .C0(n1197), 
        .Y(proc_rdata[27]) );
  OA22X1 U1348 ( .A0(n724), .A1(n1196), .B0(n721), .B1(n1195), .Y(n1197) );
  OAI221XL U1349 ( .A0(n728), .A1(n1204), .B0(n1221), .B1(n1203), .C0(n1202), 
        .Y(proc_rdata[28]) );
  OA22X1 U1350 ( .A0(n724), .A1(n1201), .B0(n721), .B1(n1200), .Y(n1202) );
  OAI221XL U1351 ( .A0(n1223), .A1(n1209), .B0(n1221), .B1(n1208), .C0(n1207), 
        .Y(proc_rdata[29]) );
  OA22X1 U1352 ( .A0(n724), .A1(n1206), .B0(n721), .B1(n1205), .Y(n1207) );
  OAI221XL U1353 ( .A0(n1223), .A1(n1214), .B0(n1221), .B1(n1213), .C0(n1212), 
        .Y(proc_rdata[30]) );
  OA22X1 U1354 ( .A0(n724), .A1(n1211), .B0(n721), .B1(n1210), .Y(n1212) );
  OAI221XL U1355 ( .A0(n1223), .A1(n1222), .B0(n1221), .B1(n1220), .C0(n1219), 
        .Y(proc_rdata[31]) );
  OA22X1 U1356 ( .A0(n724), .A1(n1217), .B0(n721), .B1(n1215), .Y(n1219) );
  INVX1 U1357 ( .A(proc_wdata[0]), .Y(n1001) );
  INVX1 U1358 ( .A(proc_wdata[1]), .Y(n999) );
  INVX1 U1359 ( .A(proc_wdata[2]), .Y(n997) );
  INVX1 U1360 ( .A(proc_wdata[3]), .Y(n995) );
  INVX1 U1361 ( .A(proc_wdata[4]), .Y(n993) );
  INVX1 U1362 ( .A(proc_wdata[5]), .Y(n991) );
  INVX1 U1363 ( .A(proc_wdata[6]), .Y(n989) );
  INVX1 U1364 ( .A(proc_wdata[7]), .Y(n987) );
  INVX1 U1365 ( .A(proc_wdata[8]), .Y(n985) );
  INVX1 U1366 ( .A(proc_wdata[9]), .Y(n983) );
  INVX1 U1367 ( .A(proc_wdata[10]), .Y(n981) );
  INVX1 U1368 ( .A(proc_wdata[11]), .Y(n979) );
  INVX1 U1369 ( .A(proc_wdata[12]), .Y(n977) );
  INVX1 U1370 ( .A(proc_wdata[13]), .Y(n975) );
  INVX1 U1371 ( .A(proc_wdata[14]), .Y(n973) );
  INVX1 U1372 ( .A(proc_wdata[15]), .Y(n971) );
  INVX1 U1373 ( .A(proc_wdata[16]), .Y(n969) );
  INVX1 U1374 ( .A(proc_wdata[17]), .Y(n967) );
  INVX1 U1375 ( .A(proc_wdata[18]), .Y(n965) );
  INVX1 U1376 ( .A(proc_wdata[19]), .Y(n963) );
  INVX1 U1377 ( .A(proc_wdata[20]), .Y(n961) );
  INVX1 U1378 ( .A(proc_wdata[21]), .Y(n959) );
  INVX1 U1379 ( .A(proc_wdata[22]), .Y(n957) );
  INVX1 U1380 ( .A(proc_wdata[23]), .Y(n955) );
  INVX1 U1381 ( .A(proc_wdata[24]), .Y(n953) );
  INVX1 U1382 ( .A(proc_wdata[25]), .Y(n951) );
  INVX1 U1383 ( .A(proc_wdata[26]), .Y(n949) );
  INVX1 U1384 ( .A(proc_wdata[27]), .Y(n947) );
  INVX1 U1385 ( .A(proc_wdata[28]), .Y(n945) );
  INVX1 U1386 ( .A(proc_wdata[29]), .Y(n943) );
  INVX1 U1387 ( .A(proc_wdata[30]), .Y(n941) );
  INVX1 U1388 ( .A(proc_wdata[31]), .Y(n939) );
  MXI2X1 U1389 ( .A(n479), .B(n77), .S0(n250), .Y(n495) );
  MXI2X1 U1390 ( .A(n480), .B(n77), .S0(n244), .Y(n496) );
  MXI2X1 U1391 ( .A(n481), .B(n77), .S0(n251), .Y(n497) );
  MXI2X1 U1392 ( .A(n482), .B(n77), .S0(n245), .Y(n498) );
  MXI2X1 U1393 ( .A(n483), .B(n77), .S0(n253), .Y(n499) );
  MXI2X1 U1394 ( .A(n484), .B(n77), .S0(n247), .Y(n500) );
  MXI2X1 U1395 ( .A(n485), .B(n77), .S0(n252), .Y(n501) );
  MXI2X1 U1396 ( .A(n486), .B(n77), .S0(n246), .Y(n503) );
  MXI2X1 U1397 ( .A(n292), .B(n293), .S0(n620), .Y(blockdata[123]) );
  MXI4X1 U1398 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n670), .S1(n651), .Y(n293) );
  MXI4X1 U1399 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n669), .S1(n652), .Y(n292) );
  MXI2X1 U1400 ( .A(n290), .B(n291), .S0(n620), .Y(blockdata[124]) );
  MXI4X1 U1401 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n680), .S1(n651), .Y(n291) );
  MXI4X1 U1402 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n668), .S1(n638), .Y(n290) );
  MXI2X1 U1403 ( .A(n288), .B(n289), .S0(n620), .Y(blockdata[125]) );
  MXI4X1 U1404 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n670), .S1(n652), .Y(n289) );
  MXI4X1 U1405 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n671), .S1(n638), .Y(n288) );
  MXI2X1 U1406 ( .A(n286), .B(n287), .S0(n626), .Y(blockdata[126]) );
  MXI4X1 U1407 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n674), .S1(n651), .Y(n287) );
  MXI4X1 U1408 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n672), .S1(n638), .Y(n286) );
  MXI2X1 U1409 ( .A(n284), .B(n285), .S0(n627), .Y(blockdata[127]) );
  MXI4X1 U1410 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n677), .S1(n638), .Y(n285) );
  MXI4X1 U1411 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n679), .S1(n638), .Y(n284) );
  CLKINVX1 U1412 ( .A(mem_ready), .Y(n1053) );
  INVXL U1413 ( .A(proc_addr[23]), .Y(n1018) );
  INVXL U1414 ( .A(proc_addr[6]), .Y(n1048) );
  INVXL U1415 ( .A(proc_addr[12]), .Y(n1040) );
  INVXL U1416 ( .A(proc_addr[11]), .Y(n1042) );
  INVXL U1417 ( .A(proc_addr[8]), .Y(n1046) );
  INVXL U1418 ( .A(proc_addr[26]), .Y(n1012) );
  INVXL U1419 ( .A(proc_addr[0]), .Y(n1225) );
  INVXL U1420 ( .A(proc_addr[1]), .Y(n1224) );
  INVXL U1421 ( .A(proc_addr[20]), .Y(n1024) );
  OAI21XL U1422 ( .A0(n1053), .A1(n1003), .B0(dirty), .Y(n1005) );
  NAND3BXL U1423 ( .AN(n835), .B(proc_write), .C(n832), .Y(n1004) );
  CLKINVX3 U1424 ( .A(n833), .Y(n868) );
  OAI221X2 U1425 ( .A0(n687), .A1(n1220), .B0(n939), .B1(n691), .C0(n836), .Y(
        block_next[127]) );
  OAI221X2 U1426 ( .A0(n687), .A1(n1213), .B0(n941), .B1(n691), .C0(n837), .Y(
        block_next[126]) );
  OAI221X2 U1427 ( .A0(n687), .A1(n1208), .B0(n943), .B1(n691), .C0(n838), .Y(
        block_next[125]) );
  OAI221X2 U1428 ( .A0(n687), .A1(n1203), .B0(n945), .B1(n691), .C0(n839), .Y(
        block_next[124]) );
  OAI221X2 U1429 ( .A0(n687), .A1(n1198), .B0(n947), .B1(n691), .C0(n840), .Y(
        block_next[123]) );
  OAI221X2 U1430 ( .A0(n687), .A1(n1193), .B0(n949), .B1(n691), .C0(n841), .Y(
        block_next[122]) );
  OAI221X2 U1431 ( .A0(n687), .A1(n1178), .B0(n955), .B1(n691), .C0(n844), .Y(
        block_next[119]) );
  OAI221X2 U1432 ( .A0(n687), .A1(n1173), .B0(n957), .B1(n691), .C0(n845), .Y(
        block_next[118]) );
  OAI221X2 U1433 ( .A0(n687), .A1(n1168), .B0(n959), .B1(n691), .C0(n846), .Y(
        block_next[117]) );
  OAI221X2 U1434 ( .A0(n687), .A1(n1163), .B0(n961), .B1(n691), .C0(n847), .Y(
        block_next[116]) );
  OAI221X2 U1435 ( .A0(n688), .A1(n1158), .B0(n963), .B1(n692), .C0(n848), .Y(
        block_next[115]) );
  OAI221X2 U1436 ( .A0(n688), .A1(n1153), .B0(n965), .B1(n692), .C0(n849), .Y(
        block_next[114]) );
  OAI221X2 U1437 ( .A0(n688), .A1(n1148), .B0(n967), .B1(n692), .C0(n850), .Y(
        block_next[113]) );
  OAI221X2 U1438 ( .A0(n688), .A1(n1143), .B0(n969), .B1(n692), .C0(n851), .Y(
        block_next[112]) );
  OAI221X2 U1439 ( .A0(n688), .A1(n1138), .B0(n971), .B1(n692), .C0(n852), .Y(
        block_next[111]) );
  OAI221X2 U1440 ( .A0(n688), .A1(n1133), .B0(n973), .B1(n692), .C0(n853), .Y(
        block_next[110]) );
  OAI221X2 U1441 ( .A0(n688), .A1(n1128), .B0(n975), .B1(n692), .C0(n854), .Y(
        block_next[109]) );
  OAI221X2 U1442 ( .A0(n688), .A1(n1123), .B0(n977), .B1(n692), .C0(n855), .Y(
        block_next[108]) );
  OAI221X2 U1443 ( .A0(n688), .A1(n1118), .B0(n979), .B1(n692), .C0(n856), .Y(
        block_next[107]) );
  OAI221X2 U1444 ( .A0(n688), .A1(n1113), .B0(n981), .B1(n692), .C0(n857), .Y(
        block_next[106]) );
  OAI221X2 U1445 ( .A0(n688), .A1(n1108), .B0(n983), .B1(n692), .C0(n858), .Y(
        block_next[105]) );
  OAI221X2 U1446 ( .A0(n689), .A1(n1098), .B0(n987), .B1(n690), .C0(n860), .Y(
        block_next[103]) );
  OAI221X2 U1447 ( .A0(n689), .A1(n1093), .B0(n989), .B1(n690), .C0(n861), .Y(
        block_next[102]) );
  OAI221X2 U1448 ( .A0(n689), .A1(n1088), .B0(n991), .B1(n690), .C0(n862), .Y(
        block_next[101]) );
  OAI221X2 U1449 ( .A0(n689), .A1(n1083), .B0(n993), .B1(n690), .C0(n863), .Y(
        block_next[100]) );
  OAI221X2 U1450 ( .A0(n689), .A1(n1078), .B0(n995), .B1(n690), .C0(n864), .Y(
        block_next[99]) );
  OAI221X2 U1451 ( .A0(n689), .A1(n1073), .B0(n997), .B1(n690), .C0(n865), .Y(
        block_next[98]) );
  OAI221X2 U1452 ( .A0(n689), .A1(n1068), .B0(n999), .B1(n691), .C0(n866), .Y(
        block_next[97]) );
  OAI221X2 U1453 ( .A0(n689), .A1(n1063), .B0(n1001), .B1(n692), .C0(n867), 
        .Y(block_next[96]) );
  CLKINVX3 U1454 ( .A(n871), .Y(n904) );
  OAI221X2 U1455 ( .A0(n693), .A1(n1217), .B0(n939), .B1(n697), .C0(n872), .Y(
        block_next[95]) );
  OAI221X2 U1456 ( .A0(n693), .A1(n1211), .B0(n941), .B1(n698), .C0(n873), .Y(
        block_next[94]) );
  OAI221X2 U1457 ( .A0(n693), .A1(n1206), .B0(n943), .B1(n696), .C0(n874), .Y(
        block_next[93]) );
  OAI221X2 U1458 ( .A0(n693), .A1(n1201), .B0(n945), .B1(n696), .C0(n875), .Y(
        block_next[92]) );
  OAI221X2 U1459 ( .A0(n693), .A1(n1196), .B0(n947), .B1(n696), .C0(n876), .Y(
        block_next[91]) );
  OAI221X2 U1460 ( .A0(n693), .A1(n1191), .B0(n949), .B1(n696), .C0(n877), .Y(
        block_next[90]) );
  OAI221X2 U1461 ( .A0(n693), .A1(n1181), .B0(n953), .B1(n696), .C0(n879), .Y(
        block_next[88]) );
  OAI221X2 U1462 ( .A0(n693), .A1(n1176), .B0(n955), .B1(n698), .C0(n880), .Y(
        block_next[87]) );
  OAI221X2 U1463 ( .A0(n693), .A1(n1171), .B0(n957), .B1(n698), .C0(n881), .Y(
        block_next[86]) );
  OAI221X2 U1464 ( .A0(n693), .A1(n1166), .B0(n959), .B1(n698), .C0(n882), .Y(
        block_next[85]) );
  OAI221X2 U1465 ( .A0(n694), .A1(n1156), .B0(n963), .B1(n698), .C0(n884), .Y(
        block_next[83]) );
  OAI221X2 U1466 ( .A0(n694), .A1(n1151), .B0(n965), .B1(n698), .C0(n885), .Y(
        block_next[82]) );
  OAI221X2 U1467 ( .A0(n694), .A1(n1146), .B0(n967), .B1(n698), .C0(n886), .Y(
        block_next[81]) );
  OAI221X2 U1468 ( .A0(n694), .A1(n1141), .B0(n969), .B1(n698), .C0(n887), .Y(
        block_next[80]) );
  OAI221X2 U1469 ( .A0(n694), .A1(n1136), .B0(n971), .B1(n698), .C0(n888), .Y(
        block_next[79]) );
  OAI221X2 U1470 ( .A0(n694), .A1(n1131), .B0(n973), .B1(n698), .C0(n889), .Y(
        block_next[78]) );
  OAI221X2 U1471 ( .A0(n694), .A1(n1126), .B0(n975), .B1(n698), .C0(n890), .Y(
        block_next[77]) );
  OAI221X2 U1472 ( .A0(n694), .A1(n1121), .B0(n977), .B1(n697), .C0(n891), .Y(
        block_next[76]) );
  OAI221X2 U1473 ( .A0(n695), .A1(n1091), .B0(n989), .B1(n697), .C0(n897), .Y(
        block_next[70]) );
  OAI221X2 U1474 ( .A0(n695), .A1(n1086), .B0(n991), .B1(n697), .C0(n898), .Y(
        block_next[69]) );
  OAI221X2 U1475 ( .A0(n695), .A1(n1081), .B0(n993), .B1(n697), .C0(n899), .Y(
        block_next[68]) );
  OAI221X2 U1476 ( .A0(n695), .A1(n1076), .B0(n995), .B1(n697), .C0(n900), .Y(
        block_next[67]) );
  OAI221X2 U1477 ( .A0(n695), .A1(n1071), .B0(n997), .B1(n697), .C0(n901), .Y(
        block_next[66]) );
  OAI221X2 U1478 ( .A0(n699), .A1(n1215), .B0(n939), .B1(n704), .C0(n906), .Y(
        block_next[63]) );
  OAI221X2 U1479 ( .A0(n699), .A1(n1210), .B0(n941), .B1(n704), .C0(n907), .Y(
        block_next[62]) );
  OAI221X2 U1480 ( .A0(n699), .A1(n1205), .B0(n943), .B1(n704), .C0(n908), .Y(
        block_next[61]) );
  OAI221X2 U1481 ( .A0(n699), .A1(n1200), .B0(n945), .B1(n704), .C0(n909), .Y(
        block_next[60]) );
  OAI221X2 U1482 ( .A0(n699), .A1(n1195), .B0(n947), .B1(n704), .C0(n910), .Y(
        block_next[59]) );
  OAI221X2 U1483 ( .A0(n699), .A1(n1190), .B0(n949), .B1(n704), .C0(n911), .Y(
        block_next[58]) );
  OAI221X2 U1484 ( .A0(n699), .A1(n1185), .B0(n951), .B1(n704), .C0(n912), .Y(
        block_next[57]) );
  OAI221X2 U1485 ( .A0(n699), .A1(n1180), .B0(n953), .B1(n704), .C0(n913), .Y(
        block_next[56]) );
  OAI221X2 U1486 ( .A0(n699), .A1(n1175), .B0(n955), .B1(n703), .C0(n914), .Y(
        block_next[55]) );
  OAI221X2 U1487 ( .A0(n699), .A1(n1170), .B0(n957), .B1(n703), .C0(n915), .Y(
        block_next[54]) );
  OAI221X2 U1488 ( .A0(n699), .A1(n1165), .B0(n959), .B1(n703), .C0(n916), .Y(
        block_next[53]) );
  OAI221X2 U1489 ( .A0(n700), .A1(n1155), .B0(n963), .B1(n703), .C0(n918), .Y(
        block_next[51]) );
  OAI221X2 U1490 ( .A0(n700), .A1(n1150), .B0(n965), .B1(n703), .C0(n919), .Y(
        block_next[50]) );
  OAI221X2 U1491 ( .A0(n700), .A1(n1145), .B0(n967), .B1(n703), .C0(n920), .Y(
        block_next[49]) );
  OAI221X2 U1492 ( .A0(n700), .A1(n1140), .B0(n969), .B1(n703), .C0(n921), .Y(
        block_next[48]) );
  OAI221X2 U1493 ( .A0(n700), .A1(n1135), .B0(n971), .B1(n703), .C0(n922), .Y(
        block_next[47]) );
  OAI221X2 U1494 ( .A0(n700), .A1(n1130), .B0(n973), .B1(n703), .C0(n923), .Y(
        block_next[46]) );
  OAI221X2 U1495 ( .A0(n700), .A1(n1125), .B0(n975), .B1(n703), .C0(n924), .Y(
        block_next[45]) );
  OAI221X2 U1496 ( .A0(n700), .A1(n1120), .B0(n977), .B1(n702), .C0(n925), .Y(
        block_next[44]) );
  OAI221X2 U1497 ( .A0(n700), .A1(n1115), .B0(n979), .B1(n702), .C0(n926), .Y(
        block_next[43]) );
  OAI221X2 U1498 ( .A0(n700), .A1(n1110), .B0(n981), .B1(n702), .C0(n927), .Y(
        block_next[42]) );
  OAI221X2 U1499 ( .A0(n700), .A1(n1105), .B0(n983), .B1(n702), .C0(n928), .Y(
        block_next[41]) );
  OAI221X2 U1500 ( .A0(n701), .A1(n1095), .B0(n987), .B1(n703), .C0(n930), .Y(
        block_next[39]) );
  OAI221X2 U1501 ( .A0(n701), .A1(n1090), .B0(n989), .B1(n702), .C0(n931), .Y(
        block_next[38]) );
  OAI221X2 U1502 ( .A0(n701), .A1(n1085), .B0(n991), .B1(n702), .C0(n932), .Y(
        block_next[37]) );
  OAI221X2 U1503 ( .A0(n701), .A1(n1080), .B0(n993), .B1(n702), .C0(n933), .Y(
        block_next[36]) );
  OAI221X2 U1504 ( .A0(n701), .A1(n1075), .B0(n995), .B1(n702), .C0(n934), .Y(
        block_next[35]) );
  OAI221X2 U1505 ( .A0(n701), .A1(n1070), .B0(n997), .B1(n702), .C0(n935), .Y(
        block_next[34]) );
  OAI221X2 U1506 ( .A0(n701), .A1(n1065), .B0(n999), .B1(n702), .C0(n936), .Y(
        block_next[33]) );
  OAI221X2 U1507 ( .A0(n701), .A1(n1060), .B0(n1001), .B1(n702), .C0(n937), 
        .Y(block_next[32]) );
  OAI221X2 U1508 ( .A0(n711), .A1(n939), .B0(n706), .B1(n1222), .C0(n938), .Y(
        block_next[31]) );
  OAI221X2 U1509 ( .A0(n711), .A1(n941), .B0(n706), .B1(n1214), .C0(n940), .Y(
        block_next[30]) );
  OAI221X2 U1510 ( .A0(n711), .A1(n943), .B0(n706), .B1(n1209), .C0(n942), .Y(
        block_next[29]) );
  OAI221X2 U1511 ( .A0(n711), .A1(n945), .B0(n706), .B1(n1204), .C0(n944), .Y(
        block_next[28]) );
  OAI221X2 U1512 ( .A0(n711), .A1(n947), .B0(n706), .B1(n1199), .C0(n946), .Y(
        block_next[27]) );
  OAI221X2 U1513 ( .A0(n711), .A1(n949), .B0(n706), .B1(n1194), .C0(n948), .Y(
        block_next[26]) );
  OAI221X2 U1514 ( .A0(n711), .A1(n951), .B0(n706), .B1(n1189), .C0(n950), .Y(
        block_next[25]) );
  OAI221X2 U1515 ( .A0(n710), .A1(n953), .B0(n706), .B1(n1184), .C0(n952), .Y(
        block_next[24]) );
  OAI221X2 U1516 ( .A0(n710), .A1(n955), .B0(n706), .B1(n1179), .C0(n954), .Y(
        block_next[23]) );
  OAI221X2 U1517 ( .A0(n710), .A1(n957), .B0(n706), .B1(n1174), .C0(n956), .Y(
        block_next[22]) );
  OAI221X2 U1518 ( .A0(n710), .A1(n963), .B0(n707), .B1(n1159), .C0(n962), .Y(
        block_next[19]) );
  OAI221X2 U1519 ( .A0(n710), .A1(n965), .B0(n707), .B1(n1154), .C0(n964), .Y(
        block_next[18]) );
  OAI221X2 U1520 ( .A0(n710), .A1(n967), .B0(n707), .B1(n1149), .C0(n966), .Y(
        block_next[17]) );
  OAI221X2 U1521 ( .A0(n710), .A1(n969), .B0(n707), .B1(n1144), .C0(n968), .Y(
        block_next[16]) );
  OAI221X2 U1522 ( .A0(n710), .A1(n971), .B0(n707), .B1(n1139), .C0(n970), .Y(
        block_next[15]) );
  OAI221X2 U1523 ( .A0(n710), .A1(n973), .B0(n707), .B1(n1134), .C0(n972), .Y(
        block_next[14]) );
  OAI221X2 U1524 ( .A0(n710), .A1(n975), .B0(n707), .B1(n1129), .C0(n974), .Y(
        block_next[13]) );
  OAI221X2 U1525 ( .A0(n709), .A1(n977), .B0(n707), .B1(n1124), .C0(n976), .Y(
        block_next[12]) );
  OAI221X2 U1526 ( .A0(n709), .A1(n979), .B0(n707), .B1(n1119), .C0(n978), .Y(
        block_next[11]) );
  OAI221X2 U1527 ( .A0(n709), .A1(n981), .B0(n707), .B1(n1114), .C0(n980), .Y(
        block_next[10]) );
  OAI221X2 U1528 ( .A0(n709), .A1(n987), .B0(n708), .B1(n1099), .C0(n986), .Y(
        block_next[7]) );
  OAI221X2 U1529 ( .A0(n709), .A1(n989), .B0(n708), .B1(n1094), .C0(n988), .Y(
        block_next[6]) );
  OAI221X2 U1530 ( .A0(n709), .A1(n991), .B0(n708), .B1(n1089), .C0(n990), .Y(
        block_next[5]) );
  OAI221X2 U1531 ( .A0(n709), .A1(n993), .B0(n708), .B1(n1084), .C0(n992), .Y(
        block_next[4]) );
  OAI221X2 U1532 ( .A0(n709), .A1(n995), .B0(n708), .B1(n1079), .C0(n994), .Y(
        block_next[3]) );
  OAI221X2 U1533 ( .A0(n709), .A1(n997), .B0(n708), .B1(n1074), .C0(n996), .Y(
        block_next[2]) );
  OAI221X2 U1534 ( .A0(n709), .A1(n999), .B0(n708), .B1(n1069), .C0(n998), .Y(
        block_next[1]) );
  OAI221X2 U1535 ( .A0(n710), .A1(n1001), .B0(n708), .B1(n1064), .C0(n1000), 
        .Y(block_next[0]) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, \blocktag[7][24] , \blocktag[7][23] , \blocktag[7][22] ,
         \blocktag[7][21] , \blocktag[7][20] , \blocktag[7][19] ,
         \blocktag[7][18] , \blocktag[7][17] , \blocktag[7][16] ,
         \blocktag[7][15] , \blocktag[7][14] , \blocktag[7][12] ,
         \blocktag[7][11] , \blocktag[7][10] , \blocktag[7][9] ,
         \blocktag[7][8] , \blocktag[7][7] , \blocktag[7][6] ,
         \blocktag[7][5] , \blocktag[7][4] , \blocktag[7][3] ,
         \blocktag[7][1] , \blocktag[6][24] , \blocktag[6][23] ,
         \blocktag[6][22] , \blocktag[6][21] , \blocktag[6][20] ,
         \blocktag[6][19] , \blocktag[6][18] , \blocktag[6][17] ,
         \blocktag[6][16] , \blocktag[6][15] , \blocktag[6][14] ,
         \blocktag[6][12] , \blocktag[6][11] , \blocktag[6][10] ,
         \blocktag[6][9] , \blocktag[6][8] , \blocktag[6][7] ,
         \blocktag[6][6] , \blocktag[6][5] , \blocktag[6][4] ,
         \blocktag[6][3] , \blocktag[6][1] , \blocktag[5][24] ,
         \blocktag[5][23] , \blocktag[5][22] , \blocktag[5][21] ,
         \blocktag[5][20] , \blocktag[5][19] , \blocktag[5][18] ,
         \blocktag[5][17] , \blocktag[5][16] , \blocktag[5][15] ,
         \blocktag[5][14] , \blocktag[5][12] , \blocktag[5][11] ,
         \blocktag[5][10] , \blocktag[5][9] , \blocktag[5][8] ,
         \blocktag[5][7] , \blocktag[5][6] , \blocktag[5][5] ,
         \blocktag[5][4] , \blocktag[5][3] , \blocktag[5][1] ,
         \blocktag[4][24] , \blocktag[4][23] , \blocktag[4][22] ,
         \blocktag[4][21] , \blocktag[4][20] , \blocktag[4][19] ,
         \blocktag[4][18] , \blocktag[4][17] , \blocktag[4][16] ,
         \blocktag[4][15] , \blocktag[4][14] , \blocktag[4][12] ,
         \blocktag[4][11] , \blocktag[4][10] , \blocktag[4][9] ,
         \blocktag[4][8] , \blocktag[4][7] , \blocktag[4][6] ,
         \blocktag[4][5] , \blocktag[4][4] , \blocktag[4][3] ,
         \blocktag[4][1] , \blocktag[3][24] , \blocktag[3][23] ,
         \blocktag[3][22] , \blocktag[3][21] , \blocktag[3][20] ,
         \blocktag[3][19] , \blocktag[3][18] , \blocktag[3][17] ,
         \blocktag[3][16] , \blocktag[3][15] , \blocktag[3][14] ,
         \blocktag[3][12] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][9] , \blocktag[3][8] , \blocktag[3][7] ,
         \blocktag[3][6] , \blocktag[3][5] , \blocktag[3][4] ,
         \blocktag[3][3] , \blocktag[3][2] , \blocktag[3][1] ,
         \blocktag[3][0] , \blocktag[2][24] , \blocktag[2][23] ,
         \blocktag[2][22] , \blocktag[2][21] , \blocktag[2][20] ,
         \blocktag[2][19] , \blocktag[2][18] , \blocktag[2][17] ,
         \blocktag[2][16] , \blocktag[2][15] , \blocktag[2][14] ,
         \blocktag[2][12] , \blocktag[2][11] , \blocktag[2][10] ,
         \blocktag[2][9] , \blocktag[2][8] , \blocktag[2][7] ,
         \blocktag[2][6] , \blocktag[2][5] , \blocktag[2][4] ,
         \blocktag[2][3] , \blocktag[2][2] , \blocktag[2][1] ,
         \blocktag[2][0] , \blocktag[1][24] , \blocktag[1][23] ,
         \blocktag[1][22] , \blocktag[1][21] , \blocktag[1][20] ,
         \blocktag[1][19] , \blocktag[1][18] , \blocktag[1][17] ,
         \blocktag[1][16] , \blocktag[1][15] , \blocktag[1][14] ,
         \blocktag[1][12] , \blocktag[1][11] , \blocktag[1][10] ,
         \blocktag[1][9] , \blocktag[1][8] , \blocktag[1][7] ,
         \blocktag[1][6] , \blocktag[1][5] , \blocktag[1][4] ,
         \blocktag[1][3] , \blocktag[1][2] , \blocktag[1][1] ,
         \blocktag[1][0] , \blocktag[0][24] , \blocktag[0][23] ,
         \blocktag[0][22] , \blocktag[0][21] , \blocktag[0][20] ,
         \blocktag[0][19] , \blocktag[0][18] , \blocktag[0][17] ,
         \blocktag[0][16] , \blocktag[0][15] , \blocktag[0][14] ,
         \blocktag[0][12] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][9] , \blocktag[0][8] , \blocktag[0][7] ,
         \blocktag[0][6] , \blocktag[0][5] , \blocktag[0][4] ,
         \blocktag[0][3] , \blocktag[0][2] , \blocktag[0][1] ,
         \blocktag[0][0] , valid, dirty, \block[7][127] , \block[7][126] ,
         \block[7][125] , \block[7][124] , \block[7][123] , \block[7][122] ,
         \block[7][121] , \block[7][120] , \block[7][119] , \block[7][118] ,
         \block[7][117] , \block[7][116] , \block[7][115] , \block[7][114] ,
         \block[7][113] , \block[7][112] , \block[7][110] , \block[7][109] ,
         \block[7][108] , \block[7][107] , \block[7][106] , \block[7][104] ,
         \block[7][103] , \block[7][102] , \block[7][101] , \block[7][100] ,
         \block[7][99] , \block[7][98] , \block[7][97] , \block[7][96] ,
         \block[7][92] , \block[7][91] , \block[7][90] , \block[7][89] ,
         \block[7][88] , \block[7][87] , \block[7][86] , \block[7][85] ,
         \block[7][84] , \block[7][83] , \block[7][82] , \block[7][81] ,
         \block[7][80] , \block[7][79] , \block[7][78] , \block[7][77] ,
         \block[7][76] , \block[7][75] , \block[7][74] , \block[7][72] ,
         \block[7][71] , \block[7][70] , \block[7][69] , \block[7][68] ,
         \block[7][67] , \block[7][66] , \block[7][65] , \block[7][64] ,
         \block[7][62] , \block[7][61] , \block[7][60] , \block[7][59] ,
         \block[7][58] , \block[7][57] , \block[7][56] , \block[7][55] ,
         \block[7][54] , \block[7][53] , \block[7][52] , \block[7][51] ,
         \block[7][50] , \block[7][49] , \block[7][48] , \block[7][46] ,
         \block[7][45] , \block[7][44] , \block[7][43] , \block[7][42] ,
         \block[7][40] , \block[7][39] , \block[7][38] , \block[7][37] ,
         \block[7][36] , \block[7][35] , \block[7][34] , \block[7][33] ,
         \block[7][32] , \block[7][31] , \block[7][30] , \block[7][29] ,
         \block[7][28] , \block[7][27] , \block[7][26] , \block[7][25] ,
         \block[7][24] , \block[7][23] , \block[7][22] , \block[7][21] ,
         \block[7][20] , \block[7][19] , \block[7][18] , \block[7][17] ,
         \block[7][16] , \block[7][15] , \block[7][14] , \block[7][13] ,
         \block[7][11] , \block[7][10] , \block[7][9] , \block[7][8] ,
         \block[7][7] , \block[7][6] , \block[7][5] , \block[7][4] ,
         \block[7][3] , \block[7][2] , \block[7][1] , \block[7][0] ,
         \block[6][127] , \block[6][126] , \block[6][125] , \block[6][124] ,
         \block[6][123] , \block[6][122] , \block[6][121] , \block[6][120] ,
         \block[6][119] , \block[6][118] , \block[6][117] , \block[6][116] ,
         \block[6][115] , \block[6][114] , \block[6][113] , \block[6][112] ,
         \block[6][110] , \block[6][109] , \block[6][108] , \block[6][107] ,
         \block[6][106] , \block[6][104] , \block[6][103] , \block[6][102] ,
         \block[6][101] , \block[6][100] , \block[6][99] , \block[6][98] ,
         \block[6][97] , \block[6][96] , \block[6][92] , \block[6][91] ,
         \block[6][90] , \block[6][89] , \block[6][88] , \block[6][87] ,
         \block[6][86] , \block[6][85] , \block[6][84] , \block[6][83] ,
         \block[6][82] , \block[6][81] , \block[6][80] , \block[6][79] ,
         \block[6][78] , \block[6][77] , \block[6][76] , \block[6][75] ,
         \block[6][74] , \block[6][72] , \block[6][71] , \block[6][70] ,
         \block[6][69] , \block[6][68] , \block[6][67] , \block[6][66] ,
         \block[6][65] , \block[6][64] , \block[6][62] , \block[6][61] ,
         \block[6][60] , \block[6][59] , \block[6][58] , \block[6][57] ,
         \block[6][56] , \block[6][55] , \block[6][54] , \block[6][53] ,
         \block[6][52] , \block[6][51] , \block[6][50] , \block[6][49] ,
         \block[6][48] , \block[6][46] , \block[6][45] , \block[6][44] ,
         \block[6][43] , \block[6][42] , \block[6][40] , \block[6][39] ,
         \block[6][38] , \block[6][37] , \block[6][36] , \block[6][35] ,
         \block[6][34] , \block[6][33] , \block[6][32] , \block[6][31] ,
         \block[6][30] , \block[6][29] , \block[6][28] , \block[6][27] ,
         \block[6][26] , \block[6][25] , \block[6][24] , \block[6][23] ,
         \block[6][22] , \block[6][21] , \block[6][20] , \block[6][19] ,
         \block[6][18] , \block[6][17] , \block[6][16] , \block[6][15] ,
         \block[6][14] , \block[6][13] , \block[6][11] , \block[6][10] ,
         \block[6][9] , \block[6][8] , \block[6][7] , \block[6][6] ,
         \block[6][5] , \block[6][4] , \block[6][3] , \block[6][2] ,
         \block[6][1] , \block[6][0] , \block[5][127] , \block[5][126] ,
         \block[5][125] , \block[5][124] , \block[5][123] , \block[5][122] ,
         \block[5][121] , \block[5][120] , \block[5][119] , \block[5][118] ,
         \block[5][117] , \block[5][116] , \block[5][115] , \block[5][114] ,
         \block[5][113] , \block[5][112] , \block[5][110] , \block[5][109] ,
         \block[5][108] , \block[5][107] , \block[5][106] , \block[5][104] ,
         \block[5][103] , \block[5][102] , \block[5][101] , \block[5][100] ,
         \block[5][99] , \block[5][98] , \block[5][97] , \block[5][96] ,
         \block[5][92] , \block[5][91] , \block[5][90] , \block[5][89] ,
         \block[5][88] , \block[5][87] , \block[5][86] , \block[5][85] ,
         \block[5][84] , \block[5][83] , \block[5][82] , \block[5][81] ,
         \block[5][80] , \block[5][79] , \block[5][78] , \block[5][77] ,
         \block[5][76] , \block[5][75] , \block[5][74] , \block[5][72] ,
         \block[5][71] , \block[5][70] , \block[5][69] , \block[5][68] ,
         \block[5][67] , \block[5][66] , \block[5][65] , \block[5][64] ,
         \block[5][62] , \block[5][61] , \block[5][60] , \block[5][59] ,
         \block[5][58] , \block[5][57] , \block[5][56] , \block[5][55] ,
         \block[5][54] , \block[5][53] , \block[5][52] , \block[5][51] ,
         \block[5][50] , \block[5][49] , \block[5][48] , \block[5][46] ,
         \block[5][45] , \block[5][44] , \block[5][43] , \block[5][42] ,
         \block[5][40] , \block[5][39] , \block[5][38] , \block[5][37] ,
         \block[5][36] , \block[5][35] , \block[5][34] , \block[5][33] ,
         \block[5][32] , \block[5][31] , \block[5][30] , \block[5][29] ,
         \block[5][28] , \block[5][27] , \block[5][26] , \block[5][25] ,
         \block[5][24] , \block[5][23] , \block[5][22] , \block[5][21] ,
         \block[5][20] , \block[5][19] , \block[5][18] , \block[5][17] ,
         \block[5][16] , \block[5][15] , \block[5][14] , \block[5][13] ,
         \block[5][11] , \block[5][10] , \block[5][9] , \block[5][8] ,
         \block[5][7] , \block[5][6] , \block[5][5] , \block[5][4] ,
         \block[5][3] , \block[5][2] , \block[5][1] , \block[5][0] ,
         \block[4][127] , \block[4][126] , \block[4][125] , \block[4][124] ,
         \block[4][123] , \block[4][122] , \block[4][121] , \block[4][120] ,
         \block[4][119] , \block[4][118] , \block[4][117] , \block[4][116] ,
         \block[4][115] , \block[4][114] , \block[4][113] , \block[4][112] ,
         \block[4][110] , \block[4][109] , \block[4][108] , \block[4][107] ,
         \block[4][106] , \block[4][104] , \block[4][103] , \block[4][102] ,
         \block[4][101] , \block[4][100] , \block[4][99] , \block[4][98] ,
         \block[4][97] , \block[4][96] , \block[4][92] , \block[4][91] ,
         \block[4][90] , \block[4][89] , \block[4][88] , \block[4][87] ,
         \block[4][86] , \block[4][85] , \block[4][84] , \block[4][83] ,
         \block[4][82] , \block[4][81] , \block[4][80] , \block[4][79] ,
         \block[4][78] , \block[4][77] , \block[4][76] , \block[4][75] ,
         \block[4][74] , \block[4][72] , \block[4][71] , \block[4][70] ,
         \block[4][69] , \block[4][68] , \block[4][67] , \block[4][66] ,
         \block[4][65] , \block[4][64] , \block[4][62] , \block[4][61] ,
         \block[4][60] , \block[4][59] , \block[4][58] , \block[4][57] ,
         \block[4][56] , \block[4][55] , \block[4][54] , \block[4][53] ,
         \block[4][52] , \block[4][51] , \block[4][50] , \block[4][49] ,
         \block[4][48] , \block[4][46] , \block[4][45] , \block[4][44] ,
         \block[4][43] , \block[4][42] , \block[4][40] , \block[4][39] ,
         \block[4][38] , \block[4][37] , \block[4][36] , \block[4][35] ,
         \block[4][34] , \block[4][33] , \block[4][32] , \block[4][31] ,
         \block[4][30] , \block[4][29] , \block[4][28] , \block[4][27] ,
         \block[4][26] , \block[4][25] , \block[4][24] , \block[4][23] ,
         \block[4][22] , \block[4][21] , \block[4][20] , \block[4][19] ,
         \block[4][18] , \block[4][17] , \block[4][16] , \block[4][15] ,
         \block[4][14] , \block[4][13] , \block[4][11] , \block[4][10] ,
         \block[4][9] , \block[4][8] , \block[4][7] , \block[4][6] ,
         \block[4][5] , \block[4][4] , \block[4][3] , \block[4][2] ,
         \block[4][1] , \block[4][0] , \block[3][127] , \block[3][126] ,
         \block[3][125] , \block[3][124] , \block[3][123] , \block[3][122] ,
         \block[3][121] , \block[3][120] , \block[3][119] , \block[3][118] ,
         \block[3][117] , \block[3][116] , \block[3][115] , \block[3][114] ,
         \block[3][113] , \block[3][112] , \block[3][111] , \block[3][110] ,
         \block[3][109] , \block[3][108] , \block[3][107] , \block[3][106] ,
         \block[3][105] , \block[3][104] , \block[3][103] , \block[3][102] ,
         \block[3][101] , \block[3][100] , \block[3][99] , \block[3][98] ,
         \block[3][97] , \block[3][96] , \block[3][92] , \block[3][91] ,
         \block[3][90] , \block[3][89] , \block[3][88] , \block[3][87] ,
         \block[3][86] , \block[3][85] , \block[3][84] , \block[3][83] ,
         \block[3][82] , \block[3][81] , \block[3][80] , \block[3][79] ,
         \block[3][78] , \block[3][77] , \block[3][76] , \block[3][75] ,
         \block[3][74] , \block[3][73] , \block[3][72] , \block[3][71] ,
         \block[3][70] , \block[3][69] , \block[3][68] , \block[3][67] ,
         \block[3][66] , \block[3][65] , \block[3][64] , \block[3][62] ,
         \block[3][61] , \block[3][60] , \block[3][59] , \block[3][58] ,
         \block[3][57] , \block[3][56] , \block[3][55] , \block[3][54] ,
         \block[3][53] , \block[3][52] , \block[3][51] , \block[3][50] ,
         \block[3][49] , \block[3][48] , \block[3][47] , \block[3][46] ,
         \block[3][45] , \block[3][44] , \block[3][43] , \block[3][42] ,
         \block[3][41] , \block[3][40] , \block[3][39] , \block[3][38] ,
         \block[3][37] , \block[3][36] , \block[3][35] , \block[3][34] ,
         \block[3][33] , \block[3][32] , \block[3][31] , \block[3][30] ,
         \block[3][29] , \block[3][28] , \block[3][27] , \block[3][26] ,
         \block[3][25] , \block[3][24] , \block[3][23] , \block[3][22] ,
         \block[3][21] , \block[3][20] , \block[3][19] , \block[3][18] ,
         \block[3][17] , \block[3][16] , \block[3][15] , \block[3][14] ,
         \block[3][13] , \block[3][11] , \block[3][10] , \block[3][9] ,
         \block[3][8] , \block[3][7] , \block[3][6] , \block[3][5] ,
         \block[3][4] , \block[3][3] , \block[3][2] , \block[3][1] ,
         \block[3][0] , \block[2][127] , \block[2][126] , \block[2][125] ,
         \block[2][124] , \block[2][123] , \block[2][122] , \block[2][121] ,
         \block[2][120] , \block[2][119] , \block[2][118] , \block[2][117] ,
         \block[2][116] , \block[2][115] , \block[2][114] , \block[2][113] ,
         \block[2][112] , \block[2][111] , \block[2][110] , \block[2][109] ,
         \block[2][108] , \block[2][107] , \block[2][106] , \block[2][105] ,
         \block[2][104] , \block[2][103] , \block[2][102] , \block[2][101] ,
         \block[2][100] , \block[2][99] , \block[2][98] , \block[2][97] ,
         \block[2][96] , \block[2][92] , \block[2][91] , \block[2][90] ,
         \block[2][89] , \block[2][88] , \block[2][87] , \block[2][86] ,
         \block[2][85] , \block[2][84] , \block[2][83] , \block[2][82] ,
         \block[2][81] , \block[2][80] , \block[2][79] , \block[2][78] ,
         \block[2][77] , \block[2][76] , \block[2][75] , \block[2][74] ,
         \block[2][73] , \block[2][72] , \block[2][71] , \block[2][70] ,
         \block[2][69] , \block[2][68] , \block[2][67] , \block[2][66] ,
         \block[2][65] , \block[2][64] , \block[2][62] , \block[2][61] ,
         \block[2][60] , \block[2][59] , \block[2][58] , \block[2][57] ,
         \block[2][56] , \block[2][55] , \block[2][54] , \block[2][53] ,
         \block[2][52] , \block[2][51] , \block[2][50] , \block[2][49] ,
         \block[2][48] , \block[2][47] , \block[2][46] , \block[2][45] ,
         \block[2][44] , \block[2][43] , \block[2][42] , \block[2][41] ,
         \block[2][40] , \block[2][39] , \block[2][38] , \block[2][37] ,
         \block[2][36] , \block[2][35] , \block[2][34] , \block[2][33] ,
         \block[2][32] , \block[2][31] , \block[2][30] , \block[2][29] ,
         \block[2][28] , \block[2][27] , \block[2][26] , \block[2][25] ,
         \block[2][24] , \block[2][23] , \block[2][22] , \block[2][21] ,
         \block[2][20] , \block[2][19] , \block[2][18] , \block[2][17] ,
         \block[2][16] , \block[2][15] , \block[2][14] , \block[2][13] ,
         \block[2][11] , \block[2][10] , \block[2][9] , \block[2][8] ,
         \block[2][7] , \block[2][6] , \block[2][5] , \block[2][4] ,
         \block[2][3] , \block[2][2] , \block[2][1] , \block[2][0] ,
         \block[1][127] , \block[1][126] , \block[1][125] , \block[1][124] ,
         \block[1][123] , \block[1][122] , \block[1][121] , \block[1][120] ,
         \block[1][119] , \block[1][118] , \block[1][117] , \block[1][116] ,
         \block[1][115] , \block[1][114] , \block[1][113] , \block[1][112] ,
         \block[1][111] , \block[1][110] , \block[1][109] , \block[1][108] ,
         \block[1][107] , \block[1][106] , \block[1][105] , \block[1][104] ,
         \block[1][103] , \block[1][102] , \block[1][101] , \block[1][100] ,
         \block[1][99] , \block[1][98] , \block[1][97] , \block[1][96] ,
         \block[1][92] , \block[1][91] , \block[1][90] , \block[1][89] ,
         \block[1][88] , \block[1][87] , \block[1][86] , \block[1][85] ,
         \block[1][84] , \block[1][83] , \block[1][82] , \block[1][81] ,
         \block[1][80] , \block[1][79] , \block[1][78] , \block[1][77] ,
         \block[1][76] , \block[1][75] , \block[1][74] , \block[1][73] ,
         \block[1][72] , \block[1][71] , \block[1][70] , \block[1][69] ,
         \block[1][68] , \block[1][67] , \block[1][66] , \block[1][65] ,
         \block[1][64] , \block[1][62] , \block[1][61] , \block[1][60] ,
         \block[1][59] , \block[1][58] , \block[1][57] , \block[1][56] ,
         \block[1][55] , \block[1][54] , \block[1][53] , \block[1][52] ,
         \block[1][51] , \block[1][50] , \block[1][49] , \block[1][48] ,
         \block[1][47] , \block[1][46] , \block[1][45] , \block[1][44] ,
         \block[1][43] , \block[1][42] , \block[1][41] , \block[1][40] ,
         \block[1][39] , \block[1][38] , \block[1][37] , \block[1][36] ,
         \block[1][35] , \block[1][34] , \block[1][33] , \block[1][32] ,
         \block[1][31] , \block[1][30] , \block[1][29] , \block[1][28] ,
         \block[1][27] , \block[1][26] , \block[1][25] , \block[1][24] ,
         \block[1][23] , \block[1][22] , \block[1][21] , \block[1][20] ,
         \block[1][19] , \block[1][18] , \block[1][17] , \block[1][16] ,
         \block[1][15] , \block[1][14] , \block[1][13] , \block[1][11] ,
         \block[1][10] , \block[1][9] , \block[1][8] , \block[1][7] ,
         \block[1][6] , \block[1][5] , \block[1][4] , \block[1][3] ,
         \block[1][2] , \block[1][1] , \block[1][0] , \block[0][127] ,
         \block[0][126] , \block[0][125] , \block[0][124] , \block[0][123] ,
         \block[0][122] , \block[0][121] , \block[0][120] , \block[0][119] ,
         \block[0][118] , \block[0][117] , \block[0][116] , \block[0][115] ,
         \block[0][114] , \block[0][113] , \block[0][112] , \block[0][111] ,
         \block[0][110] , \block[0][109] , \block[0][108] , \block[0][107] ,
         \block[0][106] , \block[0][105] , \block[0][104] , \block[0][103] ,
         \block[0][102] , \block[0][101] , \block[0][100] , \block[0][99] ,
         \block[0][98] , \block[0][97] , \block[0][96] , \block[0][92] ,
         \block[0][91] , \block[0][90] , \block[0][89] , \block[0][88] ,
         \block[0][87] , \block[0][86] , \block[0][85] , \block[0][84] ,
         \block[0][83] , \block[0][82] , \block[0][81] , \block[0][80] ,
         \block[0][79] , \block[0][78] , \block[0][77] , \block[0][76] ,
         \block[0][75] , \block[0][74] , \block[0][73] , \block[0][72] ,
         \block[0][71] , \block[0][70] , \block[0][69] , \block[0][68] ,
         \block[0][67] , \block[0][66] , \block[0][65] , \block[0][64] ,
         \block[0][62] , \block[0][61] , \block[0][60] , \block[0][59] ,
         \block[0][58] , \block[0][57] , \block[0][56] , \block[0][55] ,
         \block[0][54] , \block[0][53] , \block[0][52] , \block[0][51] ,
         \block[0][50] , \block[0][49] , \block[0][48] , \block[0][47] ,
         \block[0][46] , \block[0][45] , \block[0][44] , \block[0][43] ,
         \block[0][42] , \block[0][41] , \block[0][40] , \block[0][39] ,
         \block[0][38] , \block[0][37] , \block[0][36] , \block[0][35] ,
         \block[0][34] , \block[0][33] , \block[0][32] , \block[0][31] ,
         \block[0][30] , \block[0][29] , \block[0][28] , \block[0][27] ,
         \block[0][26] , \block[0][25] , \block[0][24] , \block[0][23] ,
         \block[0][22] , \block[0][21] , \block[0][20] , \block[0][19] ,
         \block[0][18] , \block[0][17] , \block[0][16] , \block[0][15] ,
         \block[0][14] , \block[0][13] , \block[0][11] , \block[0][10] ,
         \block[0][9] , \block[0][8] , \block[0][7] , \block[0][6] ,
         \block[0][5] , \block[0][4] , \block[0][3] , \block[0][2] ,
         \block[0][1] , \block[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n111, n113, n117, n120, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n502, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n859, n860, n861,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  EDFFX1 \block_reg[7][121]  ( .D(block_next[121]), .E(n791), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFX1 \block_reg[7][120]  ( .D(block_next[120]), .E(n792), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFX1 \block_reg[7][119]  ( .D(block_next[119]), .E(n791), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFX1 \block_reg[7][118]  ( .D(block_next[118]), .E(n798), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFX1 \block_reg[7][117]  ( .D(block_next[117]), .E(n794), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFX1 \block_reg[7][116]  ( .D(block_next[116]), .E(n795), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFX1 \block_reg[7][115]  ( .D(block_next[115]), .E(n797), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFX1 \block_reg[7][114]  ( .D(block_next[114]), .E(n798), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFX1 \block_reg[7][113]  ( .D(block_next[113]), .E(n798), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFX1 \block_reg[7][112]  ( .D(block_next[112]), .E(n792), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFX1 \block_reg[7][111]  ( .D(block_next[111]), .E(n795), .CK(clk), .QN(
        n292) );
  EDFFX1 \block_reg[7][110]  ( .D(block_next[110]), .E(n791), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFX1 \block_reg[7][109]  ( .D(block_next[109]), .E(n307), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFX1 \block_reg[7][108]  ( .D(block_next[108]), .E(n793), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFX1 \block_reg[7][107]  ( .D(block_next[107]), .E(n796), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFX1 \block_reg[7][106]  ( .D(block_next[106]), .E(n794), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFX1 \block_reg[7][105]  ( .D(block_next[105]), .E(n797), .CK(clk), .QN(
        n284) );
  EDFFX1 \block_reg[7][104]  ( .D(block_next[104]), .E(n795), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFX1 \block_reg[7][103]  ( .D(block_next[103]), .E(n794), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFX1 \block_reg[7][102]  ( .D(block_next[102]), .E(n796), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFX1 \block_reg[7][101]  ( .D(block_next[101]), .E(n793), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFX1 \block_reg[7][100]  ( .D(block_next[100]), .E(n307), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFX1 \block_reg[7][99]  ( .D(block_next[99]), .E(n791), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFX1 \block_reg[7][98]  ( .D(block_next[98]), .E(n792), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFX1 \block_reg[7][97]  ( .D(block_next[97]), .E(n798), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFX1 \block_reg[7][96]  ( .D(block_next[96]), .E(n797), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFX1 \block_reg[7][89]  ( .D(block_next[89]), .E(n798), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFX1 \block_reg[7][88]  ( .D(block_next[88]), .E(n798), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFX1 \block_reg[7][87]  ( .D(block_next[87]), .E(n798), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFX1 \block_reg[7][86]  ( .D(block_next[86]), .E(n798), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFX1 \block_reg[7][85]  ( .D(block_next[85]), .E(n798), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFX1 \block_reg[7][84]  ( .D(block_next[84]), .E(n798), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFX1 \block_reg[7][83]  ( .D(block_next[83]), .E(n798), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFX1 \block_reg[7][82]  ( .D(block_next[82]), .E(n798), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFX1 \block_reg[7][81]  ( .D(block_next[81]), .E(n798), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFX1 \block_reg[7][80]  ( .D(block_next[80]), .E(n798), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFX1 \block_reg[7][79]  ( .D(block_next[79]), .E(n798), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFX1 \block_reg[7][78]  ( .D(block_next[78]), .E(n797), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFX1 \block_reg[7][77]  ( .D(block_next[77]), .E(n797), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFX1 \block_reg[7][76]  ( .D(block_next[76]), .E(n797), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFX1 \block_reg[7][75]  ( .D(block_next[75]), .E(n797), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFX1 \block_reg[7][74]  ( .D(block_next[74]), .E(n797), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFX1 \block_reg[7][73]  ( .D(block_next[73]), .E(n797), .CK(clk), .QN(n280) );
  EDFFX1 \block_reg[7][72]  ( .D(block_next[72]), .E(n797), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFX1 \block_reg[7][71]  ( .D(block_next[71]), .E(n797), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFX1 \block_reg[7][70]  ( .D(block_next[70]), .E(n797), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFX1 \block_reg[7][69]  ( .D(block_next[69]), .E(n797), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFX1 \block_reg[7][68]  ( .D(block_next[68]), .E(n797), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFX1 \block_reg[7][67]  ( .D(block_next[67]), .E(n797), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFX1 \block_reg[7][66]  ( .D(block_next[66]), .E(n797), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFX1 \block_reg[7][65]  ( .D(block_next[65]), .E(n796), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFX1 \block_reg[7][64]  ( .D(block_next[64]), .E(n796), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFX1 \block_reg[7][57]  ( .D(block_next[57]), .E(n796), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFX1 \block_reg[7][56]  ( .D(block_next[56]), .E(n796), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFX1 \block_reg[7][55]  ( .D(block_next[55]), .E(n796), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFX1 \block_reg[7][54]  ( .D(block_next[54]), .E(n796), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n796), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n795), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[7][51]  ( .D(block_next[51]), .E(n795), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFX1 \block_reg[7][50]  ( .D(block_next[50]), .E(n795), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n795), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[7][48]  ( .D(block_next[48]), .E(n795), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFX1 \block_reg[7][47]  ( .D(block_next[47]), .E(n795), .CK(clk), .QN(n288) );
  EDFFX1 \block_reg[7][46]  ( .D(block_next[46]), .E(n795), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFX1 \block_reg[7][45]  ( .D(block_next[45]), .E(n795), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFX1 \block_reg[7][44]  ( .D(block_next[44]), .E(n795), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFX1 \block_reg[7][43]  ( .D(block_next[43]), .E(n795), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFX1 \block_reg[7][42]  ( .D(block_next[42]), .E(n795), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n795), .CK(clk), .QN(n276) );
  EDFFX1 \block_reg[7][40]  ( .D(block_next[40]), .E(n795), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFX1 \block_reg[7][39]  ( .D(block_next[39]), .E(n794), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n794), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n794), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n794), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n794), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n794), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFX1 \block_reg[7][33]  ( .D(block_next[33]), .E(n794), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n794), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[7][25]  ( .D(block_next[25]), .E(n793), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFX1 \block_reg[7][24]  ( .D(block_next[24]), .E(n793), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFX1 \block_reg[7][23]  ( .D(block_next[23]), .E(n793), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFX1 \block_reg[7][22]  ( .D(block_next[22]), .E(n793), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFX1 \block_reg[7][21]  ( .D(block_next[21]), .E(n793), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFX1 \block_reg[7][20]  ( .D(block_next[20]), .E(n793), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFX1 \block_reg[7][19]  ( .D(block_next[19]), .E(n793), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFX1 \block_reg[7][18]  ( .D(block_next[18]), .E(n793), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFX1 \block_reg[7][17]  ( .D(block_next[17]), .E(n793), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFX1 \block_reg[7][16]  ( .D(block_next[16]), .E(n793), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFX1 \block_reg[7][15]  ( .D(block_next[15]), .E(n793), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFX1 \block_reg[7][14]  ( .D(block_next[14]), .E(n793), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFX1 \block_reg[7][13]  ( .D(block_next[13]), .E(n792), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFX1 \block_reg[7][12]  ( .D(block_next[12]), .E(n792), .CK(clk), .QN(n300) );
  EDFFX1 \block_reg[7][11]  ( .D(block_next[11]), .E(n792), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFX1 \block_reg[7][10]  ( .D(block_next[10]), .E(n792), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFX1 \block_reg[7][9]  ( .D(block_next[9]), .E(n792), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFX1 \block_reg[7][8]  ( .D(block_next[8]), .E(n792), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFX1 \block_reg[7][7]  ( .D(block_next[7]), .E(n792), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFX1 \block_reg[7][6]  ( .D(block_next[6]), .E(n792), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFX1 \block_reg[7][5]  ( .D(block_next[5]), .E(n792), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFX1 \block_reg[7][4]  ( .D(block_next[4]), .E(n792), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFX1 \block_reg[7][3]  ( .D(block_next[3]), .E(n792), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFX1 \block_reg[7][2]  ( .D(block_next[2]), .E(n792), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFX1 \block_reg[7][1]  ( .D(block_next[1]), .E(n792), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFX1 \block_reg[7][0]  ( .D(block_next[0]), .E(n307), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFX1 \block_reg[3][121]  ( .D(block_next[121]), .E(n824), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFX1 \block_reg[3][120]  ( .D(block_next[120]), .E(n830), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFX1 \block_reg[3][119]  ( .D(block_next[119]), .E(n825), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFX1 \block_reg[3][118]  ( .D(block_next[118]), .E(n829), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFX1 \block_reg[3][117]  ( .D(block_next[117]), .E(n828), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFX1 \block_reg[3][116]  ( .D(block_next[116]), .E(n826), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFX1 \block_reg[3][115]  ( .D(block_next[115]), .E(n827), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFX1 \block_reg[3][114]  ( .D(block_next[114]), .E(n829), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFX1 \block_reg[3][113]  ( .D(block_next[113]), .E(n830), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFX1 \block_reg[3][112]  ( .D(block_next[112]), .E(n830), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFX1 \block_reg[3][111]  ( .D(block_next[111]), .E(n823), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFX1 \block_reg[3][110]  ( .D(block_next[110]), .E(n824), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFX1 \block_reg[3][109]  ( .D(block_next[109]), .E(n825), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFX1 \block_reg[3][108]  ( .D(block_next[108]), .E(n828), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFX1 \block_reg[3][107]  ( .D(block_next[107]), .E(n826), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFX1 \block_reg[3][106]  ( .D(block_next[106]), .E(n827), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFX1 \block_reg[3][105]  ( .D(block_next[105]), .E(n829), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFX1 \block_reg[3][104]  ( .D(block_next[104]), .E(n825), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFX1 \block_reg[3][103]  ( .D(block_next[103]), .E(n824), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFX1 \block_reg[3][102]  ( .D(block_next[102]), .E(n823), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFX1 \block_reg[3][101]  ( .D(block_next[101]), .E(n830), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFX1 \block_reg[3][100]  ( .D(block_next[100]), .E(n829), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFX1 \block_reg[3][99]  ( .D(block_next[99]), .E(n827), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFX1 \block_reg[3][98]  ( .D(block_next[98]), .E(n826), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFX1 \block_reg[3][97]  ( .D(block_next[97]), .E(n828), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFX1 \block_reg[3][96]  ( .D(block_next[96]), .E(n825), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFX1 \block_reg[3][89]  ( .D(block_next[89]), .E(n830), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFX1 \block_reg[3][88]  ( .D(block_next[88]), .E(n830), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFX1 \block_reg[3][87]  ( .D(block_next[87]), .E(n830), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFX1 \block_reg[3][86]  ( .D(block_next[86]), .E(n830), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFX1 \block_reg[3][85]  ( .D(block_next[85]), .E(n830), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFX1 \block_reg[3][84]  ( .D(block_next[84]), .E(n830), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFX1 \block_reg[3][83]  ( .D(block_next[83]), .E(n830), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFX1 \block_reg[3][82]  ( .D(block_next[82]), .E(n830), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFX1 \block_reg[3][81]  ( .D(block_next[81]), .E(n830), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFX1 \block_reg[3][80]  ( .D(block_next[80]), .E(n830), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFX1 \block_reg[3][79]  ( .D(block_next[79]), .E(n830), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFX1 \block_reg[3][78]  ( .D(block_next[78]), .E(n829), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFX1 \block_reg[3][77]  ( .D(block_next[77]), .E(n829), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFX1 \block_reg[3][76]  ( .D(block_next[76]), .E(n829), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFX1 \block_reg[3][75]  ( .D(block_next[75]), .E(n829), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFX1 \block_reg[3][74]  ( .D(block_next[74]), .E(n829), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFX1 \block_reg[3][73]  ( .D(block_next[73]), .E(n829), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFX1 \block_reg[3][72]  ( .D(block_next[72]), .E(n829), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFX1 \block_reg[3][71]  ( .D(block_next[71]), .E(n829), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFX1 \block_reg[3][70]  ( .D(block_next[70]), .E(n829), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFX1 \block_reg[3][69]  ( .D(block_next[69]), .E(n829), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFX1 \block_reg[3][68]  ( .D(block_next[68]), .E(n829), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFX1 \block_reg[3][67]  ( .D(block_next[67]), .E(n829), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFX1 \block_reg[3][66]  ( .D(block_next[66]), .E(n829), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFX1 \block_reg[3][65]  ( .D(block_next[65]), .E(n828), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFX1 \block_reg[3][64]  ( .D(block_next[64]), .E(n828), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[3][57]  ( .D(block_next[57]), .E(n828), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFX1 \block_reg[3][56]  ( .D(block_next[56]), .E(n828), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFX1 \block_reg[3][55]  ( .D(block_next[55]), .E(n828), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFX1 \block_reg[3][54]  ( .D(block_next[54]), .E(n828), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n828), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n827), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[3][51]  ( .D(block_next[51]), .E(n827), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFX1 \block_reg[3][50]  ( .D(block_next[50]), .E(n827), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n827), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[3][48]  ( .D(block_next[48]), .E(n827), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFX1 \block_reg[3][47]  ( .D(block_next[47]), .E(n827), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFX1 \block_reg[3][46]  ( .D(block_next[46]), .E(n827), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFX1 \block_reg[3][45]  ( .D(block_next[45]), .E(n827), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFX1 \block_reg[3][44]  ( .D(block_next[44]), .E(n827), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFX1 \block_reg[3][43]  ( .D(block_next[43]), .E(n827), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFX1 \block_reg[3][42]  ( .D(block_next[42]), .E(n827), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n827), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[3][40]  ( .D(block_next[40]), .E(n827), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFX1 \block_reg[3][39]  ( .D(block_next[39]), .E(n826), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n826), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n826), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n826), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n826), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n826), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[3][33]  ( .D(block_next[33]), .E(n826), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n826), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[3][25]  ( .D(block_next[25]), .E(n825), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFX1 \block_reg[3][24]  ( .D(block_next[24]), .E(n825), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFX1 \block_reg[3][23]  ( .D(block_next[23]), .E(n825), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFX1 \block_reg[3][22]  ( .D(block_next[22]), .E(n825), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFX1 \block_reg[3][21]  ( .D(block_next[21]), .E(n825), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n825), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFX1 \block_reg[3][19]  ( .D(block_next[19]), .E(n825), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFX1 \block_reg[3][18]  ( .D(block_next[18]), .E(n825), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFX1 \block_reg[3][17]  ( .D(block_next[17]), .E(n825), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFX1 \block_reg[3][16]  ( .D(block_next[16]), .E(n825), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFX1 \block_reg[3][15]  ( .D(block_next[15]), .E(n825), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFX1 \block_reg[3][14]  ( .D(block_next[14]), .E(n825), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFX1 \block_reg[3][13]  ( .D(block_next[13]), .E(n823), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFX1 \block_reg[3][12]  ( .D(block_next[12]), .E(n830), .CK(clk), .QN(n296) );
  EDFFX1 \block_reg[3][11]  ( .D(block_next[11]), .E(n306), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFX1 \block_reg[3][10]  ( .D(block_next[10]), .E(n829), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFX1 \block_reg[3][9]  ( .D(block_next[9]), .E(n827), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFX1 \block_reg[3][8]  ( .D(block_next[8]), .E(n826), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFX1 \block_reg[3][7]  ( .D(block_next[7]), .E(n828), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFX1 \block_reg[3][6]  ( .D(block_next[6]), .E(n825), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFX1 \block_reg[3][5]  ( .D(block_next[5]), .E(n306), .CK(clk), .Q(
        \block[3][5] ) );
  EDFFX1 \block_reg[3][4]  ( .D(block_next[4]), .E(n824), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFX1 \block_reg[3][3]  ( .D(block_next[3]), .E(n823), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFX1 \block_reg[3][2]  ( .D(block_next[2]), .E(n824), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFX1 \block_reg[3][1]  ( .D(block_next[1]), .E(n823), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFX1 \block_reg[3][0]  ( .D(block_next[0]), .E(n824), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFX1 \block_reg[5][121]  ( .D(block_next[121]), .E(n807), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFX1 \block_reg[5][120]  ( .D(block_next[120]), .E(n808), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFX1 \block_reg[5][119]  ( .D(block_next[119]), .E(n807), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFX1 \block_reg[5][118]  ( .D(block_next[118]), .E(n814), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFX1 \block_reg[5][117]  ( .D(block_next[117]), .E(n810), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFX1 \block_reg[5][116]  ( .D(block_next[116]), .E(n811), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFX1 \block_reg[5][115]  ( .D(block_next[115]), .E(n813), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFX1 \block_reg[5][114]  ( .D(block_next[114]), .E(n814), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFX1 \block_reg[5][113]  ( .D(block_next[113]), .E(n814), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFX1 \block_reg[5][112]  ( .D(block_next[112]), .E(n808), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFX1 \block_reg[5][111]  ( .D(block_next[111]), .E(n811), .CK(clk), .QN(
        n290) );
  EDFFX1 \block_reg[5][110]  ( .D(block_next[110]), .E(n807), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFX1 \block_reg[5][109]  ( .D(block_next[109]), .E(n305), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFX1 \block_reg[5][108]  ( .D(block_next[108]), .E(n809), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFX1 \block_reg[5][107]  ( .D(block_next[107]), .E(n812), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFX1 \block_reg[5][106]  ( .D(block_next[106]), .E(n810), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFX1 \block_reg[5][105]  ( .D(block_next[105]), .E(n813), .CK(clk), .QN(
        n282) );
  EDFFX1 \block_reg[5][104]  ( .D(block_next[104]), .E(n811), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFX1 \block_reg[5][103]  ( .D(block_next[103]), .E(n810), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFX1 \block_reg[5][102]  ( .D(block_next[102]), .E(n812), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFX1 \block_reg[5][101]  ( .D(block_next[101]), .E(n809), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFX1 \block_reg[5][100]  ( .D(block_next[100]), .E(n305), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFX1 \block_reg[5][99]  ( .D(block_next[99]), .E(n807), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFX1 \block_reg[5][98]  ( .D(block_next[98]), .E(n808), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFX1 \block_reg[5][97]  ( .D(block_next[97]), .E(n814), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFX1 \block_reg[5][96]  ( .D(block_next[96]), .E(n813), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFX1 \block_reg[5][89]  ( .D(block_next[89]), .E(n814), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFX1 \block_reg[5][88]  ( .D(block_next[88]), .E(n814), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFX1 \block_reg[5][87]  ( .D(block_next[87]), .E(n814), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFX1 \block_reg[5][86]  ( .D(block_next[86]), .E(n814), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFX1 \block_reg[5][85]  ( .D(block_next[85]), .E(n814), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFX1 \block_reg[5][84]  ( .D(block_next[84]), .E(n814), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFX1 \block_reg[5][83]  ( .D(block_next[83]), .E(n814), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFX1 \block_reg[5][82]  ( .D(block_next[82]), .E(n814), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFX1 \block_reg[5][81]  ( .D(block_next[81]), .E(n814), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFX1 \block_reg[5][80]  ( .D(block_next[80]), .E(n814), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFX1 \block_reg[5][79]  ( .D(block_next[79]), .E(n814), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFX1 \block_reg[5][78]  ( .D(block_next[78]), .E(n813), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFX1 \block_reg[5][77]  ( .D(block_next[77]), .E(n813), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFX1 \block_reg[5][76]  ( .D(block_next[76]), .E(n813), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFX1 \block_reg[5][75]  ( .D(block_next[75]), .E(n813), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFX1 \block_reg[5][74]  ( .D(block_next[74]), .E(n813), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFX1 \block_reg[5][73]  ( .D(block_next[73]), .E(n813), .CK(clk), .QN(n278) );
  EDFFX1 \block_reg[5][72]  ( .D(block_next[72]), .E(n813), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFX1 \block_reg[5][71]  ( .D(block_next[71]), .E(n813), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFX1 \block_reg[5][70]  ( .D(block_next[70]), .E(n813), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFX1 \block_reg[5][69]  ( .D(block_next[69]), .E(n813), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFX1 \block_reg[5][68]  ( .D(block_next[68]), .E(n813), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFX1 \block_reg[5][67]  ( .D(block_next[67]), .E(n813), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFX1 \block_reg[5][66]  ( .D(block_next[66]), .E(n813), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFX1 \block_reg[5][65]  ( .D(block_next[65]), .E(n812), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFX1 \block_reg[5][64]  ( .D(block_next[64]), .E(n812), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFX1 \block_reg[5][57]  ( .D(block_next[57]), .E(n812), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFX1 \block_reg[5][56]  ( .D(block_next[56]), .E(n812), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFX1 \block_reg[5][55]  ( .D(block_next[55]), .E(n812), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFX1 \block_reg[5][54]  ( .D(block_next[54]), .E(n812), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFX1 \block_reg[5][53]  ( .D(block_next[53]), .E(n812), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFX1 \block_reg[5][52]  ( .D(block_next[52]), .E(n811), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFX1 \block_reg[5][51]  ( .D(block_next[51]), .E(n811), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFX1 \block_reg[5][50]  ( .D(block_next[50]), .E(n811), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFX1 \block_reg[5][49]  ( .D(block_next[49]), .E(n811), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFX1 \block_reg[5][48]  ( .D(block_next[48]), .E(n811), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFX1 \block_reg[5][47]  ( .D(block_next[47]), .E(n811), .CK(clk), .QN(n286) );
  EDFFX1 \block_reg[5][46]  ( .D(block_next[46]), .E(n811), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFX1 \block_reg[5][45]  ( .D(block_next[45]), .E(n811), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFX1 \block_reg[5][44]  ( .D(block_next[44]), .E(n811), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFX1 \block_reg[5][43]  ( .D(block_next[43]), .E(n811), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFX1 \block_reg[5][42]  ( .D(block_next[42]), .E(n811), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n811), .CK(clk), .QN(n274) );
  EDFFX1 \block_reg[5][40]  ( .D(block_next[40]), .E(n811), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFX1 \block_reg[5][39]  ( .D(block_next[39]), .E(n810), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n810), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n810), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n810), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFX1 \block_reg[5][35]  ( .D(block_next[35]), .E(n810), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFX1 \block_reg[5][34]  ( .D(block_next[34]), .E(n810), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFX1 \block_reg[5][33]  ( .D(block_next[33]), .E(n810), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n810), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFX1 \block_reg[5][25]  ( .D(block_next[25]), .E(n809), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFX1 \block_reg[5][24]  ( .D(block_next[24]), .E(n809), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFX1 \block_reg[5][23]  ( .D(block_next[23]), .E(n809), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFX1 \block_reg[5][22]  ( .D(block_next[22]), .E(n809), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFX1 \block_reg[5][21]  ( .D(block_next[21]), .E(n809), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[5][20]  ( .D(block_next[20]), .E(n809), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFX1 \block_reg[5][19]  ( .D(block_next[19]), .E(n809), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFX1 \block_reg[5][18]  ( .D(block_next[18]), .E(n809), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFX1 \block_reg[5][17]  ( .D(block_next[17]), .E(n809), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFX1 \block_reg[5][16]  ( .D(block_next[16]), .E(n809), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFX1 \block_reg[5][15]  ( .D(block_next[15]), .E(n809), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[5][14]  ( .D(block_next[14]), .E(n809), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFX1 \block_reg[5][13]  ( .D(block_next[13]), .E(n808), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFX1 \block_reg[5][12]  ( .D(block_next[12]), .E(n808), .CK(clk), .QN(n298) );
  EDFFX1 \block_reg[5][11]  ( .D(block_next[11]), .E(n808), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFX1 \block_reg[5][10]  ( .D(block_next[10]), .E(n808), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFX1 \block_reg[5][9]  ( .D(block_next[9]), .E(n808), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFX1 \block_reg[5][8]  ( .D(block_next[8]), .E(n808), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFX1 \block_reg[5][7]  ( .D(block_next[7]), .E(n808), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFX1 \block_reg[5][6]  ( .D(block_next[6]), .E(n808), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFX1 \block_reg[5][5]  ( .D(block_next[5]), .E(n808), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFX1 \block_reg[5][4]  ( .D(block_next[4]), .E(n808), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFX1 \block_reg[5][3]  ( .D(block_next[3]), .E(n808), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFX1 \block_reg[5][2]  ( .D(block_next[2]), .E(n808), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFX1 \block_reg[5][1]  ( .D(block_next[1]), .E(n808), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFX1 \block_reg[5][0]  ( .D(block_next[0]), .E(n305), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFX1 \block_reg[1][121]  ( .D(block_next[121]), .E(n840), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFX1 \block_reg[1][120]  ( .D(block_next[120]), .E(n846), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFX1 \block_reg[1][119]  ( .D(block_next[119]), .E(n841), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFX1 \block_reg[1][118]  ( .D(block_next[118]), .E(n845), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFX1 \block_reg[1][117]  ( .D(block_next[117]), .E(n845), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFX1 \block_reg[1][116]  ( .D(block_next[116]), .E(n843), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFX1 \block_reg[1][115]  ( .D(block_next[115]), .E(n842), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFX1 \block_reg[1][114]  ( .D(block_next[114]), .E(n844), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFX1 \block_reg[1][113]  ( .D(block_next[113]), .E(n841), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFX1 \block_reg[1][112]  ( .D(block_next[112]), .E(n840), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFX1 \block_reg[1][111]  ( .D(block_next[111]), .E(n839), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFX1 \block_reg[1][110]  ( .D(block_next[110]), .E(n846), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFX1 \block_reg[1][109]  ( .D(block_next[109]), .E(n846), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFX1 \block_reg[1][108]  ( .D(block_next[108]), .E(n845), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFX1 \block_reg[1][107]  ( .D(block_next[107]), .E(n843), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFX1 \block_reg[1][106]  ( .D(block_next[106]), .E(n842), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFX1 \block_reg[1][105]  ( .D(block_next[105]), .E(n844), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFX1 \block_reg[1][104]  ( .D(block_next[104]), .E(n841), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFX1 \block_reg[1][103]  ( .D(block_next[103]), .E(n840), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFX1 \block_reg[1][102]  ( .D(block_next[102]), .E(n839), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFX1 \block_reg[1][101]  ( .D(block_next[101]), .E(n846), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFX1 \block_reg[1][100]  ( .D(block_next[100]), .E(n845), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFX1 \block_reg[1][99]  ( .D(block_next[99]), .E(n843), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFX1 \block_reg[1][98]  ( .D(block_next[98]), .E(n842), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFX1 \block_reg[1][97]  ( .D(block_next[97]), .E(n844), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFX1 \block_reg[1][96]  ( .D(block_next[96]), .E(n841), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFX1 \block_reg[1][89]  ( .D(block_next[89]), .E(n846), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFX1 \block_reg[1][88]  ( .D(block_next[88]), .E(n846), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFX1 \block_reg[1][87]  ( .D(block_next[87]), .E(n846), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFX1 \block_reg[1][86]  ( .D(block_next[86]), .E(n846), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFX1 \block_reg[1][85]  ( .D(block_next[85]), .E(n846), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFX1 \block_reg[1][84]  ( .D(block_next[84]), .E(n846), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFX1 \block_reg[1][83]  ( .D(block_next[83]), .E(n846), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFX1 \block_reg[1][82]  ( .D(block_next[82]), .E(n846), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFX1 \block_reg[1][81]  ( .D(block_next[81]), .E(n846), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFX1 \block_reg[1][80]  ( .D(block_next[80]), .E(n846), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFX1 \block_reg[1][79]  ( .D(block_next[79]), .E(n846), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFX1 \block_reg[1][78]  ( .D(block_next[78]), .E(n845), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFX1 \block_reg[1][77]  ( .D(block_next[77]), .E(n845), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFX1 \block_reg[1][76]  ( .D(block_next[76]), .E(n845), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFX1 \block_reg[1][75]  ( .D(block_next[75]), .E(n845), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFX1 \block_reg[1][74]  ( .D(block_next[74]), .E(n845), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFX1 \block_reg[1][73]  ( .D(block_next[73]), .E(n845), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFX1 \block_reg[1][72]  ( .D(block_next[72]), .E(n845), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFX1 \block_reg[1][71]  ( .D(block_next[71]), .E(n845), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFX1 \block_reg[1][70]  ( .D(block_next[70]), .E(n845), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFX1 \block_reg[1][69]  ( .D(block_next[69]), .E(n845), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFX1 \block_reg[1][68]  ( .D(block_next[68]), .E(n845), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFX1 \block_reg[1][67]  ( .D(block_next[67]), .E(n845), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFX1 \block_reg[1][66]  ( .D(block_next[66]), .E(n845), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFX1 \block_reg[1][65]  ( .D(block_next[65]), .E(n844), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFX1 \block_reg[1][64]  ( .D(block_next[64]), .E(n844), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[1][57]  ( .D(block_next[57]), .E(n844), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFX1 \block_reg[1][56]  ( .D(block_next[56]), .E(n844), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFX1 \block_reg[1][55]  ( .D(block_next[55]), .E(n844), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFX1 \block_reg[1][54]  ( .D(block_next[54]), .E(n844), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n844), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n843), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[1][51]  ( .D(block_next[51]), .E(n843), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFX1 \block_reg[1][50]  ( .D(block_next[50]), .E(n843), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n843), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[1][48]  ( .D(block_next[48]), .E(n843), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFX1 \block_reg[1][47]  ( .D(block_next[47]), .E(n843), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFX1 \block_reg[1][46]  ( .D(block_next[46]), .E(n843), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFX1 \block_reg[1][45]  ( .D(block_next[45]), .E(n843), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFX1 \block_reg[1][44]  ( .D(block_next[44]), .E(n843), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFX1 \block_reg[1][43]  ( .D(block_next[43]), .E(n843), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFX1 \block_reg[1][42]  ( .D(block_next[42]), .E(n843), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFX1 \block_reg[1][41]  ( .D(block_next[41]), .E(n843), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[1][40]  ( .D(block_next[40]), .E(n843), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFX1 \block_reg[1][39]  ( .D(block_next[39]), .E(n842), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFX1 \block_reg[1][38]  ( .D(block_next[38]), .E(n842), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFX1 \block_reg[1][37]  ( .D(block_next[37]), .E(n842), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[1][36]  ( .D(block_next[36]), .E(n842), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(n842), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFX1 \block_reg[1][34]  ( .D(block_next[34]), .E(n842), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFX1 \block_reg[1][33]  ( .D(block_next[33]), .E(n842), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFX1 \block_reg[1][32]  ( .D(block_next[32]), .E(n842), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[1][25]  ( .D(block_next[25]), .E(n841), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFX1 \block_reg[1][24]  ( .D(block_next[24]), .E(n841), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFX1 \block_reg[1][23]  ( .D(block_next[23]), .E(n841), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFX1 \block_reg[1][22]  ( .D(block_next[22]), .E(n841), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFX1 \block_reg[1][21]  ( .D(block_next[21]), .E(n841), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n841), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFX1 \block_reg[1][19]  ( .D(block_next[19]), .E(n841), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFX1 \block_reg[1][18]  ( .D(block_next[18]), .E(n841), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFX1 \block_reg[1][17]  ( .D(block_next[17]), .E(n841), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFX1 \block_reg[1][16]  ( .D(block_next[16]), .E(n841), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFX1 \block_reg[1][15]  ( .D(block_next[15]), .E(n841), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFX1 \block_reg[1][14]  ( .D(block_next[14]), .E(n841), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFX1 \block_reg[1][13]  ( .D(block_next[13]), .E(n839), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFX1 \block_reg[1][12]  ( .D(block_next[12]), .E(n846), .CK(clk), .QN(n294) );
  EDFFX1 \block_reg[1][11]  ( .D(block_next[11]), .E(n304), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFX1 \block_reg[1][10]  ( .D(block_next[10]), .E(n845), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFX1 \block_reg[1][9]  ( .D(block_next[9]), .E(n843), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFX1 \block_reg[1][8]  ( .D(block_next[8]), .E(n842), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFX1 \block_reg[1][7]  ( .D(block_next[7]), .E(n844), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFX1 \block_reg[1][6]  ( .D(block_next[6]), .E(n841), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFX1 \block_reg[1][5]  ( .D(block_next[5]), .E(n304), .CK(clk), .Q(
        \block[1][5] ) );
  EDFFX1 \block_reg[1][4]  ( .D(block_next[4]), .E(n840), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFX1 \block_reg[1][3]  ( .D(block_next[3]), .E(n839), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFX1 \block_reg[1][2]  ( .D(block_next[2]), .E(n840), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFX1 \block_reg[1][1]  ( .D(block_next[1]), .E(n839), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFX1 \block_reg[1][0]  ( .D(block_next[0]), .E(n840), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFX1 \block_reg[4][121]  ( .D(block_next[121]), .E(n819), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFX1 \block_reg[4][120]  ( .D(block_next[120]), .E(n819), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFX1 \block_reg[4][119]  ( .D(block_next[119]), .E(n818), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFX1 \block_reg[4][118]  ( .D(block_next[118]), .E(n820), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFX1 \block_reg[4][117]  ( .D(block_next[117]), .E(n815), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFX1 \block_reg[4][116]  ( .D(block_next[116]), .E(n816), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFX1 \block_reg[4][115]  ( .D(block_next[115]), .E(n821), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFX1 \block_reg[4][114]  ( .D(block_next[114]), .E(n820), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFX1 \block_reg[4][113]  ( .D(block_next[113]), .E(n818), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFX1 \block_reg[4][112]  ( .D(block_next[112]), .E(n819), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFX1 \block_reg[4][111]  ( .D(block_next[111]), .E(n816), .CK(clk), .QN(
        n289) );
  EDFFX1 \block_reg[4][110]  ( .D(block_next[110]), .E(n820), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFX1 \block_reg[4][109]  ( .D(block_next[109]), .E(n311), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFX1 \block_reg[4][108]  ( .D(block_next[108]), .E(n822), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFX1 \block_reg[4][107]  ( .D(block_next[107]), .E(n817), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFX1 \block_reg[4][106]  ( .D(block_next[106]), .E(n815), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFX1 \block_reg[4][105]  ( .D(block_next[105]), .E(n821), .CK(clk), .QN(
        n281) );
  EDFFX1 \block_reg[4][104]  ( .D(block_next[104]), .E(n822), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFX1 \block_reg[4][103]  ( .D(block_next[103]), .E(n822), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFX1 \block_reg[4][102]  ( .D(block_next[102]), .E(n822), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFX1 \block_reg[4][101]  ( .D(block_next[101]), .E(n822), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFX1 \block_reg[4][100]  ( .D(block_next[100]), .E(n822), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFX1 \block_reg[4][99]  ( .D(block_next[99]), .E(n822), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFX1 \block_reg[4][98]  ( .D(block_next[98]), .E(n822), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFX1 \block_reg[4][97]  ( .D(block_next[97]), .E(n822), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFX1 \block_reg[4][96]  ( .D(block_next[96]), .E(n822), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFX1 \block_reg[4][89]  ( .D(block_next[89]), .E(n821), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFX1 \block_reg[4][88]  ( .D(block_next[88]), .E(n821), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFX1 \block_reg[4][87]  ( .D(block_next[87]), .E(n821), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFX1 \block_reg[4][86]  ( .D(block_next[86]), .E(n821), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFX1 \block_reg[4][85]  ( .D(block_next[85]), .E(n821), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFX1 \block_reg[4][84]  ( .D(block_next[84]), .E(n821), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFX1 \block_reg[4][83]  ( .D(block_next[83]), .E(n821), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFX1 \block_reg[4][82]  ( .D(block_next[82]), .E(n821), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFX1 \block_reg[4][81]  ( .D(block_next[81]), .E(n821), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFX1 \block_reg[4][80]  ( .D(block_next[80]), .E(n821), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFX1 \block_reg[4][79]  ( .D(block_next[79]), .E(n821), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFX1 \block_reg[4][78]  ( .D(block_next[78]), .E(n816), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFX1 \block_reg[4][77]  ( .D(block_next[77]), .E(n815), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFX1 \block_reg[4][76]  ( .D(block_next[76]), .E(n817), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFX1 \block_reg[4][75]  ( .D(block_next[75]), .E(n822), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFX1 \block_reg[4][74]  ( .D(block_next[74]), .E(n311), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFX1 \block_reg[4][73]  ( .D(block_next[73]), .E(n822), .CK(clk), .QN(n277) );
  EDFFX1 \block_reg[4][72]  ( .D(block_next[72]), .E(n819), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFX1 \block_reg[4][71]  ( .D(block_next[71]), .E(n818), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFX1 \block_reg[4][70]  ( .D(block_next[70]), .E(n820), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFX1 \block_reg[4][69]  ( .D(block_next[69]), .E(n821), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFX1 \block_reg[4][68]  ( .D(block_next[68]), .E(n816), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFX1 \block_reg[4][67]  ( .D(block_next[67]), .E(n815), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFX1 \block_reg[4][66]  ( .D(block_next[66]), .E(n817), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFX1 \block_reg[4][65]  ( .D(block_next[65]), .E(n820), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFX1 \block_reg[4][64]  ( .D(block_next[64]), .E(n820), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFX1 \block_reg[4][57]  ( .D(block_next[57]), .E(n820), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFX1 \block_reg[4][56]  ( .D(block_next[56]), .E(n820), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFX1 \block_reg[4][55]  ( .D(block_next[55]), .E(n820), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFX1 \block_reg[4][54]  ( .D(block_next[54]), .E(n820), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n820), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n819), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[4][51]  ( .D(block_next[51]), .E(n819), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFX1 \block_reg[4][50]  ( .D(block_next[50]), .E(n819), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n819), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[4][48]  ( .D(block_next[48]), .E(n819), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFX1 \block_reg[4][47]  ( .D(block_next[47]), .E(n819), .CK(clk), .QN(n285) );
  EDFFX1 \block_reg[4][46]  ( .D(block_next[46]), .E(n819), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFX1 \block_reg[4][45]  ( .D(block_next[45]), .E(n819), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFX1 \block_reg[4][44]  ( .D(block_next[44]), .E(n819), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFX1 \block_reg[4][43]  ( .D(block_next[43]), .E(n819), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFX1 \block_reg[4][42]  ( .D(block_next[42]), .E(n819), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n819), .CK(clk), .QN(n273) );
  EDFFX1 \block_reg[4][40]  ( .D(block_next[40]), .E(n819), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFX1 \block_reg[4][39]  ( .D(block_next[39]), .E(n818), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n818), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n818), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n818), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n818), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFX1 \block_reg[4][34]  ( .D(block_next[34]), .E(n818), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFX1 \block_reg[4][33]  ( .D(block_next[33]), .E(n818), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n818), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[4][25]  ( .D(block_next[25]), .E(n311), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFX1 \block_reg[4][24]  ( .D(block_next[24]), .E(n311), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFX1 \block_reg[4][23]  ( .D(block_next[23]), .E(n311), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFX1 \block_reg[4][22]  ( .D(block_next[22]), .E(n818), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFX1 \block_reg[4][21]  ( .D(block_next[21]), .E(n819), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n818), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFX1 \block_reg[4][19]  ( .D(block_next[19]), .E(n820), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFX1 \block_reg[4][18]  ( .D(block_next[18]), .E(n821), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFX1 \block_reg[4][17]  ( .D(block_next[17]), .E(n816), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFX1 \block_reg[4][16]  ( .D(block_next[16]), .E(n815), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFX1 \block_reg[4][15]  ( .D(block_next[15]), .E(n817), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFX1 \block_reg[4][14]  ( .D(block_next[14]), .E(n822), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFX1 \block_reg[4][13]  ( .D(block_next[13]), .E(n817), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFX1 \block_reg[4][12]  ( .D(block_next[12]), .E(n817), .CK(clk), .QN(n297) );
  EDFFX1 \block_reg[4][11]  ( .D(block_next[11]), .E(n817), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFX1 \block_reg[4][10]  ( .D(block_next[10]), .E(n817), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFX1 \block_reg[4][9]  ( .D(block_next[9]), .E(n817), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFX1 \block_reg[4][8]  ( .D(block_next[8]), .E(n817), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFX1 \block_reg[4][7]  ( .D(block_next[7]), .E(n817), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFX1 \block_reg[4][6]  ( .D(block_next[6]), .E(n817), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFX1 \block_reg[4][5]  ( .D(block_next[5]), .E(n817), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFX1 \block_reg[4][4]  ( .D(block_next[4]), .E(n817), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFX1 \block_reg[4][3]  ( .D(block_next[3]), .E(n817), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFX1 \block_reg[4][2]  ( .D(block_next[2]), .E(n817), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFX1 \block_reg[4][1]  ( .D(block_next[1]), .E(n817), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFX1 \block_reg[4][0]  ( .D(block_next[0]), .E(n816), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFX1 \block_reg[0][121]  ( .D(block_next[121]), .E(n854), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFX1 \block_reg[0][120]  ( .D(block_next[120]), .E(n854), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFX1 \block_reg[0][119]  ( .D(block_next[119]), .E(n852), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFX1 \block_reg[0][118]  ( .D(block_next[118]), .E(n853), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFX1 \block_reg[0][117]  ( .D(block_next[117]), .E(n847), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFX1 \block_reg[0][116]  ( .D(block_next[116]), .E(n849), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFX1 \block_reg[0][115]  ( .D(block_next[115]), .E(n850), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFX1 \block_reg[0][114]  ( .D(block_next[114]), .E(n852), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFX1 \block_reg[0][113]  ( .D(block_next[113]), .E(n851), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFX1 \block_reg[0][112]  ( .D(block_next[112]), .E(n310), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFX1 \block_reg[0][111]  ( .D(block_next[111]), .E(n848), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFX1 \block_reg[0][110]  ( .D(block_next[110]), .E(n854), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFX1 \block_reg[0][109]  ( .D(block_next[109]), .E(n853), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFX1 \block_reg[0][108]  ( .D(block_next[108]), .E(n848), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFX1 \block_reg[0][107]  ( .D(block_next[107]), .E(n847), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFX1 \block_reg[0][106]  ( .D(block_next[106]), .E(n849), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFX1 \block_reg[0][105]  ( .D(block_next[105]), .E(n850), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFX1 \block_reg[0][104]  ( .D(block_next[104]), .E(n849), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFX1 \block_reg[0][103]  ( .D(block_next[103]), .E(n850), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFX1 \block_reg[0][102]  ( .D(block_next[102]), .E(n852), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFX1 \block_reg[0][101]  ( .D(block_next[101]), .E(n851), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFX1 \block_reg[0][100]  ( .D(block_next[100]), .E(n310), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFX1 \block_reg[0][99]  ( .D(block_next[99]), .E(n854), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFX1 \block_reg[0][98]  ( .D(block_next[98]), .E(n853), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFX1 \block_reg[0][97]  ( .D(block_next[97]), .E(n848), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFX1 \block_reg[0][96]  ( .D(block_next[96]), .E(n847), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFX1 \block_reg[0][89]  ( .D(block_next[89]), .E(n854), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFX1 \block_reg[0][88]  ( .D(block_next[88]), .E(n854), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFX1 \block_reg[0][87]  ( .D(block_next[87]), .E(n854), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFX1 \block_reg[0][86]  ( .D(block_next[86]), .E(n854), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFX1 \block_reg[0][85]  ( .D(block_next[85]), .E(n854), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFX1 \block_reg[0][84]  ( .D(block_next[84]), .E(n854), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFX1 \block_reg[0][83]  ( .D(block_next[83]), .E(n854), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFX1 \block_reg[0][82]  ( .D(block_next[82]), .E(n854), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFX1 \block_reg[0][81]  ( .D(block_next[81]), .E(n854), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFX1 \block_reg[0][80]  ( .D(block_next[80]), .E(n854), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFX1 \block_reg[0][79]  ( .D(block_next[79]), .E(n854), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFX1 \block_reg[0][78]  ( .D(block_next[78]), .E(n853), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFX1 \block_reg[0][77]  ( .D(block_next[77]), .E(n853), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFX1 \block_reg[0][76]  ( .D(block_next[76]), .E(n853), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFX1 \block_reg[0][75]  ( .D(block_next[75]), .E(n853), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFX1 \block_reg[0][74]  ( .D(block_next[74]), .E(n853), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFX1 \block_reg[0][73]  ( .D(block_next[73]), .E(n853), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFX1 \block_reg[0][72]  ( .D(block_next[72]), .E(n853), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFX1 \block_reg[0][71]  ( .D(block_next[71]), .E(n853), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFX1 \block_reg[0][70]  ( .D(block_next[70]), .E(n853), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFX1 \block_reg[0][69]  ( .D(block_next[69]), .E(n853), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFX1 \block_reg[0][68]  ( .D(block_next[68]), .E(n853), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFX1 \block_reg[0][67]  ( .D(block_next[67]), .E(n853), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFX1 \block_reg[0][66]  ( .D(block_next[66]), .E(n853), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFX1 \block_reg[0][65]  ( .D(block_next[65]), .E(n852), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFX1 \block_reg[0][64]  ( .D(block_next[64]), .E(n852), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[0][57]  ( .D(block_next[57]), .E(n852), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFX1 \block_reg[0][56]  ( .D(block_next[56]), .E(n852), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFX1 \block_reg[0][55]  ( .D(block_next[55]), .E(n852), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFX1 \block_reg[0][54]  ( .D(block_next[54]), .E(n852), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n852), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n851), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[0][51]  ( .D(block_next[51]), .E(n851), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFX1 \block_reg[0][50]  ( .D(block_next[50]), .E(n851), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n851), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[0][48]  ( .D(block_next[48]), .E(n851), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFX1 \block_reg[0][47]  ( .D(block_next[47]), .E(n851), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFX1 \block_reg[0][46]  ( .D(block_next[46]), .E(n851), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFX1 \block_reg[0][45]  ( .D(block_next[45]), .E(n851), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFX1 \block_reg[0][44]  ( .D(block_next[44]), .E(n851), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFX1 \block_reg[0][43]  ( .D(block_next[43]), .E(n851), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFX1 \block_reg[0][42]  ( .D(block_next[42]), .E(n851), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n851), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[0][40]  ( .D(block_next[40]), .E(n851), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFX1 \block_reg[0][39]  ( .D(block_next[39]), .E(n850), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n850), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n850), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n850), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n850), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[0][34]  ( .D(block_next[34]), .E(n850), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFX1 \block_reg[0][33]  ( .D(block_next[33]), .E(n850), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n850), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[0][25]  ( .D(block_next[25]), .E(n310), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFX1 \block_reg[0][24]  ( .D(block_next[24]), .E(n310), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFX1 \block_reg[0][23]  ( .D(block_next[23]), .E(n310), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFX1 \block_reg[0][22]  ( .D(block_next[22]), .E(n853), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFX1 \block_reg[0][21]  ( .D(block_next[21]), .E(n854), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n851), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFX1 \block_reg[0][19]  ( .D(block_next[19]), .E(n853), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFX1 \block_reg[0][18]  ( .D(block_next[18]), .E(n848), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFX1 \block_reg[0][17]  ( .D(block_next[17]), .E(n847), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFX1 \block_reg[0][16]  ( .D(block_next[16]), .E(n849), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFX1 \block_reg[0][15]  ( .D(block_next[15]), .E(n850), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFX1 \block_reg[0][14]  ( .D(block_next[14]), .E(n852), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFX1 \block_reg[0][13]  ( .D(block_next[13]), .E(n849), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFX1 \block_reg[0][12]  ( .D(block_next[12]), .E(n849), .CK(clk), .QN(n293) );
  EDFFX1 \block_reg[0][11]  ( .D(block_next[11]), .E(n849), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFX1 \block_reg[0][10]  ( .D(block_next[10]), .E(n849), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFX1 \block_reg[0][9]  ( .D(block_next[9]), .E(n849), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFX1 \block_reg[0][8]  ( .D(block_next[8]), .E(n849), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFX1 \block_reg[0][7]  ( .D(block_next[7]), .E(n849), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFX1 \block_reg[0][6]  ( .D(block_next[6]), .E(n849), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFX1 \block_reg[0][5]  ( .D(block_next[5]), .E(n849), .CK(clk), .Q(
        \block[0][5] ) );
  EDFFX1 \block_reg[0][4]  ( .D(block_next[4]), .E(n849), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFX1 \block_reg[0][3]  ( .D(block_next[3]), .E(n849), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFX1 \block_reg[0][2]  ( .D(block_next[2]), .E(n849), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFX1 \block_reg[0][1]  ( .D(block_next[1]), .E(n849), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFX1 \block_reg[0][0]  ( .D(block_next[0]), .E(n848), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFX1 \block_reg[6][121]  ( .D(block_next[121]), .E(n803), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFX1 \block_reg[6][120]  ( .D(block_next[120]), .E(n803), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFX1 \block_reg[6][119]  ( .D(block_next[119]), .E(n802), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFX1 \block_reg[6][118]  ( .D(block_next[118]), .E(n804), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFX1 \block_reg[6][117]  ( .D(block_next[117]), .E(n799), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFX1 \block_reg[6][116]  ( .D(block_next[116]), .E(n800), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFX1 \block_reg[6][115]  ( .D(block_next[115]), .E(n805), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFX1 \block_reg[6][114]  ( .D(block_next[114]), .E(n804), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFX1 \block_reg[6][113]  ( .D(block_next[113]), .E(n802), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFX1 \block_reg[6][112]  ( .D(block_next[112]), .E(n803), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFX1 \block_reg[6][111]  ( .D(block_next[111]), .E(n800), .CK(clk), .QN(
        n291) );
  EDFFX1 \block_reg[6][110]  ( .D(block_next[110]), .E(n804), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFX1 \block_reg[6][109]  ( .D(block_next[109]), .E(n316), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFX1 \block_reg[6][108]  ( .D(block_next[108]), .E(n806), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFX1 \block_reg[6][107]  ( .D(block_next[107]), .E(n801), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFX1 \block_reg[6][106]  ( .D(block_next[106]), .E(n799), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFX1 \block_reg[6][105]  ( .D(block_next[105]), .E(n805), .CK(clk), .QN(
        n283) );
  EDFFX1 \block_reg[6][104]  ( .D(block_next[104]), .E(n806), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFX1 \block_reg[6][103]  ( .D(block_next[103]), .E(n806), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFX1 \block_reg[6][102]  ( .D(block_next[102]), .E(n806), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFX1 \block_reg[6][101]  ( .D(block_next[101]), .E(n806), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFX1 \block_reg[6][100]  ( .D(block_next[100]), .E(n806), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFX1 \block_reg[6][99]  ( .D(block_next[99]), .E(n806), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFX1 \block_reg[6][98]  ( .D(block_next[98]), .E(n806), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFX1 \block_reg[6][97]  ( .D(block_next[97]), .E(n806), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFX1 \block_reg[6][96]  ( .D(block_next[96]), .E(n806), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFX1 \block_reg[6][89]  ( .D(block_next[89]), .E(n805), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFX1 \block_reg[6][88]  ( .D(block_next[88]), .E(n805), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFX1 \block_reg[6][87]  ( .D(block_next[87]), .E(n805), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFX1 \block_reg[6][86]  ( .D(block_next[86]), .E(n805), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFX1 \block_reg[6][85]  ( .D(block_next[85]), .E(n805), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFX1 \block_reg[6][84]  ( .D(block_next[84]), .E(n805), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFX1 \block_reg[6][83]  ( .D(block_next[83]), .E(n805), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFX1 \block_reg[6][82]  ( .D(block_next[82]), .E(n805), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFX1 \block_reg[6][81]  ( .D(block_next[81]), .E(n805), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFX1 \block_reg[6][80]  ( .D(block_next[80]), .E(n805), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFX1 \block_reg[6][79]  ( .D(block_next[79]), .E(n805), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFX1 \block_reg[6][78]  ( .D(block_next[78]), .E(n800), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFX1 \block_reg[6][77]  ( .D(block_next[77]), .E(n799), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFX1 \block_reg[6][76]  ( .D(block_next[76]), .E(n801), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFX1 \block_reg[6][75]  ( .D(block_next[75]), .E(n806), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFX1 \block_reg[6][74]  ( .D(block_next[74]), .E(n316), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFX1 \block_reg[6][73]  ( .D(block_next[73]), .E(n806), .CK(clk), .QN(n279) );
  EDFFX1 \block_reg[6][72]  ( .D(block_next[72]), .E(n803), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFX1 \block_reg[6][71]  ( .D(block_next[71]), .E(n802), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFX1 \block_reg[6][70]  ( .D(block_next[70]), .E(n804), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFX1 \block_reg[6][69]  ( .D(block_next[69]), .E(n805), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFX1 \block_reg[6][68]  ( .D(block_next[68]), .E(n800), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFX1 \block_reg[6][67]  ( .D(block_next[67]), .E(n799), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFX1 \block_reg[6][66]  ( .D(block_next[66]), .E(n801), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFX1 \block_reg[6][65]  ( .D(block_next[65]), .E(n804), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFX1 \block_reg[6][64]  ( .D(block_next[64]), .E(n804), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFX1 \block_reg[6][57]  ( .D(block_next[57]), .E(n804), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFX1 \block_reg[6][56]  ( .D(block_next[56]), .E(n804), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFX1 \block_reg[6][55]  ( .D(block_next[55]), .E(n804), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFX1 \block_reg[6][54]  ( .D(block_next[54]), .E(n804), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n804), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n803), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[6][51]  ( .D(block_next[51]), .E(n803), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFX1 \block_reg[6][50]  ( .D(block_next[50]), .E(n803), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFX1 \block_reg[6][49]  ( .D(block_next[49]), .E(n803), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFX1 \block_reg[6][48]  ( .D(block_next[48]), .E(n803), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFX1 \block_reg[6][47]  ( .D(block_next[47]), .E(n803), .CK(clk), .QN(n287) );
  EDFFX1 \block_reg[6][46]  ( .D(block_next[46]), .E(n803), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFX1 \block_reg[6][45]  ( .D(block_next[45]), .E(n803), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFX1 \block_reg[6][44]  ( .D(block_next[44]), .E(n803), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFX1 \block_reg[6][43]  ( .D(block_next[43]), .E(n803), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFX1 \block_reg[6][42]  ( .D(block_next[42]), .E(n803), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n803), .CK(clk), .QN(n275) );
  EDFFX1 \block_reg[6][40]  ( .D(block_next[40]), .E(n803), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFX1 \block_reg[6][39]  ( .D(block_next[39]), .E(n802), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n802), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n802), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n802), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n802), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFX1 \block_reg[6][34]  ( .D(block_next[34]), .E(n802), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFX1 \block_reg[6][33]  ( .D(block_next[33]), .E(n802), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n802), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[6][25]  ( .D(block_next[25]), .E(n316), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFX1 \block_reg[6][24]  ( .D(block_next[24]), .E(n316), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFX1 \block_reg[6][23]  ( .D(block_next[23]), .E(n316), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFX1 \block_reg[6][22]  ( .D(block_next[22]), .E(n802), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFX1 \block_reg[6][21]  ( .D(block_next[21]), .E(n803), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n802), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFX1 \block_reg[6][19]  ( .D(block_next[19]), .E(n804), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFX1 \block_reg[6][18]  ( .D(block_next[18]), .E(n805), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFX1 \block_reg[6][17]  ( .D(block_next[17]), .E(n800), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFX1 \block_reg[6][16]  ( .D(block_next[16]), .E(n799), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFX1 \block_reg[6][15]  ( .D(block_next[15]), .E(n801), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFX1 \block_reg[6][14]  ( .D(block_next[14]), .E(n806), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFX1 \block_reg[6][13]  ( .D(block_next[13]), .E(n801), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFX1 \block_reg[6][12]  ( .D(block_next[12]), .E(n801), .CK(clk), .QN(n299) );
  EDFFX1 \block_reg[6][11]  ( .D(block_next[11]), .E(n801), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFX1 \block_reg[6][10]  ( .D(block_next[10]), .E(n801), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFX1 \block_reg[6][9]  ( .D(block_next[9]), .E(n801), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFX1 \block_reg[6][8]  ( .D(block_next[8]), .E(n801), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFX1 \block_reg[6][7]  ( .D(block_next[7]), .E(n801), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFX1 \block_reg[6][6]  ( .D(block_next[6]), .E(n801), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFX1 \block_reg[6][5]  ( .D(block_next[5]), .E(n801), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFX1 \block_reg[6][4]  ( .D(block_next[4]), .E(n801), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFX1 \block_reg[6][3]  ( .D(block_next[3]), .E(n801), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFX1 \block_reg[6][2]  ( .D(block_next[2]), .E(n801), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFX1 \block_reg[6][1]  ( .D(block_next[1]), .E(n801), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFX1 \block_reg[6][0]  ( .D(block_next[0]), .E(n800), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFX1 \block_reg[2][121]  ( .D(block_next[121]), .E(n838), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFX1 \block_reg[2][120]  ( .D(block_next[120]), .E(n838), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFX1 \block_reg[2][119]  ( .D(block_next[119]), .E(n836), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFX1 \block_reg[2][118]  ( .D(block_next[118]), .E(n837), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFX1 \block_reg[2][117]  ( .D(block_next[117]), .E(n831), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFX1 \block_reg[2][116]  ( .D(block_next[116]), .E(n833), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFX1 \block_reg[2][115]  ( .D(block_next[115]), .E(n834), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFX1 \block_reg[2][114]  ( .D(block_next[114]), .E(n836), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFX1 \block_reg[2][113]  ( .D(block_next[113]), .E(n835), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFX1 \block_reg[2][112]  ( .D(block_next[112]), .E(n315), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFX1 \block_reg[2][111]  ( .D(block_next[111]), .E(n832), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFX1 \block_reg[2][110]  ( .D(block_next[110]), .E(n838), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFX1 \block_reg[2][109]  ( .D(block_next[109]), .E(n837), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFX1 \block_reg[2][108]  ( .D(block_next[108]), .E(n832), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFX1 \block_reg[2][107]  ( .D(block_next[107]), .E(n831), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFX1 \block_reg[2][106]  ( .D(block_next[106]), .E(n833), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFX1 \block_reg[2][105]  ( .D(block_next[105]), .E(n834), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFX1 \block_reg[2][104]  ( .D(block_next[104]), .E(n833), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFX1 \block_reg[2][103]  ( .D(block_next[103]), .E(n834), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFX1 \block_reg[2][102]  ( .D(block_next[102]), .E(n836), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFX1 \block_reg[2][101]  ( .D(block_next[101]), .E(n835), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFX1 \block_reg[2][100]  ( .D(block_next[100]), .E(n315), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFX1 \block_reg[2][99]  ( .D(block_next[99]), .E(n838), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFX1 \block_reg[2][98]  ( .D(block_next[98]), .E(n837), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFX1 \block_reg[2][97]  ( .D(block_next[97]), .E(n832), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFX1 \block_reg[2][96]  ( .D(block_next[96]), .E(n831), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFX1 \block_reg[2][89]  ( .D(block_next[89]), .E(n838), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFX1 \block_reg[2][88]  ( .D(block_next[88]), .E(n838), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFX1 \block_reg[2][87]  ( .D(block_next[87]), .E(n838), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFX1 \block_reg[2][86]  ( .D(block_next[86]), .E(n838), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFX1 \block_reg[2][85]  ( .D(block_next[85]), .E(n838), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFX1 \block_reg[2][84]  ( .D(block_next[84]), .E(n838), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFX1 \block_reg[2][83]  ( .D(block_next[83]), .E(n838), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFX1 \block_reg[2][82]  ( .D(block_next[82]), .E(n838), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFX1 \block_reg[2][81]  ( .D(block_next[81]), .E(n838), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFX1 \block_reg[2][80]  ( .D(block_next[80]), .E(n838), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFX1 \block_reg[2][79]  ( .D(block_next[79]), .E(n838), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFX1 \block_reg[2][78]  ( .D(block_next[78]), .E(n837), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFX1 \block_reg[2][77]  ( .D(block_next[77]), .E(n837), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFX1 \block_reg[2][76]  ( .D(block_next[76]), .E(n837), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFX1 \block_reg[2][75]  ( .D(block_next[75]), .E(n837), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFX1 \block_reg[2][74]  ( .D(block_next[74]), .E(n837), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFX1 \block_reg[2][73]  ( .D(block_next[73]), .E(n837), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFX1 \block_reg[2][72]  ( .D(block_next[72]), .E(n837), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFX1 \block_reg[2][71]  ( .D(block_next[71]), .E(n837), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFX1 \block_reg[2][70]  ( .D(block_next[70]), .E(n837), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFX1 \block_reg[2][69]  ( .D(block_next[69]), .E(n837), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFX1 \block_reg[2][68]  ( .D(block_next[68]), .E(n837), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFX1 \block_reg[2][67]  ( .D(block_next[67]), .E(n837), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFX1 \block_reg[2][66]  ( .D(block_next[66]), .E(n837), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFX1 \block_reg[2][65]  ( .D(block_next[65]), .E(n836), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFX1 \block_reg[2][64]  ( .D(block_next[64]), .E(n836), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFX1 \block_reg[2][57]  ( .D(block_next[57]), .E(n836), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFX1 \block_reg[2][56]  ( .D(block_next[56]), .E(n836), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFX1 \block_reg[2][55]  ( .D(block_next[55]), .E(n836), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFX1 \block_reg[2][54]  ( .D(block_next[54]), .E(n836), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFX1 \block_reg[2][53]  ( .D(block_next[53]), .E(n836), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFX1 \block_reg[2][52]  ( .D(block_next[52]), .E(n835), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFX1 \block_reg[2][51]  ( .D(block_next[51]), .E(n835), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFX1 \block_reg[2][50]  ( .D(block_next[50]), .E(n835), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFX1 \block_reg[2][49]  ( .D(block_next[49]), .E(n835), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFX1 \block_reg[2][48]  ( .D(block_next[48]), .E(n835), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFX1 \block_reg[2][47]  ( .D(block_next[47]), .E(n835), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFX1 \block_reg[2][46]  ( .D(block_next[46]), .E(n835), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFX1 \block_reg[2][45]  ( .D(block_next[45]), .E(n835), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFX1 \block_reg[2][44]  ( .D(block_next[44]), .E(n835), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFX1 \block_reg[2][43]  ( .D(block_next[43]), .E(n835), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFX1 \block_reg[2][42]  ( .D(block_next[42]), .E(n835), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFX1 \block_reg[2][41]  ( .D(block_next[41]), .E(n835), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFX1 \block_reg[2][40]  ( .D(block_next[40]), .E(n835), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFX1 \block_reg[2][39]  ( .D(block_next[39]), .E(n834), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFX1 \block_reg[2][38]  ( .D(block_next[38]), .E(n834), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFX1 \block_reg[2][37]  ( .D(block_next[37]), .E(n834), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFX1 \block_reg[2][36]  ( .D(block_next[36]), .E(n834), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFX1 \block_reg[2][35]  ( .D(block_next[35]), .E(n834), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFX1 \block_reg[2][34]  ( .D(block_next[34]), .E(n834), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFX1 \block_reg[2][33]  ( .D(block_next[33]), .E(n834), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFX1 \block_reg[2][32]  ( .D(block_next[32]), .E(n834), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFX1 \block_reg[2][25]  ( .D(block_next[25]), .E(n315), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFX1 \block_reg[2][24]  ( .D(block_next[24]), .E(n315), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFX1 \block_reg[2][23]  ( .D(block_next[23]), .E(n315), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFX1 \block_reg[2][22]  ( .D(block_next[22]), .E(n837), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFX1 \block_reg[2][21]  ( .D(block_next[21]), .E(n838), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFX1 \block_reg[2][20]  ( .D(block_next[20]), .E(n835), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFX1 \block_reg[2][19]  ( .D(block_next[19]), .E(n837), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFX1 \block_reg[2][18]  ( .D(block_next[18]), .E(n832), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFX1 \block_reg[2][17]  ( .D(block_next[17]), .E(n831), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFX1 \block_reg[2][16]  ( .D(block_next[16]), .E(n833), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFX1 \block_reg[2][15]  ( .D(block_next[15]), .E(n834), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFX1 \block_reg[2][14]  ( .D(block_next[14]), .E(n836), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFX1 \block_reg[2][13]  ( .D(block_next[13]), .E(n833), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFX1 \block_reg[2][12]  ( .D(block_next[12]), .E(n833), .CK(clk), .QN(n295) );
  EDFFX1 \block_reg[2][11]  ( .D(block_next[11]), .E(n833), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFX1 \block_reg[2][10]  ( .D(block_next[10]), .E(n833), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFX1 \block_reg[2][9]  ( .D(block_next[9]), .E(n833), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFX1 \block_reg[2][8]  ( .D(block_next[8]), .E(n833), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFX1 \block_reg[2][7]  ( .D(block_next[7]), .E(n833), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFX1 \block_reg[2][6]  ( .D(block_next[6]), .E(n833), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFX1 \block_reg[2][5]  ( .D(block_next[5]), .E(n833), .CK(clk), .Q(
        \block[2][5] ) );
  EDFFX1 \block_reg[2][4]  ( .D(block_next[4]), .E(n833), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFX1 \block_reg[2][3]  ( .D(block_next[3]), .E(n833), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFX1 \block_reg[2][2]  ( .D(block_next[2]), .E(n833), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFX1 \block_reg[2][1]  ( .D(block_next[1]), .E(n833), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFX1 \block_reg[2][0]  ( .D(block_next[0]), .E(n832), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFX1 \block_reg[7][127]  ( .D(block_next[127]), .E(n796), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFX1 \block_reg[7][126]  ( .D(block_next[126]), .E(n797), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFX1 \block_reg[7][125]  ( .D(block_next[125]), .E(n795), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFX1 \block_reg[7][124]  ( .D(block_next[124]), .E(n794), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFX1 \block_reg[7][123]  ( .D(block_next[123]), .E(n796), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFX1 \block_reg[7][122]  ( .D(block_next[122]), .E(n793), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFX1 \block_reg[7][95]  ( .D(block_next[95]), .E(n793), .CK(clk), .QN(n256) );
  EDFFX1 \block_reg[7][94]  ( .D(block_next[94]), .E(n796), .CK(clk), .QN(n272) );
  EDFFX1 \block_reg[7][93]  ( .D(block_next[93]), .E(n794), .CK(clk), .QN(n264) );
  EDFFX1 \block_reg[7][92]  ( .D(block_next[92]), .E(n795), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFX1 \block_reg[7][91]  ( .D(block_next[91]), .E(n798), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFX1 \block_reg[7][90]  ( .D(block_next[90]), .E(n798), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFX1 \block_reg[7][63]  ( .D(block_next[63]), .E(n796), .CK(clk), .QN(n248) );
  EDFFX1 \block_reg[7][62]  ( .D(block_next[62]), .E(n796), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFX1 \block_reg[7][61]  ( .D(block_next[61]), .E(n796), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFX1 \block_reg[7][60]  ( .D(block_next[60]), .E(n796), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFX1 \block_reg[7][59]  ( .D(block_next[59]), .E(n796), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFX1 \block_reg[7][58]  ( .D(block_next[58]), .E(n796), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFX1 \block_reg[7][31]  ( .D(block_next[31]), .E(n794), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFX1 \block_reg[7][30]  ( .D(block_next[30]), .E(n794), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFX1 \block_reg[7][29]  ( .D(block_next[29]), .E(n794), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFX1 \block_reg[7][28]  ( .D(block_next[28]), .E(n794), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFX1 \block_reg[7][27]  ( .D(block_next[27]), .E(n794), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFX1 \block_reg[7][26]  ( .D(block_next[26]), .E(n793), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFX1 \block_reg[3][127]  ( .D(block_next[127]), .E(n827), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFX1 \block_reg[3][126]  ( .D(block_next[126]), .E(n826), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFX1 \block_reg[3][125]  ( .D(block_next[125]), .E(n828), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFX1 \block_reg[3][124]  ( .D(block_next[124]), .E(n825), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFX1 \block_reg[3][123]  ( .D(block_next[123]), .E(n306), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFX1 \block_reg[3][122]  ( .D(block_next[122]), .E(n306), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFX1 \block_reg[3][95]  ( .D(block_next[95]), .E(n830), .CK(clk), .QN(n252) );
  EDFFX1 \block_reg[3][94]  ( .D(block_next[94]), .E(n823), .CK(clk), .QN(n268) );
  EDFFX1 \block_reg[3][93]  ( .D(block_next[93]), .E(n824), .CK(clk), .QN(n260) );
  EDFFX1 \block_reg[3][92]  ( .D(block_next[92]), .E(n306), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFX1 \block_reg[3][91]  ( .D(block_next[91]), .E(n830), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFX1 \block_reg[3][90]  ( .D(block_next[90]), .E(n830), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFX1 \block_reg[3][63]  ( .D(block_next[63]), .E(n828), .CK(clk), .QN(n244) );
  EDFFX1 \block_reg[3][62]  ( .D(block_next[62]), .E(n828), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFX1 \block_reg[3][61]  ( .D(block_next[61]), .E(n828), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFX1 \block_reg[3][60]  ( .D(block_next[60]), .E(n828), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFX1 \block_reg[3][59]  ( .D(block_next[59]), .E(n828), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFX1 \block_reg[3][58]  ( .D(block_next[58]), .E(n828), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFX1 \block_reg[3][31]  ( .D(block_next[31]), .E(n826), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFX1 \block_reg[3][30]  ( .D(block_next[30]), .E(n826), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFX1 \block_reg[3][29]  ( .D(block_next[29]), .E(n826), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFX1 \block_reg[3][28]  ( .D(block_next[28]), .E(n826), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFX1 \block_reg[3][27]  ( .D(block_next[27]), .E(n826), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFX1 \block_reg[3][26]  ( .D(block_next[26]), .E(n825), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFX1 \block_reg[5][127]  ( .D(block_next[127]), .E(n812), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFX1 \block_reg[5][126]  ( .D(block_next[126]), .E(n813), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFX1 \block_reg[5][125]  ( .D(block_next[125]), .E(n811), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFX1 \block_reg[5][124]  ( .D(block_next[124]), .E(n810), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFX1 \block_reg[5][123]  ( .D(block_next[123]), .E(n812), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFX1 \block_reg[5][122]  ( .D(block_next[122]), .E(n809), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFX1 \block_reg[5][95]  ( .D(block_next[95]), .E(n809), .CK(clk), .QN(n254) );
  EDFFX1 \block_reg[5][94]  ( .D(block_next[94]), .E(n812), .CK(clk), .QN(n270) );
  EDFFX1 \block_reg[5][93]  ( .D(block_next[93]), .E(n810), .CK(clk), .QN(n262) );
  EDFFX1 \block_reg[5][92]  ( .D(block_next[92]), .E(n811), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFX1 \block_reg[5][91]  ( .D(block_next[91]), .E(n814), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFX1 \block_reg[5][90]  ( .D(block_next[90]), .E(n814), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFX1 \block_reg[5][63]  ( .D(block_next[63]), .E(n812), .CK(clk), .QN(n246) );
  EDFFX1 \block_reg[5][62]  ( .D(block_next[62]), .E(n812), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFX1 \block_reg[5][61]  ( .D(block_next[61]), .E(n812), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFX1 \block_reg[5][60]  ( .D(block_next[60]), .E(n812), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFX1 \block_reg[5][59]  ( .D(block_next[59]), .E(n812), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFX1 \block_reg[5][58]  ( .D(block_next[58]), .E(n812), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFX1 \block_reg[5][31]  ( .D(block_next[31]), .E(n810), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFX1 \block_reg[5][30]  ( .D(block_next[30]), .E(n810), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFX1 \block_reg[5][29]  ( .D(block_next[29]), .E(n810), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFX1 \block_reg[5][28]  ( .D(block_next[28]), .E(n810), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFX1 \block_reg[5][27]  ( .D(block_next[27]), .E(n810), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFX1 \block_reg[5][26]  ( .D(block_next[26]), .E(n809), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFX1 \block_reg[1][127]  ( .D(block_next[127]), .E(n843), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFX1 \block_reg[1][126]  ( .D(block_next[126]), .E(n842), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFX1 \block_reg[1][125]  ( .D(block_next[125]), .E(n844), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFX1 \block_reg[1][124]  ( .D(block_next[124]), .E(n841), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFX1 \block_reg[1][123]  ( .D(block_next[123]), .E(n304), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFX1 \block_reg[1][122]  ( .D(block_next[122]), .E(n304), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFX1 \block_reg[1][95]  ( .D(block_next[95]), .E(n846), .CK(clk), .QN(n250) );
  EDFFX1 \block_reg[1][94]  ( .D(block_next[94]), .E(n839), .CK(clk), .QN(n266) );
  EDFFX1 \block_reg[1][93]  ( .D(block_next[93]), .E(n840), .CK(clk), .QN(n258) );
  EDFFX1 \block_reg[1][92]  ( .D(block_next[92]), .E(n304), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFX1 \block_reg[1][91]  ( .D(block_next[91]), .E(n846), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFX1 \block_reg[1][90]  ( .D(block_next[90]), .E(n846), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFX1 \block_reg[1][63]  ( .D(block_next[63]), .E(n844), .CK(clk), .QN(n242) );
  EDFFX1 \block_reg[1][62]  ( .D(block_next[62]), .E(n844), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFX1 \block_reg[1][61]  ( .D(block_next[61]), .E(n844), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFX1 \block_reg[1][60]  ( .D(block_next[60]), .E(n844), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFX1 \block_reg[1][59]  ( .D(block_next[59]), .E(n844), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFX1 \block_reg[1][58]  ( .D(block_next[58]), .E(n844), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFX1 \block_reg[1][31]  ( .D(block_next[31]), .E(n842), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFX1 \block_reg[1][30]  ( .D(block_next[30]), .E(n842), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFX1 \block_reg[1][29]  ( .D(block_next[29]), .E(n842), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFX1 \block_reg[1][28]  ( .D(block_next[28]), .E(n842), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFX1 \block_reg[1][27]  ( .D(block_next[27]), .E(n842), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFX1 \block_reg[1][26]  ( .D(block_next[26]), .E(n841), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFX1 \block_reg[4][127]  ( .D(block_next[127]), .E(n821), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFX1 \block_reg[4][126]  ( .D(block_next[126]), .E(n816), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFX1 \block_reg[4][125]  ( .D(block_next[125]), .E(n815), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFX1 \block_reg[4][124]  ( .D(block_next[124]), .E(n817), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFX1 \block_reg[4][123]  ( .D(block_next[123]), .E(n822), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFX1 \block_reg[4][122]  ( .D(block_next[122]), .E(n817), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFX1 \block_reg[4][95]  ( .D(block_next[95]), .E(n822), .CK(clk), .QN(n253) );
  EDFFX1 \block_reg[4][94]  ( .D(block_next[94]), .E(n822), .CK(clk), .QN(n269) );
  EDFFX1 \block_reg[4][93]  ( .D(block_next[93]), .E(n822), .CK(clk), .QN(n261) );
  EDFFX1 \block_reg[4][92]  ( .D(block_next[92]), .E(n822), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFX1 \block_reg[4][91]  ( .D(block_next[91]), .E(n821), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFX1 \block_reg[4][90]  ( .D(block_next[90]), .E(n821), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFX1 \block_reg[4][63]  ( .D(block_next[63]), .E(n820), .CK(clk), .QN(n245) );
  EDFFX1 \block_reg[4][62]  ( .D(block_next[62]), .E(n820), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFX1 \block_reg[4][61]  ( .D(block_next[61]), .E(n820), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFX1 \block_reg[4][60]  ( .D(block_next[60]), .E(n820), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFX1 \block_reg[4][59]  ( .D(block_next[59]), .E(n820), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFX1 \block_reg[4][58]  ( .D(block_next[58]), .E(n820), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFX1 \block_reg[4][31]  ( .D(block_next[31]), .E(n818), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFX1 \block_reg[4][30]  ( .D(block_next[30]), .E(n818), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFX1 \block_reg[4][29]  ( .D(block_next[29]), .E(n818), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFX1 \block_reg[4][28]  ( .D(block_next[28]), .E(n818), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFX1 \block_reg[4][27]  ( .D(block_next[27]), .E(n818), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFX1 \block_reg[4][26]  ( .D(block_next[26]), .E(n822), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFX1 \block_reg[0][127]  ( .D(block_next[127]), .E(n848), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFX1 \block_reg[0][126]  ( .D(block_next[126]), .E(n847), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFX1 \block_reg[0][125]  ( .D(block_next[125]), .E(n849), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFX1 \block_reg[0][124]  ( .D(block_next[124]), .E(n850), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFX1 \block_reg[0][123]  ( .D(block_next[123]), .E(n852), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFX1 \block_reg[0][122]  ( .D(block_next[122]), .E(n851), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFX1 \block_reg[0][95]  ( .D(block_next[95]), .E(n851), .CK(clk), .QN(n249) );
  EDFFX1 \block_reg[0][94]  ( .D(block_next[94]), .E(n852), .CK(clk), .QN(n265) );
  EDFFX1 \block_reg[0][93]  ( .D(block_next[93]), .E(n850), .CK(clk), .QN(n257) );
  EDFFX1 \block_reg[0][92]  ( .D(block_next[92]), .E(n849), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFX1 \block_reg[0][91]  ( .D(block_next[91]), .E(n854), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFX1 \block_reg[0][90]  ( .D(block_next[90]), .E(n854), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFX1 \block_reg[0][63]  ( .D(block_next[63]), .E(n852), .CK(clk), .QN(n241) );
  EDFFX1 \block_reg[0][62]  ( .D(block_next[62]), .E(n852), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFX1 \block_reg[0][61]  ( .D(block_next[61]), .E(n852), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFX1 \block_reg[0][60]  ( .D(block_next[60]), .E(n852), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFX1 \block_reg[0][59]  ( .D(block_next[59]), .E(n852), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFX1 \block_reg[0][58]  ( .D(block_next[58]), .E(n852), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFX1 \block_reg[0][31]  ( .D(block_next[31]), .E(n850), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFX1 \block_reg[0][30]  ( .D(block_next[30]), .E(n850), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFX1 \block_reg[0][29]  ( .D(block_next[29]), .E(n850), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFX1 \block_reg[0][28]  ( .D(block_next[28]), .E(n850), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFX1 \block_reg[0][27]  ( .D(block_next[27]), .E(n850), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFX1 \block_reg[0][26]  ( .D(block_next[26]), .E(n851), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFX1 \block_reg[6][127]  ( .D(block_next[127]), .E(n805), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFX1 \block_reg[6][126]  ( .D(block_next[126]), .E(n800), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFX1 \block_reg[6][125]  ( .D(block_next[125]), .E(n799), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFX1 \block_reg[6][124]  ( .D(block_next[124]), .E(n801), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFX1 \block_reg[6][123]  ( .D(block_next[123]), .E(n806), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFX1 \block_reg[6][122]  ( .D(block_next[122]), .E(n801), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFX1 \block_reg[6][95]  ( .D(block_next[95]), .E(n806), .CK(clk), .QN(n255) );
  EDFFX1 \block_reg[6][94]  ( .D(block_next[94]), .E(n806), .CK(clk), .QN(n271) );
  EDFFX1 \block_reg[6][93]  ( .D(block_next[93]), .E(n806), .CK(clk), .QN(n263) );
  EDFFX1 \block_reg[6][92]  ( .D(block_next[92]), .E(n806), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFX1 \block_reg[6][91]  ( .D(block_next[91]), .E(n805), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFX1 \block_reg[6][90]  ( .D(block_next[90]), .E(n805), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFX1 \block_reg[6][63]  ( .D(block_next[63]), .E(n804), .CK(clk), .QN(n247) );
  EDFFX1 \block_reg[6][62]  ( .D(block_next[62]), .E(n804), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFX1 \block_reg[6][61]  ( .D(block_next[61]), .E(n804), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFX1 \block_reg[6][60]  ( .D(block_next[60]), .E(n804), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFX1 \block_reg[6][59]  ( .D(block_next[59]), .E(n804), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFX1 \block_reg[6][58]  ( .D(block_next[58]), .E(n804), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFX1 \block_reg[6][31]  ( .D(block_next[31]), .E(n802), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFX1 \block_reg[6][30]  ( .D(block_next[30]), .E(n802), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFX1 \block_reg[6][29]  ( .D(block_next[29]), .E(n802), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFX1 \block_reg[6][28]  ( .D(block_next[28]), .E(n802), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFX1 \block_reg[6][27]  ( .D(block_next[27]), .E(n802), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFX1 \block_reg[6][26]  ( .D(block_next[26]), .E(n806), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFX1 \block_reg[2][127]  ( .D(block_next[127]), .E(n832), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFX1 \block_reg[2][126]  ( .D(block_next[126]), .E(n831), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFX1 \block_reg[2][125]  ( .D(block_next[125]), .E(n833), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFX1 \block_reg[2][124]  ( .D(block_next[124]), .E(n834), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFX1 \block_reg[2][123]  ( .D(block_next[123]), .E(n836), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFX1 \block_reg[2][122]  ( .D(block_next[122]), .E(n835), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFX1 \block_reg[2][95]  ( .D(block_next[95]), .E(n835), .CK(clk), .QN(n251) );
  EDFFX1 \block_reg[2][94]  ( .D(block_next[94]), .E(n836), .CK(clk), .QN(n267) );
  EDFFX1 \block_reg[2][93]  ( .D(block_next[93]), .E(n834), .CK(clk), .QN(n259) );
  EDFFX1 \block_reg[2][92]  ( .D(block_next[92]), .E(n833), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFX1 \block_reg[2][91]  ( .D(block_next[91]), .E(n838), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFX1 \block_reg[2][90]  ( .D(block_next[90]), .E(n838), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFX1 \block_reg[2][63]  ( .D(block_next[63]), .E(n836), .CK(clk), .QN(n243) );
  EDFFX1 \block_reg[2][62]  ( .D(block_next[62]), .E(n836), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFX1 \block_reg[2][61]  ( .D(block_next[61]), .E(n836), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFX1 \block_reg[2][60]  ( .D(block_next[60]), .E(n836), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFX1 \block_reg[2][59]  ( .D(block_next[59]), .E(n836), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFX1 \block_reg[2][58]  ( .D(block_next[58]), .E(n836), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFX1 \block_reg[2][31]  ( .D(block_next[31]), .E(n834), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFX1 \block_reg[2][30]  ( .D(block_next[30]), .E(n834), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFX1 \block_reg[2][29]  ( .D(block_next[29]), .E(n834), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFX1 \block_reg[2][28]  ( .D(block_next[28]), .E(n834), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFX1 \block_reg[2][27]  ( .D(block_next[27]), .E(n834), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFX1 \block_reg[2][26]  ( .D(block_next[26]), .E(n835), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(n78), .E(n816), .CK(clk), .Q(
        \blocktag[4][22] ) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(n11), .E(n816), .CK(clk), .Q(
        \blocktag[4][21] ) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(n10), .E(n816), .CK(clk), .Q(
        \blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(n77), .E(n816), .CK(clk), .Q(
        \blocktag[4][19] ) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(n816), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(n9), .E(n816), .CK(clk), .QN(n343) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n815), .CK(clk), .QN(
        n232) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(n78), .E(n848), .CK(clk), .Q(
        \blocktag[0][22] ) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(n11), .E(n848), .CK(clk), .Q(
        \blocktag[0][21] ) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(n10), .E(n848), .CK(clk), .Q(
        \blocktag[0][20] ) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(n77), .E(n848), .CK(clk), .Q(
        \blocktag[0][19] ) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(n848), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(n76), .E(n848), .CK(clk), .Q(
        \blocktag[0][14] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(n9), .E(n848), .CK(clk), .QN(n339) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n847), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(n78), .E(n307), .CK(clk), .Q(
        \blocktag[7][22] ) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(n11), .E(n307), .CK(clk), .Q(
        \blocktag[7][21] ) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(n10), .E(n791), .CK(clk), .Q(
        \blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(n77), .E(n792), .CK(clk), .Q(
        \blocktag[7][19] ) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(n792), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(n9), .E(n793), .CK(clk), .QN(n346) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n791), .CK(clk), .QN(
        n235) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(n78), .E(n824), .CK(clk), .Q(
        \blocktag[3][22] ) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(n11), .E(n824), .CK(clk), .Q(
        \blocktag[3][21] ) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(n10), .E(n824), .CK(clk), .Q(
        \blocktag[3][20] ) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(n77), .E(n824), .CK(clk), .Q(
        \blocktag[3][19] ) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(n824), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(n76), .E(n824), .CK(clk), .Q(
        \blocktag[3][14] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(n9), .E(n824), .CK(clk), .QN(n342) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n823), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(n78), .E(n305), .CK(clk), .Q(
        \blocktag[5][22] ) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(n11), .E(n305), .CK(clk), .Q(
        \blocktag[5][21] ) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(n10), .E(n807), .CK(clk), .Q(
        \blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(n77), .E(n808), .CK(clk), .Q(
        \blocktag[5][19] ) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(n808), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(n9), .E(n809), .CK(clk), .QN(n344) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(n807), .CK(clk), .QN(
        n233) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(n78), .E(n840), .CK(clk), .Q(
        \blocktag[1][22] ) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(n11), .E(n840), .CK(clk), .Q(
        \blocktag[1][21] ) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(n10), .E(n840), .CK(clk), .Q(
        \blocktag[1][20] ) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(n77), .E(n840), .CK(clk), .Q(
        \blocktag[1][19] ) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n840), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(n76), .E(n840), .CK(clk), .Q(
        \blocktag[1][14] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(n9), .E(n840), .CK(clk), .QN(n340) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n839), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(n78), .E(n800), .CK(clk), .Q(
        \blocktag[6][22] ) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(n11), .E(n800), .CK(clk), .Q(
        \blocktag[6][21] ) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(n10), .E(n800), .CK(clk), .Q(
        \blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(n77), .E(n800), .CK(clk), .Q(
        \blocktag[6][19] ) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n800), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(n9), .E(n800), .CK(clk), .QN(n345) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n799), .CK(clk), .QN(
        n234) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(n78), .E(n832), .CK(clk), .Q(
        \blocktag[2][22] ) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(n11), .E(n832), .CK(clk), .Q(
        \blocktag[2][21] ) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(n10), .E(n832), .CK(clk), .Q(
        \blocktag[2][20] ) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(n77), .E(n832), .CK(clk), .Q(
        \blocktag[2][19] ) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(n832), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(n76), .E(n832), .CK(clk), .Q(
        \blocktag[2][14] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(n9), .E(n832), .CK(clk), .QN(n341) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n831), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(n75), .E(n798), .CK(clk), .Q(
        \blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(n74), .E(n793), .CK(clk), .Q(
        \blocktag[7][23] ) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(n375), .E(n797), .CK(clk), .Q(
        \blocktag[7][18] ) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(n73), .E(n795), .CK(clk), .Q(
        \blocktag[7][16] ) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(n76), .E(n794), .CK(clk), .Q(
        \blocktag[7][14] ) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(n71), .E(n791), .CK(clk), .Q(
        \blocktag[7][12] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(n70), .E(n791), .CK(clk), .Q(
        \blocktag[7][11] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(n69), .E(n791), .CK(clk), .Q(
        \blocktag[7][10] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(n68), .E(n791), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(n67), .E(n791), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(n66), .E(n791), .CK(clk), .Q(
        \blocktag[7][7] ) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(n65), .E(n791), .CK(clk), .Q(
        \blocktag[7][6] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(n374), .E(n791), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(n64), .E(n791), .CK(clk), .Q(
        \blocktag[7][4] ) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(n373), .E(n791), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(n372), .E(n791), .CK(clk), .QN(n191) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(n63), .E(n791), .CK(clk), .Q(
        \blocktag[7][1] ) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(n75), .E(n824), .CK(clk), .Q(
        \blocktag[3][24] ) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(n74), .E(n824), .CK(clk), .Q(
        \blocktag[3][23] ) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(n375), .E(n824), .CK(clk), .Q(
        \blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(n72), .E(n824), .CK(clk), .Q(
        \blocktag[3][17] ) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(n73), .E(n824), .CK(clk), .Q(
        \blocktag[3][16] ) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(n71), .E(n823), .CK(clk), .Q(
        \blocktag[3][12] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(n70), .E(n823), .CK(clk), .Q(
        \blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(n69), .E(n823), .CK(clk), .Q(
        \blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[3][9]  ( .D(n68), .E(n823), .CK(clk), .Q(
        \blocktag[3][9] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(n67), .E(n823), .CK(clk), .Q(
        \blocktag[3][8] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(n66), .E(n823), .CK(clk), .Q(
        \blocktag[3][7] ) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(n65), .E(n823), .CK(clk), .Q(
        \blocktag[3][6] ) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(n374), .E(n823), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(n64), .E(n823), .CK(clk), .Q(
        \blocktag[3][4] ) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(n373), .E(n823), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(n372), .E(n823), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(n63), .E(n823), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(n75), .E(n814), .CK(clk), .Q(
        \blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(n74), .E(n809), .CK(clk), .Q(
        \blocktag[5][23] ) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(n375), .E(n813), .CK(clk), .Q(
        \blocktag[5][18] ) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(n73), .E(n811), .CK(clk), .Q(
        \blocktag[5][16] ) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(n76), .E(n810), .CK(clk), .Q(
        \blocktag[5][14] ) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(n71), .E(n807), .CK(clk), .Q(
        \blocktag[5][12] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(n70), .E(n807), .CK(clk), .Q(
        \blocktag[5][11] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(n69), .E(n807), .CK(clk), .Q(
        \blocktag[5][10] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(n68), .E(n807), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(n67), .E(n807), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(n66), .E(n807), .CK(clk), .Q(
        \blocktag[5][7] ) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(n65), .E(n807), .CK(clk), .Q(
        \blocktag[5][6] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(n374), .E(n807), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(n64), .E(n807), .CK(clk), .Q(
        \blocktag[5][4] ) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(n373), .E(n807), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(n372), .E(n807), .CK(clk), .QN(n189) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(n63), .E(n807), .CK(clk), .Q(
        \blocktag[5][1] ) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(n75), .E(n840), .CK(clk), .Q(
        \blocktag[1][24] ) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(n74), .E(n840), .CK(clk), .Q(
        \blocktag[1][23] ) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(n375), .E(n840), .CK(clk), .Q(
        \blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(n72), .E(n840), .CK(clk), .Q(
        \blocktag[1][17] ) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(n73), .E(n840), .CK(clk), .Q(
        \blocktag[1][16] ) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(n71), .E(n839), .CK(clk), .Q(
        \blocktag[1][12] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(n70), .E(n839), .CK(clk), .Q(
        \blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(n69), .E(n839), .CK(clk), .Q(
        \blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[1][9]  ( .D(n68), .E(n839), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(n67), .E(n839), .CK(clk), .Q(
        \blocktag[1][8] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(n66), .E(n839), .CK(clk), .Q(
        \blocktag[1][7] ) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(n65), .E(n839), .CK(clk), .Q(
        \blocktag[1][6] ) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(n374), .E(n839), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(n64), .E(n839), .CK(clk), .Q(
        \blocktag[1][4] ) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(n373), .E(n839), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(n372), .E(n839), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(n63), .E(n839), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(n75), .E(n816), .CK(clk), .Q(
        \blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(n74), .E(n816), .CK(clk), .Q(
        \blocktag[4][23] ) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(n375), .E(n816), .CK(clk), .Q(
        \blocktag[4][18] ) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(n73), .E(n816), .CK(clk), .Q(
        \blocktag[4][16] ) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(n76), .E(n816), .CK(clk), .Q(
        \blocktag[4][14] ) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(n71), .E(n815), .CK(clk), .Q(
        \blocktag[4][12] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(n70), .E(n815), .CK(clk), .Q(
        \blocktag[4][11] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(n69), .E(n815), .CK(clk), .Q(
        \blocktag[4][10] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(n68), .E(n815), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(n67), .E(n815), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(n66), .E(n815), .CK(clk), .Q(
        \blocktag[4][7] ) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(n65), .E(n815), .CK(clk), .Q(
        \blocktag[4][6] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(n374), .E(n815), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(n64), .E(n815), .CK(clk), .Q(
        \blocktag[4][4] ) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(n373), .E(n815), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(n372), .E(n815), .CK(clk), .QN(n188) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(n63), .E(n815), .CK(clk), .Q(
        \blocktag[4][1] ) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(n75), .E(n848), .CK(clk), .Q(
        \blocktag[0][24] ) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(n74), .E(n848), .CK(clk), .Q(
        \blocktag[0][23] ) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(n375), .E(n848), .CK(clk), .Q(
        \blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(n72), .E(n848), .CK(clk), .Q(
        \blocktag[0][17] ) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(n73), .E(n848), .CK(clk), .Q(
        \blocktag[0][16] ) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(n71), .E(n847), .CK(clk), .Q(
        \blocktag[0][12] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(n70), .E(n847), .CK(clk), .Q(
        \blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(n69), .E(n847), .CK(clk), .Q(
        \blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[0][9]  ( .D(n68), .E(n847), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(n67), .E(n847), .CK(clk), .Q(
        \blocktag[0][8] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(n66), .E(n847), .CK(clk), .Q(
        \blocktag[0][7] ) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(n65), .E(n847), .CK(clk), .Q(
        \blocktag[0][6] ) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(n374), .E(n847), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(n64), .E(n847), .CK(clk), .Q(
        \blocktag[0][4] ) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(n373), .E(n847), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(n372), .E(n847), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(n63), .E(n847), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(n75), .E(n800), .CK(clk), .Q(
        \blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(n74), .E(n800), .CK(clk), .Q(
        \blocktag[6][23] ) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(n375), .E(n800), .CK(clk), .Q(
        \blocktag[6][18] ) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(n73), .E(n800), .CK(clk), .Q(
        \blocktag[6][16] ) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(n76), .E(n800), .CK(clk), .Q(
        \blocktag[6][14] ) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(n71), .E(n799), .CK(clk), .Q(
        \blocktag[6][12] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(n70), .E(n799), .CK(clk), .Q(
        \blocktag[6][11] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(n69), .E(n799), .CK(clk), .Q(
        \blocktag[6][10] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(n68), .E(n799), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(n67), .E(n799), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(n66), .E(n799), .CK(clk), .Q(
        \blocktag[6][7] ) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(n65), .E(n799), .CK(clk), .Q(
        \blocktag[6][6] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(n374), .E(n799), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(n64), .E(n799), .CK(clk), .Q(
        \blocktag[6][4] ) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(n373), .E(n799), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(n372), .E(n799), .CK(clk), .QN(n190) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(n63), .E(n799), .CK(clk), .Q(
        \blocktag[6][1] ) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(n75), .E(n832), .CK(clk), .Q(
        \blocktag[2][24] ) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(n74), .E(n832), .CK(clk), .Q(
        \blocktag[2][23] ) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(n375), .E(n832), .CK(clk), .Q(
        \blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(n72), .E(n832), .CK(clk), .Q(
        \blocktag[2][17] ) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(n73), .E(n832), .CK(clk), .Q(
        \blocktag[2][16] ) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(n71), .E(n831), .CK(clk), .Q(
        \blocktag[2][12] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(n70), .E(n831), .CK(clk), .Q(
        \blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(n69), .E(n831), .CK(clk), .Q(
        \blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[2][9]  ( .D(n68), .E(n831), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(n67), .E(n831), .CK(clk), .Q(
        \blocktag[2][8] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(n66), .E(n831), .CK(clk), .Q(
        \blocktag[2][7] ) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(n65), .E(n831), .CK(clk), .Q(
        \blocktag[2][6] ) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(n374), .E(n831), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(n64), .E(n831), .CK(clk), .Q(
        \blocktag[2][4] ) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(n373), .E(n831), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(n372), .E(n831), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(n63), .E(n831), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(n72), .E(n812), .CK(clk), .Q(
        \blocktag[5][17] ) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(n72), .E(n800), .CK(clk), .Q(
        \blocktag[6][17] ) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(n72), .E(n796), .CK(clk), .Q(
        \blocktag[7][17] ) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(n72), .E(n816), .CK(clk), .Q(
        \blocktag[4][17] ) );
  DFFRX1 \blockvalid_reg[7]  ( .D(n1278), .CK(clk), .RN(n865), .Q(
        blockvalid[7]), .QN(n1294) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n1280), .CK(clk), .RN(n865), .Q(
        blockvalid[5]), .QN(n1296) );
  DFFRX1 \blockvalid_reg[3]  ( .D(n1282), .CK(clk), .RN(n865), .Q(
        blockvalid[3]), .QN(n1298) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n1284), .CK(clk), .RN(n865), .Q(
        blockvalid[1]), .QN(n1300) );
  DFFRX1 \blockvalid_reg[6]  ( .D(n1279), .CK(clk), .RN(n865), .Q(
        blockvalid[6]), .QN(n1295) );
  DFFRX1 \blockvalid_reg[4]  ( .D(n1281), .CK(clk), .RN(n865), .Q(
        blockvalid[4]), .QN(n1297) );
  DFFRX1 \blockvalid_reg[2]  ( .D(n1283), .CK(clk), .RN(n865), .Q(
        blockvalid[2]), .QN(n1299) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n1285), .CK(clk), .RN(n865), .Q(
        blockvalid[0]), .QN(n1301) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n1286), .CK(clk), .RN(n865), .Q(
        blockdirty[7]), .QN(n1302) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n1288), .CK(clk), .RN(n865), .Q(
        blockdirty[5]), .QN(n1304) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n1290), .CK(clk), .RN(n865), .Q(
        blockdirty[3]), .QN(n1306) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n1292), .CK(clk), .RN(n865), .Q(
        blockdirty[1]), .QN(n1308) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n1287), .CK(clk), .RN(n865), .Q(
        blockdirty[6]), .QN(n1303) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n1289), .CK(clk), .RN(n865), .Q(
        blockdirty[4]), .QN(n1305) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n1291), .CK(clk), .RN(n865), .Q(
        blockdirty[2]), .QN(n1307) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n1293), .CK(clk), .RN(n865), .Q(
        blockdirty[0]), .QN(n1309) );
  CLKINVX4 U3 ( .A(n1113), .Y(n1110) );
  MX4X2 U4 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n199), .S1(n729), .Y(
        n332) );
  AND3X6 U5 ( .A(n888), .B(n887), .C(n886), .Y(n889) );
  BUFX16 U6 ( .A(n1270), .Y(n1) );
  NOR2X6 U7 ( .A(n1), .B(n1269), .Y(n196) );
  BUFX20 U8 ( .A(n1277), .Y(n2) );
  BUFX6 U9 ( .A(n1), .Y(n4) );
  CLKBUFX3 U10 ( .A(n4), .Y(n7) );
  CLKBUFX3 U11 ( .A(n4), .Y(n8) );
  CLKBUFX3 U12 ( .A(n8), .Y(n784) );
  BUFX20 U13 ( .A(n1272), .Y(n3) );
  NOR2X4 U14 ( .A(n3), .B(n1271), .Y(n195) );
  OA22X2 U15 ( .A0(n3), .A1(n1250), .B0(n1), .B1(n1249), .Y(n1251) );
  OA22X4 U16 ( .A0(n3), .A1(n1245), .B0(n4), .B1(n1244), .Y(n1246) );
  OA22X4 U17 ( .A0(n3), .A1(n1255), .B0(n4), .B1(n1254), .Y(n1256) );
  NAND2X6 U18 ( .A(n376), .B(n1110), .Y(n1275) );
  CLKBUFX2 U19 ( .A(n784), .Y(n785) );
  CLKBUFX3 U20 ( .A(n2), .Y(n5) );
  CLKBUFX2 U21 ( .A(n2), .Y(n6) );
  NAND2X6 U22 ( .A(n228), .B(n229), .Y(n239) );
  NAND2X6 U23 ( .A(n223), .B(proc_addr[5]), .Y(n228) );
  XOR2X4 U24 ( .A(n1074), .B(proc_addr[24]), .Y(n884) );
  XOR2X4 U25 ( .A(proc_addr[10]), .B(tag[5]), .Y(n876) );
  CLKMX2X12 U26 ( .A(n367), .B(n368), .S0(n698), .Y(tag[5]) );
  MX4X2 U27 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n199), .S1(n727), .Y(
        n327) );
  MX4XL U28 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n731), .S1(n727), .Y(
        n328) );
  MX4X2 U29 ( .A(\blocktag[0][23] ), .B(\blocktag[1][23] ), .C(
        \blocktag[2][23] ), .D(\blocktag[3][23] ), .S0(n198), .S1(n727), .Y(
        n357) );
  MX4X2 U30 ( .A(\blocktag[4][23] ), .B(\blocktag[5][23] ), .C(
        \blocktag[6][23] ), .D(\blocktag[7][23] ), .S0(n198), .S1(n727), .Y(
        n358) );
  CLKBUFX20 U31 ( .A(n702), .Y(n727) );
  XOR2X2 U32 ( .A(n1089), .B(proc_addr[14]), .Y(n879) );
  NAND4X2 U33 ( .A(n873), .B(n872), .C(n871), .D(n870), .Y(n892) );
  NAND4X2 U34 ( .A(n881), .B(n880), .C(n879), .D(n878), .Y(n891) );
  NOR4X4 U35 ( .A(n877), .B(n876), .C(n875), .D(n874), .Y(n878) );
  INVX20 U36 ( .A(n197), .Y(n200) );
  CLKINVX20 U37 ( .A(n753), .Y(n197) );
  AND4X8 U38 ( .A(n885), .B(n884), .C(n883), .D(n882), .Y(n230) );
  XNOR2X2 U39 ( .A(n1070), .B(proc_addr[28]), .Y(n240) );
  MX4X2 U40 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n198), .S1(n726), .Y(
        n331) );
  INVX12 U41 ( .A(n197), .Y(n198) );
  XNOR2X4 U42 ( .A(n1068), .B(proc_addr[29]), .Y(n238) );
  MX4X2 U43 ( .A(\blocktag[4][17] ), .B(\blocktag[6][17] ), .C(
        \blocktag[5][17] ), .D(\blocktag[7][17] ), .S0(n726), .S1(n200), .Y(
        n338) );
  MX4X2 U44 ( .A(\blocktag[0][12] ), .B(\blocktag[1][12] ), .C(
        \blocktag[2][12] ), .D(\blocktag[3][12] ), .S0(n755), .S1(n726), .Y(
        n333) );
  MX4X2 U45 ( .A(\blocktag[4][12] ), .B(\blocktag[5][12] ), .C(
        \blocktag[6][12] ), .D(\blocktag[7][12] ), .S0(n731), .S1(n726), .Y(
        n334) );
  BUFX20 U46 ( .A(n728), .Y(n726) );
  NOR2X2 U47 ( .A(n195), .B(n196), .Y(n1273) );
  OA22X4 U48 ( .A0(n3), .A1(n1265), .B0(n1), .B1(n1264), .Y(n1266) );
  XOR2X2 U49 ( .A(n1081), .B(proc_addr[19]), .Y(n867) );
  AND3X6 U50 ( .A(n869), .B(n868), .C(n867), .Y(n870) );
  CLKXOR2X2 U51 ( .A(n1078), .B(proc_addr[21]), .Y(n869) );
  XOR2X4 U52 ( .A(n1076), .B(proc_addr[22]), .Y(n887) );
  CLKINVX6 U53 ( .A(tag[17]), .Y(n1076) );
  NOR3X4 U54 ( .A(n238), .B(n239), .C(n240), .Y(n882) );
  XOR2X4 U55 ( .A(n1083), .B(proc_addr[17]), .Y(n868) );
  INVX6 U56 ( .A(tag[12]), .Y(n1083) );
  OAI221X2 U57 ( .A0(n2), .A1(n1263), .B0(n1275), .B1(n1262), .C0(n1261), .Y(
        proc_rdata[29]) );
  INVX8 U58 ( .A(tag[22]), .Y(n1072) );
  MXI2X4 U59 ( .A(n672), .B(n673), .S0(n697), .Y(tag[22]) );
  NAND4BBX4 U60 ( .AN(n892), .BN(n891), .C(n230), .D(n231), .Y(n1104) );
  AND3X8 U61 ( .A(n889), .B(n890), .C(n371), .Y(n231) );
  CLKINVX1 U62 ( .A(blockdata[107]), .Y(n1172) );
  OA22X2 U63 ( .A0(n789), .A1(n1190), .B0(n784), .B1(n1189), .Y(n1191) );
  XOR2X1 U64 ( .A(proc_addr[8]), .B(tag[3]), .Y(n875) );
  XNOR2X1 U65 ( .A(n192), .B(tag[2]), .Y(n877) );
  CLKINVX1 U66 ( .A(proc_addr[7]), .Y(n192) );
  XOR2X1 U67 ( .A(n1095), .B(proc_addr[11]), .Y(n881) );
  AND2X2 U68 ( .A(n236), .B(n237), .Y(n371) );
  XOR2X1 U69 ( .A(n1099), .B(proc_addr[6]), .Y(n236) );
  XOR2X1 U70 ( .A(n15), .B(proc_addr[20]), .Y(n237) );
  XOR2X1 U71 ( .A(n1072), .B(proc_addr[27]), .Y(n886) );
  XOR2X1 U72 ( .A(n1087), .B(proc_addr[15]), .Y(n888) );
  XOR2X1 U73 ( .A(n12), .B(proc_addr[18]), .Y(n890) );
  XOR2X1 U74 ( .A(n1091), .B(proc_addr[13]), .Y(n872) );
  XOR2X1 U75 ( .A(n1085), .B(proc_addr[16]), .Y(n871) );
  XOR2X1 U76 ( .A(n1093), .B(proc_addr[12]), .Y(n873) );
  XOR2X1 U77 ( .A(n13), .B(proc_addr[25]), .Y(n885) );
  XOR2X1 U78 ( .A(n1097), .B(proc_addr[9]), .Y(n880) );
  CLKBUFX3 U79 ( .A(proc_read), .Y(n863) );
  CLKINVX6 U80 ( .A(n1104), .Y(n893) );
  MXI2X1 U81 ( .A(n670), .B(n671), .S0(n689), .Y(dirty) );
  CLKMX2X2 U82 ( .A(n325), .B(n326), .S0(n696), .Y(valid) );
  MX4X1 U83 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n752), .S1(n705), .Y(n326) );
  NAND2X1 U84 ( .A(n866), .B(n1108), .Y(n1103) );
  MX4X1 U85 ( .A(n232), .B(n233), .C(n234), .D(n235), .S0(n754), .S1(n728), 
        .Y(n685) );
  MXI4X2 U86 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(\blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n754), .S1(n728), .Y(n684) );
  CLKINVX1 U87 ( .A(n1064), .Y(proc_stall) );
  MXI2X1 U88 ( .A(n612), .B(n613), .S0(n696), .Y(blockdata[28]) );
  MXI2X1 U89 ( .A(n548), .B(n549), .S0(n693), .Y(blockdata[60]) );
  MXI2X1 U90 ( .A(n448), .B(n449), .S0(n691), .Y(blockdata[92]) );
  MXI2X1 U91 ( .A(n384), .B(n385), .S0(n690), .Y(blockdata[124]) );
  CLKMX2X2 U92 ( .A(n355), .B(n356), .S0(n698), .Y(tag[1]) );
  MX4X1 U93 ( .A(\blocktag[4][1] ), .B(\blocktag[5][1] ), .C(\blocktag[6][1] ), 
        .D(\blocktag[7][1] ), .S0(n754), .S1(n728), .Y(n356) );
  CLKMX2X2 U94 ( .A(n361), .B(n362), .S0(n698), .Y(tag[4]) );
  CLKMX2X2 U95 ( .A(n363), .B(n364), .S0(n698), .Y(tag[6]) );
  MX4X1 U96 ( .A(\blocktag[0][6] ), .B(\blocktag[1][6] ), .C(\blocktag[2][6] ), 
        .D(\blocktag[3][6] ), .S0(n754), .S1(n727), .Y(n363) );
  CLKMX2X2 U97 ( .A(n353), .B(n354), .S0(n698), .Y(tag[7]) );
  CLKMX2X2 U98 ( .A(n351), .B(n352), .S0(n698), .Y(tag[8]) );
  CLKMX2X2 U99 ( .A(n359), .B(n360), .S0(n698), .Y(tag[9]) );
  CLKMX2X2 U100 ( .A(n327), .B(n328), .S0(n698), .Y(tag[10]) );
  CLKMX2X2 U101 ( .A(n349), .B(n350), .S0(n698), .Y(tag[11]) );
  CLKMX2X2 U102 ( .A(n333), .B(n334), .S0(n686), .Y(tag[12]) );
  CLKMX2X2 U103 ( .A(n331), .B(n332), .S0(n686), .Y(tag[14]) );
  CLKMX2X2 U104 ( .A(n335), .B(n336), .S0(n686), .Y(tag[16]) );
  MX4X1 U105 ( .A(\blocktag[4][16] ), .B(\blocktag[5][16] ), .C(
        \blocktag[6][16] ), .D(\blocktag[7][16] ), .S0(n200), .S1(n726), .Y(
        n336) );
  MX4X1 U106 ( .A(\blocktag[0][16] ), .B(\blocktag[1][16] ), .C(
        \blocktag[2][16] ), .D(\blocktag[3][16] ), .S0(n200), .S1(n726), .Y(
        n335) );
  CLKMX2X2 U107 ( .A(n337), .B(n338), .S0(n686), .Y(tag[17]) );
  MX4X1 U108 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n199), .S1(n726), .Y(
        n337) );
  CLKMX2X2 U109 ( .A(n347), .B(n348), .S0(n697), .Y(tag[19]) );
  MXI4X1 U110 ( .A(\blocktag[0][22] ), .B(\blocktag[1][22] ), .C(
        \blocktag[2][22] ), .D(\blocktag[3][22] ), .S0(n199), .S1(n730), .Y(
        n672) );
  MXI4X1 U111 ( .A(\blocktag[4][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[7][22] ), .S0(n199), .S1(n727), .Y(
        n673) );
  CLKMX2X2 U112 ( .A(n357), .B(n358), .S0(n686), .Y(tag[23]) );
  CLKMX2X2 U113 ( .A(n329), .B(n330), .S0(n698), .Y(tag[24]) );
  MX4X1 U114 ( .A(\blocktag[0][24] ), .B(\blocktag[1][24] ), .C(
        \blocktag[2][24] ), .D(\blocktag[3][24] ), .S0(n199), .S1(n730), .Y(
        n329) );
  MX4X1 U115 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n200), .S1(n730), .Y(
        n330) );
  INVX3 U116 ( .A(tag[1]), .Y(n1099) );
  CLKINVX1 U117 ( .A(tag[4]), .Y(n1097) );
  MX4X1 U118 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(\blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n754), .S1(n728), .Y(n367) );
  MX4X1 U119 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(\blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n754), .S1(n728), .Y(n368) );
  INVX6 U120 ( .A(tag[6]), .Y(n1095) );
  INVX3 U121 ( .A(tag[7]), .Y(n1093) );
  INVX3 U122 ( .A(tag[8]), .Y(n1091) );
  INVX3 U123 ( .A(tag[9]), .Y(n1089) );
  INVX3 U124 ( .A(tag[10]), .Y(n1087) );
  INVX3 U125 ( .A(tag[11]), .Y(n1085) );
  INVX3 U126 ( .A(tag[16]), .Y(n1078) );
  MX2X6 U127 ( .A(n369), .B(n370), .S0(n686), .Y(tag[18]) );
  MX4X2 U128 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n198), .S1(n703), .Y(
        n369) );
  INVX3 U129 ( .A(tag[23]), .Y(n1070) );
  INVX3 U130 ( .A(tag[24]), .Y(n1068) );
  INVX3 U131 ( .A(tag[14]), .Y(n1081) );
  CLKINVX1 U132 ( .A(tag[19]), .Y(n1074) );
  CLKMX2X2 U133 ( .A(n676), .B(n677), .S0(n697), .Y(n13) );
  MXI4X1 U134 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n198), .S1(n727), .Y(
        n677) );
  MXI4X1 U135 ( .A(\blocktag[0][20] ), .B(\blocktag[1][20] ), .C(
        \blocktag[2][20] ), .D(\blocktag[3][20] ), .S0(n200), .S1(n730), .Y(
        n676) );
  CLKMX2X2 U136 ( .A(n674), .B(n675), .S0(n697), .Y(n14) );
  MXI4X1 U137 ( .A(\blocktag[0][21] ), .B(\blocktag[1][21] ), .C(
        \blocktag[2][21] ), .D(\blocktag[3][21] ), .S0(n199), .S1(n730), .Y(
        n674) );
  CLKINVX1 U138 ( .A(blockdata[27]), .Y(n1253) );
  CLKINVX1 U139 ( .A(blockdata[31]), .Y(n1276) );
  CLKINVX1 U140 ( .A(blockdata[59]), .Y(n1249) );
  CLKINVX1 U141 ( .A(blockdata[91]), .Y(n1250) );
  CLKINVX1 U142 ( .A(blockdata[123]), .Y(n1252) );
  CLKINVX1 U143 ( .A(blockdata[127]), .Y(n1274) );
  NAND3BX1 U144 ( .AN(n769), .B(n320), .C(n774), .Y(n931) );
  OR2X1 U145 ( .A(n2), .B(n1248), .Y(n193) );
  OR2X1 U146 ( .A(n1275), .B(n1247), .Y(n194) );
  BUFX4 U147 ( .A(n755), .Y(n741) );
  BUFX12 U148 ( .A(N31), .Y(n731) );
  INVX16 U149 ( .A(n197), .Y(n199) );
  CLKBUFX3 U150 ( .A(N31), .Y(n755) );
  CLKBUFX3 U151 ( .A(N32), .Y(n730) );
  BUFX12 U152 ( .A(n702), .Y(n728) );
  CLKBUFX8 U153 ( .A(n686), .Y(n687) );
  CLKBUFX2 U154 ( .A(n198), .Y(n733) );
  BUFX6 U155 ( .A(n686), .Y(n688) );
  BUFX4 U156 ( .A(n688), .Y(n697) );
  AND2X2 U157 ( .A(n377), .B(proc_stall), .Y(n319) );
  CLKBUFX3 U158 ( .A(n687), .Y(n690) );
  BUFX4 U159 ( .A(n1275), .Y(n790) );
  CLKINVX1 U160 ( .A(N31), .Y(n855) );
  CLKINVX1 U161 ( .A(N32), .Y(n856) );
  MXI2X2 U162 ( .A(n12), .B(n204), .S0(n775), .Y(n9) );
  MXI2X2 U163 ( .A(n13), .B(n219), .S0(n775), .Y(n10) );
  MXI2X2 U164 ( .A(n14), .B(n215), .S0(n775), .Y(n11) );
  BUFX8 U165 ( .A(N32), .Y(n702) );
  CLKMX2X2 U166 ( .A(n680), .B(n681), .S0(n697), .Y(n12) );
  MX2X2 U167 ( .A(n678), .B(n679), .S0(n697), .Y(n15) );
  INVXL U168 ( .A(N33), .Y(n857) );
  CLKBUFX2 U169 ( .A(n755), .Y(n734) );
  NAND2XL U170 ( .A(n861), .B(blockdata[8]), .Y(n16) );
  NAND2X1 U171 ( .A(n861), .B(blockdata[16]), .Y(n17) );
  NAND2X1 U172 ( .A(n861), .B(blockdata[17]), .Y(n18) );
  NAND2X1 U173 ( .A(n861), .B(blockdata[18]), .Y(n19) );
  NAND2X1 U174 ( .A(n861), .B(blockdata[19]), .Y(n20) );
  NAND2X1 U175 ( .A(n861), .B(blockdata[20]), .Y(n21) );
  NAND2X1 U176 ( .A(n861), .B(blockdata[21]), .Y(n22) );
  NAND2X1 U177 ( .A(n861), .B(blockdata[22]), .Y(n23) );
  NAND2X1 U178 ( .A(n861), .B(blockdata[23]), .Y(n24) );
  NAND2X1 U179 ( .A(n861), .B(blockdata[24]), .Y(n25) );
  NAND2X1 U180 ( .A(n861), .B(blockdata[25]), .Y(n26) );
  NAND2X1 U181 ( .A(n861), .B(blockdata[32]), .Y(n27) );
  NAND2X1 U182 ( .A(n860), .B(blockdata[48]), .Y(n28) );
  NAND2X1 U183 ( .A(n860), .B(blockdata[49]), .Y(n29) );
  NAND2X1 U184 ( .A(n860), .B(blockdata[50]), .Y(n30) );
  NAND2X1 U185 ( .A(n860), .B(blockdata[51]), .Y(n31) );
  NAND2X1 U186 ( .A(n860), .B(blockdata[52]), .Y(n32) );
  NAND2X1 U187 ( .A(n860), .B(blockdata[53]), .Y(n33) );
  NAND2X1 U188 ( .A(n860), .B(blockdata[54]), .Y(n34) );
  NAND2X1 U189 ( .A(n860), .B(blockdata[55]), .Y(n35) );
  NAND2X1 U190 ( .A(n860), .B(blockdata[56]), .Y(n36) );
  NAND2X1 U191 ( .A(n860), .B(blockdata[57]), .Y(n37) );
  NAND2X1 U192 ( .A(n860), .B(blockdata[64]), .Y(n38) );
  NAND2X1 U193 ( .A(n860), .B(blockdata[65]), .Y(n39) );
  NAND2X1 U194 ( .A(n860), .B(blockdata[66]), .Y(n40) );
  NAND2X1 U195 ( .A(n860), .B(blockdata[67]), .Y(n41) );
  NAND2X1 U196 ( .A(n860), .B(blockdata[68]), .Y(n42) );
  NAND2X1 U197 ( .A(n860), .B(blockdata[80]), .Y(n43) );
  NAND2X1 U198 ( .A(n860), .B(blockdata[81]), .Y(n44) );
  NAND2X1 U199 ( .A(n860), .B(blockdata[82]), .Y(n45) );
  NAND2X1 U200 ( .A(n860), .B(blockdata[83]), .Y(n46) );
  AOI22X1 U201 ( .A0(tag[1]), .A1(mem_write), .B0(proc_addr[6]), .B1(mem_read), 
        .Y(n47) );
  AOI22X1 U202 ( .A0(tag[2]), .A1(mem_write), .B0(proc_addr[7]), .B1(mem_read), 
        .Y(n48) );
  AOI22X1 U203 ( .A0(tag[5]), .A1(mem_write), .B0(proc_addr[10]), .B1(mem_read), .Y(n49) );
  AOI22X1 U204 ( .A0(tag[6]), .A1(mem_write), .B0(proc_addr[11]), .B1(mem_read), .Y(n50) );
  AOI22X1 U205 ( .A0(tag[8]), .A1(mem_write), .B0(proc_addr[13]), .B1(mem_read), .Y(n51) );
  AOI22X1 U206 ( .A0(tag[10]), .A1(mem_write), .B0(proc_addr[15]), .B1(
        mem_read), .Y(n52) );
  AOI22X1 U207 ( .A0(tag[11]), .A1(mem_write), .B0(proc_addr[16]), .B1(
        mem_read), .Y(n53) );
  AOI22X1 U208 ( .A0(tag[12]), .A1(mem_write), .B0(proc_addr[17]), .B1(
        mem_read), .Y(n54) );
  AOI22X1 U209 ( .A0(tag[14]), .A1(mem_write), .B0(proc_addr[19]), .B1(
        mem_read), .Y(n55) );
  AOI22X1 U210 ( .A0(tag[16]), .A1(mem_write), .B0(proc_addr[21]), .B1(
        mem_read), .Y(n56) );
  AOI22X1 U211 ( .A0(tag[17]), .A1(mem_write), .B0(proc_addr[22]), .B1(
        mem_read), .Y(n57) );
  AOI22X1 U212 ( .A0(tag[18]), .A1(mem_write), .B0(proc_addr[23]), .B1(
        mem_read), .Y(n58) );
  AOI22X1 U213 ( .A0(tag[19]), .A1(mem_write), .B0(proc_addr[24]), .B1(
        mem_read), .Y(n59) );
  AOI22X1 U214 ( .A0(tag[22]), .A1(mem_write), .B0(proc_addr[27]), .B1(
        mem_read), .Y(n60) );
  AOI22X1 U215 ( .A0(tag[23]), .A1(mem_write), .B0(proc_addr[28]), .B1(
        mem_read), .Y(n61) );
  AOI22X1 U216 ( .A0(tag[24]), .A1(mem_write), .B0(proc_addr[29]), .B1(
        mem_read), .Y(n62) );
  MXI2X2 U217 ( .A(n1099), .B(n1098), .S0(n781), .Y(n63) );
  MXI2X2 U218 ( .A(n1097), .B(n1096), .S0(n782), .Y(n64) );
  MXI2X2 U219 ( .A(n1095), .B(n1094), .S0(n781), .Y(n65) );
  MXI2X2 U220 ( .A(n1093), .B(n1092), .S0(n782), .Y(n66) );
  MXI2X2 U221 ( .A(n1091), .B(n1090), .S0(n777), .Y(n67) );
  MXI2X2 U222 ( .A(n1089), .B(n1088), .S0(n319), .Y(n68) );
  MXI2X2 U223 ( .A(n1087), .B(n1086), .S0(n779), .Y(n69) );
  MXI2X2 U224 ( .A(n1085), .B(n1084), .S0(n780), .Y(n70) );
  MXI2X2 U225 ( .A(n1083), .B(n1082), .S0(n776), .Y(n71) );
  MXI2X2 U226 ( .A(n1076), .B(n1075), .S0(n775), .Y(n72) );
  MXI2X2 U227 ( .A(n1078), .B(n1077), .S0(n775), .Y(n73) );
  MXI2X2 U228 ( .A(n1070), .B(n1069), .S0(n775), .Y(n74) );
  MXI2X2 U229 ( .A(n1068), .B(n1067), .S0(n775), .Y(n75) );
  MXI2X2 U230 ( .A(n1081), .B(n1080), .S0(n775), .Y(n76) );
  MXI2X2 U231 ( .A(n1074), .B(n1073), .S0(n775), .Y(n77) );
  MXI2X2 U232 ( .A(n1072), .B(n1071), .S0(n775), .Y(n78) );
  BUFX4 U233 ( .A(n1314), .Y(mem_read) );
  NAND2X6 U234 ( .A(valid), .B(n893), .Y(n1109) );
  INVX3 U235 ( .A(tag[0]), .Y(n223) );
  NAND2X1 U236 ( .A(mem_write), .B(blockdata[0]), .Y(n79) );
  NAND2XL U237 ( .A(n859), .B(blockdata[84]), .Y(n80) );
  NAND2XL U238 ( .A(n859), .B(blockdata[85]), .Y(n81) );
  NAND2XL U239 ( .A(n859), .B(blockdata[86]), .Y(n82) );
  NAND2X1 U240 ( .A(n859), .B(blockdata[87]), .Y(n83) );
  NAND2XL U241 ( .A(n859), .B(blockdata[88]), .Y(n84) );
  NAND2XL U242 ( .A(n859), .B(blockdata[89]), .Y(n85) );
  NAND2XL U243 ( .A(n859), .B(blockdata[96]), .Y(n86) );
  NAND2XL U244 ( .A(n859), .B(blockdata[97]), .Y(n87) );
  NAND2X1 U245 ( .A(n859), .B(blockdata[98]), .Y(n88) );
  NAND2XL U246 ( .A(n859), .B(blockdata[99]), .Y(n89) );
  NAND2X1 U247 ( .A(n859), .B(blockdata[100]), .Y(n90) );
  NAND2X1 U248 ( .A(n859), .B(blockdata[101]), .Y(n91) );
  NAND2X1 U249 ( .A(n859), .B(blockdata[102]), .Y(n92) );
  NAND2X1 U250 ( .A(n859), .B(blockdata[103]), .Y(n93) );
  NAND2X1 U251 ( .A(n859), .B(blockdata[104]), .Y(n94) );
  NAND2X1 U252 ( .A(n859), .B(blockdata[112]), .Y(n95) );
  NAND2X1 U253 ( .A(n859), .B(blockdata[113]), .Y(n96) );
  NAND2X1 U254 ( .A(n859), .B(blockdata[114]), .Y(n97) );
  NAND2X1 U255 ( .A(n859), .B(blockdata[115]), .Y(n98) );
  NAND2X1 U256 ( .A(n859), .B(blockdata[116]), .Y(n99) );
  NAND2X1 U257 ( .A(n859), .B(blockdata[117]), .Y(n100) );
  NAND2X1 U258 ( .A(n859), .B(blockdata[118]), .Y(n101) );
  NAND2X1 U259 ( .A(n859), .B(blockdata[119]), .Y(n102) );
  NAND2X1 U260 ( .A(n859), .B(blockdata[120]), .Y(n103) );
  NAND2X1 U261 ( .A(n859), .B(blockdata[121]), .Y(n104) );
  CLKBUFX3 U262 ( .A(n728), .Y(n703) );
  AND4X1 U263 ( .A(n930), .B(n965), .C(n998), .D(n772), .Y(n105) );
  AOI21X2 U264 ( .A0(mem_ready), .A1(n1103), .B0(valid), .Y(n106) );
  MXI2X1 U265 ( .A(n666), .B(n667), .S0(n689), .Y(blockdata[1]) );
  MXI2X1 U266 ( .A(n662), .B(n663), .S0(n689), .Y(blockdata[3]) );
  CLKMX2X2 U267 ( .A(tag[3]), .B(proc_addr[8]), .S0(n775), .Y(n373) );
  CLKMX2X2 U268 ( .A(tag[18]), .B(proc_addr[23]), .S0(n775), .Y(n375) );
  CLKMX2X2 U269 ( .A(tag[2]), .B(proc_addr[7]), .S0(n778), .Y(n372) );
  INVX12 U270 ( .A(n48), .Y(mem_addr[5]) );
  INVX12 U271 ( .A(n47), .Y(mem_addr[4]) );
  INVX12 U272 ( .A(n57), .Y(mem_addr[20]) );
  INVX12 U273 ( .A(n60), .Y(mem_addr[25]) );
  INVXL U274 ( .A(n1319), .Y(n111) );
  INVX12 U275 ( .A(n111), .Y(mem_addr[6]) );
  AO22X1 U276 ( .A0(tag[3]), .A1(mem_write), .B0(proc_addr[8]), .B1(mem_read), 
        .Y(n1319) );
  INVXL U277 ( .A(n1318), .Y(n113) );
  INVX12 U278 ( .A(n113), .Y(mem_addr[7]) );
  AO22X1 U279 ( .A0(tag[4]), .A1(mem_write), .B0(proc_addr[9]), .B1(mem_read), 
        .Y(n1318) );
  INVX12 U280 ( .A(n49), .Y(mem_addr[8]) );
  INVX12 U281 ( .A(n50), .Y(mem_addr[9]) );
  INVXL U282 ( .A(n1317), .Y(n117) );
  INVX12 U283 ( .A(n117), .Y(mem_addr[10]) );
  AO22X1 U284 ( .A0(tag[7]), .A1(mem_write), .B0(proc_addr[12]), .B1(mem_read), 
        .Y(n1317) );
  INVX12 U285 ( .A(n51), .Y(mem_addr[11]) );
  INVXL U286 ( .A(n1316), .Y(n120) );
  INVX12 U287 ( .A(n120), .Y(mem_addr[12]) );
  AO22X1 U288 ( .A0(tag[9]), .A1(mem_write), .B0(proc_addr[14]), .B1(mem_read), 
        .Y(n1316) );
  INVX12 U289 ( .A(n52), .Y(mem_addr[13]) );
  INVX12 U290 ( .A(n53), .Y(mem_addr[14]) );
  INVX12 U291 ( .A(n54), .Y(mem_addr[15]) );
  INVX12 U292 ( .A(n55), .Y(mem_addr[17]) );
  INVX12 U293 ( .A(n56), .Y(mem_addr[19]) );
  INVX12 U294 ( .A(n58), .Y(mem_addr[21]) );
  INVX12 U295 ( .A(n59), .Y(mem_addr[22]) );
  INVX12 U296 ( .A(n61), .Y(mem_addr[26]) );
  INVX12 U297 ( .A(n62), .Y(mem_addr[27]) );
  INVX12 U298 ( .A(n79), .Y(mem_wdata[0]) );
  INVX12 U299 ( .A(n16), .Y(mem_wdata[8]) );
  CLKAND2X12 U300 ( .A(n861), .B(blockdata[9]), .Y(mem_wdata[9]) );
  CLKAND2X12 U301 ( .A(n861), .B(blockdata[10]), .Y(mem_wdata[10]) );
  CLKAND2X12 U302 ( .A(n861), .B(blockdata[11]), .Y(mem_wdata[11]) );
  CLKAND2X12 U303 ( .A(n861), .B(blockdata[12]), .Y(mem_wdata[12]) );
  CLKAND2X12 U304 ( .A(n861), .B(blockdata[13]), .Y(mem_wdata[13]) );
  CLKAND2X12 U305 ( .A(n861), .B(blockdata[14]), .Y(mem_wdata[14]) );
  CLKAND2X12 U306 ( .A(n861), .B(blockdata[15]), .Y(mem_wdata[15]) );
  INVX12 U307 ( .A(n17), .Y(mem_wdata[16]) );
  INVX12 U308 ( .A(n18), .Y(mem_wdata[17]) );
  INVX12 U309 ( .A(n19), .Y(mem_wdata[18]) );
  INVX12 U310 ( .A(n20), .Y(mem_wdata[19]) );
  INVX12 U311 ( .A(n21), .Y(mem_wdata[20]) );
  INVX12 U312 ( .A(n22), .Y(mem_wdata[21]) );
  INVX12 U313 ( .A(n23), .Y(mem_wdata[22]) );
  INVX12 U314 ( .A(n24), .Y(mem_wdata[23]) );
  INVX12 U315 ( .A(n25), .Y(mem_wdata[24]) );
  INVX12 U316 ( .A(n26), .Y(mem_wdata[25]) );
  CLKAND2X12 U317 ( .A(n861), .B(blockdata[27]), .Y(mem_wdata[27]) );
  CLKAND2X12 U318 ( .A(n861), .B(blockdata[28]), .Y(mem_wdata[28]) );
  CLKAND2X12 U319 ( .A(n861), .B(blockdata[29]), .Y(mem_wdata[29]) );
  CLKAND2X12 U320 ( .A(n861), .B(blockdata[30]), .Y(mem_wdata[30]) );
  CLKAND2X12 U321 ( .A(n861), .B(blockdata[31]), .Y(mem_wdata[31]) );
  INVX12 U322 ( .A(n27), .Y(mem_wdata[32]) );
  CLKAND2X12 U323 ( .A(n861), .B(blockdata[33]), .Y(mem_wdata[33]) );
  CLKAND2X12 U324 ( .A(n861), .B(blockdata[34]), .Y(mem_wdata[34]) );
  CLKAND2X12 U325 ( .A(n861), .B(blockdata[35]), .Y(mem_wdata[35]) );
  CLKAND2X12 U326 ( .A(n861), .B(blockdata[36]), .Y(mem_wdata[36]) );
  CLKAND2X12 U327 ( .A(n860), .B(blockdata[37]), .Y(mem_wdata[37]) );
  CLKAND2X12 U328 ( .A(n861), .B(blockdata[38]), .Y(mem_wdata[38]) );
  CLKAND2X12 U329 ( .A(n861), .B(blockdata[39]), .Y(mem_wdata[39]) );
  CLKAND2X12 U330 ( .A(n861), .B(blockdata[40]), .Y(mem_wdata[40]) );
  CLKAND2X12 U331 ( .A(n861), .B(blockdata[41]), .Y(mem_wdata[41]) );
  CLKAND2X12 U332 ( .A(n861), .B(blockdata[42]), .Y(mem_wdata[42]) );
  CLKAND2X12 U333 ( .A(n861), .B(blockdata[43]), .Y(mem_wdata[43]) );
  CLKAND2X12 U334 ( .A(n861), .B(blockdata[44]), .Y(mem_wdata[44]) );
  CLKAND2X12 U335 ( .A(n861), .B(blockdata[45]), .Y(mem_wdata[45]) );
  CLKAND2X12 U336 ( .A(n861), .B(blockdata[46]), .Y(mem_wdata[46]) );
  CLKBUFX8 U337 ( .A(mem_write), .Y(n861) );
  CLKAND2X12 U338 ( .A(n860), .B(blockdata[47]), .Y(mem_wdata[47]) );
  INVX12 U339 ( .A(n28), .Y(mem_wdata[48]) );
  INVX12 U340 ( .A(n29), .Y(mem_wdata[49]) );
  INVX12 U341 ( .A(n30), .Y(mem_wdata[50]) );
  INVX12 U342 ( .A(n31), .Y(mem_wdata[51]) );
  INVX12 U343 ( .A(n32), .Y(mem_wdata[52]) );
  INVX12 U344 ( .A(n33), .Y(mem_wdata[53]) );
  INVX12 U345 ( .A(n34), .Y(mem_wdata[54]) );
  INVX12 U346 ( .A(n35), .Y(mem_wdata[55]) );
  INVX12 U347 ( .A(n36), .Y(mem_wdata[56]) );
  INVX12 U348 ( .A(n37), .Y(mem_wdata[57]) );
  CLKAND2X12 U349 ( .A(n860), .B(blockdata[58]), .Y(mem_wdata[58]) );
  CLKAND2X12 U350 ( .A(n860), .B(blockdata[59]), .Y(mem_wdata[59]) );
  CLKAND2X12 U351 ( .A(n860), .B(blockdata[61]), .Y(mem_wdata[61]) );
  CLKAND2X12 U352 ( .A(n860), .B(blockdata[62]), .Y(mem_wdata[62]) );
  CLKAND2X12 U353 ( .A(n860), .B(blockdata[63]), .Y(mem_wdata[63]) );
  INVX12 U354 ( .A(n38), .Y(mem_wdata[64]) );
  INVX12 U355 ( .A(n39), .Y(mem_wdata[65]) );
  INVX12 U356 ( .A(n40), .Y(mem_wdata[66]) );
  INVX12 U357 ( .A(n41), .Y(mem_wdata[67]) );
  INVX12 U358 ( .A(n42), .Y(mem_wdata[68]) );
  CLKAND2X12 U359 ( .A(n860), .B(blockdata[69]), .Y(mem_wdata[69]) );
  CLKAND2X12 U360 ( .A(n860), .B(blockdata[70]), .Y(mem_wdata[70]) );
  CLKAND2X12 U361 ( .A(n860), .B(blockdata[71]), .Y(mem_wdata[71]) );
  CLKAND2X12 U362 ( .A(n860), .B(blockdata[72]), .Y(mem_wdata[72]) );
  CLKAND2X12 U363 ( .A(n860), .B(blockdata[73]), .Y(mem_wdata[73]) );
  CLKAND2X12 U364 ( .A(n860), .B(blockdata[74]), .Y(mem_wdata[74]) );
  CLKAND2X12 U365 ( .A(n860), .B(blockdata[75]), .Y(mem_wdata[75]) );
  CLKAND2X12 U366 ( .A(n860), .B(blockdata[76]), .Y(mem_wdata[76]) );
  CLKAND2X12 U367 ( .A(n860), .B(blockdata[77]), .Y(mem_wdata[77]) );
  CLKAND2X12 U368 ( .A(n860), .B(blockdata[78]), .Y(mem_wdata[78]) );
  CLKAND2X12 U369 ( .A(n860), .B(blockdata[79]), .Y(mem_wdata[79]) );
  CLKBUFX8 U370 ( .A(n1315), .Y(n860) );
  INVX12 U371 ( .A(n43), .Y(mem_wdata[80]) );
  INVX12 U372 ( .A(n44), .Y(mem_wdata[81]) );
  INVX12 U373 ( .A(n45), .Y(mem_wdata[82]) );
  INVX12 U374 ( .A(n46), .Y(mem_wdata[83]) );
  INVX12 U375 ( .A(n80), .Y(mem_wdata[84]) );
  INVX12 U376 ( .A(n81), .Y(mem_wdata[85]) );
  INVX12 U377 ( .A(n82), .Y(mem_wdata[86]) );
  INVX12 U378 ( .A(n83), .Y(mem_wdata[87]) );
  INVX12 U379 ( .A(n84), .Y(mem_wdata[88]) );
  INVX12 U380 ( .A(n85), .Y(mem_wdata[89]) );
  CLKAND2X12 U381 ( .A(n859), .B(blockdata[90]), .Y(mem_wdata[90]) );
  CLKAND2X12 U382 ( .A(n859), .B(blockdata[91]), .Y(mem_wdata[91]) );
  CLKAND2X12 U383 ( .A(n859), .B(blockdata[93]), .Y(mem_wdata[93]) );
  CLKAND2X12 U384 ( .A(n859), .B(blockdata[94]), .Y(mem_wdata[94]) );
  CLKAND2X12 U385 ( .A(n859), .B(blockdata[95]), .Y(mem_wdata[95]) );
  INVX12 U386 ( .A(n86), .Y(mem_wdata[96]) );
  INVX12 U387 ( .A(n87), .Y(mem_wdata[97]) );
  INVX12 U388 ( .A(n88), .Y(mem_wdata[98]) );
  INVX12 U389 ( .A(n89), .Y(mem_wdata[99]) );
  INVX12 U390 ( .A(n90), .Y(mem_wdata[100]) );
  INVX12 U391 ( .A(n91), .Y(mem_wdata[101]) );
  INVX12 U392 ( .A(n92), .Y(mem_wdata[102]) );
  INVX12 U393 ( .A(n93), .Y(mem_wdata[103]) );
  INVX12 U394 ( .A(n94), .Y(mem_wdata[104]) );
  CLKAND2X12 U395 ( .A(n859), .B(blockdata[105]), .Y(mem_wdata[105]) );
  CLKAND2X12 U396 ( .A(n859), .B(blockdata[106]), .Y(mem_wdata[106]) );
  CLKAND2X12 U397 ( .A(n859), .B(blockdata[107]), .Y(mem_wdata[107]) );
  CLKAND2X12 U398 ( .A(n859), .B(blockdata[108]), .Y(mem_wdata[108]) );
  CLKAND2X12 U399 ( .A(n859), .B(blockdata[109]), .Y(mem_wdata[109]) );
  CLKAND2X12 U400 ( .A(n859), .B(blockdata[110]), .Y(mem_wdata[110]) );
  CLKBUFX8 U401 ( .A(mem_write), .Y(n859) );
  CLKAND2X12 U402 ( .A(n859), .B(blockdata[111]), .Y(mem_wdata[111]) );
  INVX12 U403 ( .A(n95), .Y(mem_wdata[112]) );
  INVX12 U404 ( .A(n96), .Y(mem_wdata[113]) );
  INVX12 U405 ( .A(n97), .Y(mem_wdata[114]) );
  INVX12 U406 ( .A(n98), .Y(mem_wdata[115]) );
  INVX12 U407 ( .A(n99), .Y(mem_wdata[116]) );
  INVX12 U408 ( .A(n100), .Y(mem_wdata[117]) );
  INVX12 U409 ( .A(n101), .Y(mem_wdata[118]) );
  INVX12 U410 ( .A(n102), .Y(mem_wdata[119]) );
  INVX12 U411 ( .A(n103), .Y(mem_wdata[120]) );
  INVX12 U412 ( .A(n104), .Y(mem_wdata[121]) );
  CLKAND2X12 U413 ( .A(mem_write), .B(blockdata[123]), .Y(mem_wdata[123]) );
  CLKAND2X12 U414 ( .A(mem_write), .B(blockdata[125]), .Y(mem_wdata[125]) );
  CLKAND2X12 U415 ( .A(mem_write), .B(blockdata[126]), .Y(mem_wdata[126]) );
  CLKAND2X12 U416 ( .A(mem_write), .B(blockdata[127]), .Y(mem_wdata[127]) );
  INVX3 U417 ( .A(proc_reset), .Y(n865) );
  NAND2XL U418 ( .A(n1103), .B(n1109), .Y(n1064) );
  XOR2X2 U419 ( .A(n14), .B(proc_addr[26]), .Y(n883) );
  MX4X1 U420 ( .A(\blocktag[0][7] ), .B(\blocktag[1][7] ), .C(\blocktag[2][7] ), .D(\blocktag[3][7] ), .S0(n731), .S1(n727), .Y(n353) );
  MX4X1 U421 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n731), .S1(n727), .Y(
        n350) );
  MX4X1 U422 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n199), .S1(n727), .Y(
        n349) );
  MX4X1 U423 ( .A(\blocktag[4][8] ), .B(\blocktag[5][8] ), .C(\blocktag[6][8] ), .D(\blocktag[7][8] ), .S0(n731), .S1(n727), .Y(n352) );
  MX4X1 U424 ( .A(\blocktag[0][8] ), .B(\blocktag[1][8] ), .C(\blocktag[2][8] ), .D(\blocktag[3][8] ), .S0(n199), .S1(n727), .Y(n351) );
  MX4X1 U425 ( .A(\blocktag[4][7] ), .B(\blocktag[5][7] ), .C(\blocktag[6][7] ), .D(\blocktag[7][7] ), .S0(n199), .S1(n727), .Y(n354) );
  CLKMX2X6 U426 ( .A(n365), .B(n366), .S0(n698), .Y(tag[3]) );
  MX4X2 U427 ( .A(\blocktag[4][3] ), .B(\blocktag[5][3] ), .C(\blocktag[6][3] ), .D(\blocktag[7][3] ), .S0(n754), .S1(n728), .Y(n366) );
  MX4X2 U428 ( .A(\blocktag[0][3] ), .B(\blocktag[1][3] ), .C(\blocktag[2][3] ), .D(\blocktag[3][3] ), .S0(n754), .S1(n728), .Y(n365) );
  MX4X1 U429 ( .A(\blocktag[4][4] ), .B(\blocktag[5][4] ), .C(\blocktag[6][4] ), .D(\blocktag[7][4] ), .S0(n754), .S1(n728), .Y(n362) );
  MX4X1 U430 ( .A(\blocktag[0][4] ), .B(\blocktag[1][4] ), .C(\blocktag[2][4] ), .D(\blocktag[3][4] ), .S0(n754), .S1(n728), .Y(n361) );
  MXI4X4 U431 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(
        \blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n754), .S1(n728), .Y(n682) );
  BUFX8 U432 ( .A(N31), .Y(n732) );
  MX4X1 U433 ( .A(n343), .B(n344), .C(n345), .D(n346), .S0(n199), .S1(n726), 
        .Y(n681) );
  MX4X1 U434 ( .A(n339), .B(n340), .C(n341), .D(n342), .S0(n199), .S1(n726), 
        .Y(n680) );
  MX4X2 U435 ( .A(\blocktag[4][18] ), .B(\blocktag[6][18] ), .C(
        \blocktag[5][18] ), .D(\blocktag[7][18] ), .S0(N32), .S1(n200), .Y(
        n370) );
  MX4XL U436 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(\blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n731), .S1(n727), .Y(n360) );
  MX4X1 U437 ( .A(n188), .B(n189), .C(n190), .D(n191), .S0(n754), .S1(n728), 
        .Y(n683) );
  MX4X1 U438 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n754), .S1(n701), .Y(n325) );
  NOR2XL U439 ( .A(n857), .B(n856), .Y(n1313) );
  NAND3X6 U440 ( .A(n301), .B(n302), .C(n1256), .Y(proc_rdata[28]) );
  OR2X2 U441 ( .A(n1275), .B(n1257), .Y(n302) );
  OAI221X2 U442 ( .A0(n2), .A1(n1268), .B0(n1275), .B1(n1267), .C0(n1266), .Y(
        proc_rdata[30]) );
  OA22X4 U443 ( .A0(n3), .A1(n1260), .B0(n1), .B1(n1259), .Y(n1261) );
  OAI221X2 U444 ( .A0(n2), .A1(n1276), .B0(n1275), .B1(n1274), .C0(n1273), .Y(
        proc_rdata[31]) );
  NAND3X2 U445 ( .A(n193), .B(n194), .C(n1246), .Y(proc_rdata[26]) );
  OAI221X4 U446 ( .A0(n2), .A1(n1253), .B0(n1275), .B1(n1252), .C0(n1251), .Y(
        proc_rdata[27]) );
  CLKINVX1 U447 ( .A(blockdata[95]), .Y(n1271) );
  CLKINVX1 U448 ( .A(blockdata[63]), .Y(n1269) );
  MX4X1 U449 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(\blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n754), .S1(n728), .Y(n355) );
  MXI4X2 U450 ( .A(\blocktag[4][21] ), .B(\blocktag[5][21] ), .C(
        \blocktag[6][21] ), .D(\blocktag[7][21] ), .S0(n200), .S1(n727), .Y(
        n675) );
  MXI4X2 U451 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n200), .S1(n726), .Y(
        n679) );
  MX4X1 U452 ( .A(\blocktag[4][19] ), .B(\blocktag[5][19] ), .C(
        \blocktag[6][19] ), .D(\blocktag[7][19] ), .S0(n199), .S1(n727), .Y(
        n348) );
  XNOR2X4 U453 ( .A(n756), .B(tag[18]), .Y(n874) );
  MX4X1 U454 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(\blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n199), .S1(n727), .Y(n359) );
  MX4X1 U455 ( .A(\blocktag[4][6] ), .B(\blocktag[5][6] ), .C(\blocktag[6][6] ), .D(\blocktag[7][6] ), .S0(n731), .S1(n727), .Y(n364) );
  MXI2X4 U456 ( .A(n682), .B(n683), .S0(n698), .Y(tag[2]) );
  MXI2X1 U457 ( .A(n654), .B(n655), .S0(n695), .Y(blockdata[7]) );
  MXI2X1 U458 ( .A(n656), .B(n657), .S0(n691), .Y(blockdata[6]) );
  CLKAND2X12 U459 ( .A(n859), .B(blockdata[7]), .Y(mem_wdata[7]) );
  INVX1 U460 ( .A(blockdata[5]), .Y(n1143) );
  MXI2X1 U461 ( .A(n658), .B(n659), .S0(n689), .Y(blockdata[5]) );
  CLKAND2X12 U462 ( .A(n859), .B(blockdata[6]), .Y(mem_wdata[6]) );
  MXI2X1 U463 ( .A(n660), .B(n661), .S0(n695), .Y(blockdata[4]) );
  CLKAND2X12 U464 ( .A(n859), .B(blockdata[5]), .Y(mem_wdata[5]) );
  BUFX12 U465 ( .A(n1320), .Y(mem_addr[2]) );
  NOR2XL U466 ( .A(n318), .B(n857), .Y(n1320) );
  CLKAND2X12 U467 ( .A(n859), .B(blockdata[4]), .Y(mem_wdata[4]) );
  MXI2X1 U468 ( .A(n664), .B(n665), .S0(n691), .Y(blockdata[2]) );
  BUFX12 U469 ( .A(n1321), .Y(mem_addr[1]) );
  NOR2XL U470 ( .A(n318), .B(n856), .Y(n1321) );
  CLKAND2X12 U471 ( .A(n859), .B(blockdata[3]), .Y(mem_wdata[3]) );
  INVX12 U472 ( .A(n203), .Y(mem_addr[16]) );
  INVXL U473 ( .A(proc_addr[18]), .Y(n204) );
  INVXL U474 ( .A(mem_write), .Y(n205) );
  NOR2X1 U475 ( .A(n209), .B(n204), .Y(n206) );
  NOR2XL U476 ( .A(n205), .B(n12), .Y(n207) );
  NOR2XL U477 ( .A(n206), .B(n207), .Y(n203) );
  INVX12 U478 ( .A(n208), .Y(mem_addr[18]) );
  INVX1 U479 ( .A(mem_read), .Y(n209) );
  INVXL U480 ( .A(proc_addr[20]), .Y(n210) );
  INVXL U481 ( .A(mem_write), .Y(n211) );
  NOR2X1 U482 ( .A(n209), .B(n210), .Y(n212) );
  NOR2XL U483 ( .A(n211), .B(n15), .Y(n213) );
  NOR2XL U484 ( .A(n212), .B(n213), .Y(n208) );
  INVX12 U485 ( .A(n214), .Y(mem_addr[24]) );
  INVXL U486 ( .A(proc_addr[26]), .Y(n215) );
  NOR2X1 U487 ( .A(n209), .B(n215), .Y(n216) );
  NOR2XL U488 ( .A(n205), .B(n14), .Y(n217) );
  NOR2XL U489 ( .A(n216), .B(n217), .Y(n214) );
  INVX12 U490 ( .A(n218), .Y(mem_addr[23]) );
  INVXL U491 ( .A(proc_addr[25]), .Y(n219) );
  NOR2X1 U492 ( .A(n209), .B(n219), .Y(n220) );
  NOR2XL U493 ( .A(n211), .B(n13), .Y(n221) );
  NOR2XL U494 ( .A(n220), .B(n221), .Y(n218) );
  INVX12 U495 ( .A(n222), .Y(mem_addr[3]) );
  NOR2X1 U496 ( .A(n209), .B(n227), .Y(n224) );
  NOR2XL U497 ( .A(n205), .B(n223), .Y(n225) );
  NOR2XL U498 ( .A(n224), .B(n225), .Y(n222) );
  MXI2X4 U499 ( .A(n684), .B(n685), .S0(n698), .Y(tag[0]) );
  BUFX12 U500 ( .A(n1322), .Y(mem_addr[0]) );
  NOR2XL U501 ( .A(n318), .B(n855), .Y(n1322) );
  CLKAND2X12 U502 ( .A(n860), .B(blockdata[2]), .Y(mem_wdata[2]) );
  CLKAND2X12 U503 ( .A(n860), .B(blockdata[1]), .Y(mem_wdata[1]) );
  CLKAND2X12 U504 ( .A(n860), .B(blockdata[60]), .Y(mem_wdata[60]) );
  CLKAND2X12 U505 ( .A(n861), .B(blockdata[26]), .Y(mem_wdata[26]) );
  CLKAND2X12 U506 ( .A(mem_write), .B(blockdata[124]), .Y(mem_wdata[124]) );
  CLKAND2X12 U507 ( .A(mem_write), .B(blockdata[122]), .Y(mem_wdata[122]) );
  CLKAND2X12 U508 ( .A(n859), .B(blockdata[92]), .Y(mem_wdata[92]) );
  BUFX20 U509 ( .A(n731), .Y(n754) );
  BUFX20 U510 ( .A(N33), .Y(n686) );
  NAND2X2 U511 ( .A(tag[0]), .B(n227), .Y(n229) );
  INVXL U512 ( .A(proc_addr[5]), .Y(n227) );
  CLKBUFX2 U513 ( .A(n732), .Y(n752) );
  BUFX20 U514 ( .A(n732), .Y(n753) );
  CLKBUFX4 U515 ( .A(n200), .Y(n749) );
  MXI4XL U516 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n736), .S1(n709), .Y(n378) );
  MXI4X1 U517 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n736), .S1(n709), .Y(n379) );
  BUFX4 U518 ( .A(n752), .Y(n736) );
  AND2X2 U519 ( .A(n320), .B(n965), .Y(n308) );
  INVX1 U520 ( .A(proc_addr[1]), .Y(n1112) );
  CLKBUFX3 U521 ( .A(n741), .Y(n751) );
  BUFX4 U522 ( .A(n733), .Y(n747) );
  CLKBUFX3 U523 ( .A(n703), .Y(n725) );
  BUFX4 U524 ( .A(n708), .Y(n709) );
  OA22XL U525 ( .A0(n788), .A1(n1130), .B0(n7), .B1(n1129), .Y(n1131) );
  INVX1 U526 ( .A(blockdata[73]), .Y(n1160) );
  MXI2X2 U527 ( .A(n616), .B(n617), .S0(n696), .Y(blockdata[26]) );
  MX4XL U528 ( .A(n249), .B(n250), .C(n251), .D(n252), .S0(n741), .S1(n713), 
        .Y(n442) );
  MX4XL U529 ( .A(n253), .B(n254), .C(n255), .D(n256), .S0(n741), .S1(n713), 
        .Y(n443) );
  MXI4XL U530 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n742), .S1(n715), .Y(n510) );
  MXI4XL U531 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n742), .S1(n715), .Y(n511) );
  CLKBUFX3 U532 ( .A(n752), .Y(n743) );
  BUFX20 U533 ( .A(n687), .Y(n698) );
  CLKBUFX2 U534 ( .A(n319), .Y(n783) );
  OAI221X1 U535 ( .A0(n6), .A1(n1163), .B0(n790), .B1(n1162), .C0(n1161), .Y(
        proc_rdata[9]) );
  OA22XL U536 ( .A0(n788), .A1(n1160), .B0(n8), .B1(n1159), .Y(n1161) );
  OAI221XL U537 ( .A0(n5), .A1(n1238), .B0(n1275), .B1(n1237), .C0(n1236), .Y(
        proc_rdata[24]) );
  OA22X1 U538 ( .A0(n788), .A1(n1235), .B0(n785), .B1(n1234), .Y(n1236) );
  OAI221XL U539 ( .A0(n5), .A1(n1243), .B0(n1275), .B1(n1242), .C0(n1241), .Y(
        proc_rdata[25]) );
  OA22X1 U540 ( .A0(n789), .A1(n1240), .B0(n786), .B1(n1239), .Y(n1241) );
  MXI4X1 U541 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n749), .S1(n724), .Y(n617) );
  MXI4X1 U542 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n749), .S1(n724), .Y(n616) );
  MXI2X1 U543 ( .A(n452), .B(n453), .S0(n691), .Y(blockdata[90]) );
  MXI2X2 U544 ( .A(n388), .B(n389), .S0(n690), .Y(blockdata[122]) );
  MXI4X1 U545 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n736), .S1(n710), .Y(n389) );
  MXI4X1 U546 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n737), .S1(n710), .Y(n388) );
  MX4X1 U547 ( .A(n245), .B(n246), .C(n247), .D(n248), .S0(n745), .S1(n717), 
        .Y(n543) );
  MX4X1 U548 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n745), .S1(n717), 
        .Y(n542) );
  MXI4X1 U549 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n749), .S1(n723), .Y(n609) );
  MXI4X1 U550 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n749), .S1(n723), .Y(n608) );
  MXI2X1 U551 ( .A(n552), .B(n553), .S0(n693), .Y(blockdata[58]) );
  MXI4XL U552 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n745), .S1(n718), .Y(n549) );
  MXI4XL U553 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n749), .S1(n723), .Y(n613) );
  MXI4XL U554 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n736), .S1(n709), .Y(n385) );
  MX4XL U555 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(n739), .S1(n711), 
        .Y(n423) );
  MXI4XL U556 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n739), .S1(n711), .Y(n422) );
  MXI4X1 U557 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n739), .S1(n711), .Y(n419) );
  MXI4X1 U558 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n739), .S1(n711), .Y(n418) );
  MX4XL U559 ( .A(n273), .B(n274), .C(n275), .D(n276), .S0(n747), .S1(n721), 
        .Y(n587) );
  MXI4XL U560 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n747), .S1(n721), .Y(n586) );
  MX4XL U561 ( .A(n277), .B(n278), .C(n279), .D(n280), .S0(n743), .S1(n716), 
        .Y(n523) );
  MXI4XL U562 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n743), .S1(n716), .Y(n522) );
  MXI4X1 U563 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n747), .S1(n721), .Y(n583) );
  MXI4X1 U564 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n747), .S1(n721), .Y(n582) );
  MXI4X1 U565 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n743), .S1(n715), .Y(n519) );
  MXI4X1 U566 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n743), .S1(n715), .Y(n518) );
  BUFX8 U567 ( .A(n733), .Y(n745) );
  CLKBUFX2 U568 ( .A(n700), .Y(n706) );
  CLKBUFX2 U569 ( .A(n730), .Y(n707) );
  CLKBUFX2 U570 ( .A(n701), .Y(n704) );
  BUFX4 U571 ( .A(n735), .Y(n739) );
  CLKBUFX2 U572 ( .A(n729), .Y(n705) );
  CLKBUFX2 U573 ( .A(n303), .Y(n771) );
  CLKBUFX2 U574 ( .A(n687), .Y(n689) );
  CLKBUFX2 U575 ( .A(n702), .Y(n729) );
  CLKBUFX2 U576 ( .A(n964), .Y(n762) );
  OA22XL U577 ( .A0(n788), .A1(n1135), .B0(n8), .B1(n1134), .Y(n1136) );
  OA22XL U578 ( .A0(n788), .A1(n1150), .B0(n7), .B1(n1149), .Y(n1151) );
  OA22XL U579 ( .A0(n788), .A1(n1115), .B0(n8), .B1(n1114), .Y(n1116) );
  OA22XL U580 ( .A0(n788), .A1(n1120), .B0(n7), .B1(n1119), .Y(n1121) );
  CLKBUFX2 U581 ( .A(n784), .Y(n786) );
  OA22XL U582 ( .A0(n789), .A1(n1195), .B0(n785), .B1(n1194), .Y(n1196) );
  OA22XL U583 ( .A0(n789), .A1(n1200), .B0(n785), .B1(n1199), .Y(n1201) );
  OA22XL U584 ( .A0(n789), .A1(n1205), .B0(n786), .B1(n1204), .Y(n1206) );
  OA22XL U585 ( .A0(n789), .A1(n1210), .B0(n785), .B1(n1209), .Y(n1211) );
  OA22XL U586 ( .A0(n789), .A1(n1215), .B0(n786), .B1(n1214), .Y(n1216) );
  OA22XL U587 ( .A0(n789), .A1(n1220), .B0(n785), .B1(n1219), .Y(n1221) );
  OA22XL U588 ( .A0(n789), .A1(n1225), .B0(n785), .B1(n1224), .Y(n1226) );
  OA22XL U589 ( .A0(n789), .A1(n1230), .B0(n786), .B1(n1229), .Y(n1231) );
  NAND3BX4 U590 ( .AN(n1109), .B(n863), .C(n1108), .Y(n1113) );
  INVX3 U591 ( .A(blockdata[29]), .Y(n1263) );
  INVX3 U592 ( .A(blockdata[30]), .Y(n1268) );
  INVX3 U593 ( .A(blockdata[125]), .Y(n1262) );
  INVX3 U594 ( .A(blockdata[126]), .Y(n1267) );
  INVX3 U595 ( .A(blockdata[93]), .Y(n1260) );
  INVX3 U596 ( .A(blockdata[94]), .Y(n1265) );
  INVX3 U597 ( .A(blockdata[61]), .Y(n1259) );
  INVX3 U598 ( .A(blockdata[62]), .Y(n1264) );
  CLKBUFX2 U599 ( .A(n3), .Y(n787) );
  NAND4BXL U600 ( .AN(n1105), .B(n1104), .C(n1103), .D(n1102), .Y(n1106) );
  INVX1 U601 ( .A(blockdata[105]), .Y(n1162) );
  INVX1 U602 ( .A(blockdata[72]), .Y(n1155) );
  INVX1 U603 ( .A(blockdata[41]), .Y(n1159) );
  INVX1 U604 ( .A(blockdata[40]), .Y(n1154) );
  INVX1 U605 ( .A(blockdata[43]), .Y(n1169) );
  AND2X1 U606 ( .A(n1106), .B(n1107), .Y(n318) );
  INVX1 U607 ( .A(blockdata[9]), .Y(n1163) );
  INVX1 U608 ( .A(blockdata[11]), .Y(n1173) );
  INVX1 U609 ( .A(blockdata[10]), .Y(n1168) );
  INVX1 U610 ( .A(blockdata[15]), .Y(n1193) );
  INVX1 U611 ( .A(blockdata[12]), .Y(n1178) );
  INVX1 U612 ( .A(blockdata[14]), .Y(n1188) );
  INVX1 U613 ( .A(blockdata[13]), .Y(n1183) );
  INVX1 U614 ( .A(blockdata[106]), .Y(n1167) );
  INVX1 U615 ( .A(blockdata[111]), .Y(n1192) );
  INVX1 U616 ( .A(blockdata[108]), .Y(n1177) );
  INVX1 U617 ( .A(blockdata[110]), .Y(n1187) );
  INVX1 U618 ( .A(blockdata[109]), .Y(n1182) );
  INVX1 U619 ( .A(blockdata[75]), .Y(n1170) );
  INVX1 U620 ( .A(blockdata[74]), .Y(n1165) );
  INVX1 U621 ( .A(blockdata[79]), .Y(n1190) );
  INVX1 U622 ( .A(blockdata[76]), .Y(n1175) );
  INVX1 U623 ( .A(blockdata[78]), .Y(n1185) );
  INVX1 U624 ( .A(blockdata[69]), .Y(n1140) );
  INVX1 U625 ( .A(blockdata[77]), .Y(n1180) );
  INVX1 U626 ( .A(blockdata[70]), .Y(n1145) );
  INVX1 U627 ( .A(blockdata[71]), .Y(n1150) );
  INVX1 U628 ( .A(blockdata[42]), .Y(n1164) );
  INVX1 U629 ( .A(blockdata[47]), .Y(n1189) );
  INVX1 U630 ( .A(blockdata[35]), .Y(n1129) );
  INVX1 U631 ( .A(blockdata[46]), .Y(n1184) );
  INVX1 U632 ( .A(blockdata[44]), .Y(n1174) );
  INVX1 U633 ( .A(blockdata[34]), .Y(n1124) );
  INVX1 U634 ( .A(blockdata[45]), .Y(n1179) );
  INVX1 U635 ( .A(blockdata[36]), .Y(n1134) );
  INVX1 U636 ( .A(blockdata[37]), .Y(n1139) );
  INVX1 U637 ( .A(blockdata[33]), .Y(n1119) );
  INVX1 U638 ( .A(blockdata[38]), .Y(n1144) );
  INVX1 U639 ( .A(blockdata[39]), .Y(n1149) );
  NOR2XL U640 ( .A(n856), .B(N33), .Y(n1311) );
  AND2XL U641 ( .A(n1310), .B(n855), .Y(n321) );
  AND2XL U642 ( .A(n1312), .B(n855), .Y(n322) );
  AND2XL U643 ( .A(n1311), .B(n855), .Y(n323) );
  AND2XL U644 ( .A(n1313), .B(n855), .Y(n324) );
  INVX1 U645 ( .A(proc_addr[23]), .Y(n756) );
  MXI4XL U646 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n749), .S1(n723), .Y(n614) );
  MXI4XL U647 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n749), .S1(n723), .Y(n615) );
  MX4XL U648 ( .A(n257), .B(n258), .C(n259), .D(n260), .S0(n741), .S1(n713), 
        .Y(n446) );
  MX4XL U649 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n741), .S1(n713), 
        .Y(n447) );
  MX4XL U650 ( .A(n265), .B(n266), .C(n267), .D(n268), .S0(n741), .S1(n713), 
        .Y(n444) );
  MX4XL U651 ( .A(n269), .B(n270), .C(n271), .D(n272), .S0(n741), .S1(n713), 
        .Y(n445) );
  MXI4XL U652 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n741), .S1(n714), .Y(n453) );
  MXI4XL U653 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n741), .S1(n714), .Y(n452) );
  MXI4XL U654 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n736), .S1(n709), .Y(n386) );
  MXI4XL U655 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n736), .S1(n709), .Y(n387) );
  MXI4XL U656 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n736), .S1(n709), .Y(n382) );
  MXI4XL U657 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n736), .S1(n709), .Y(n383) );
  MXI4XL U658 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n736), .S1(n709), .Y(n380) );
  MXI4XL U659 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n736), .S1(n709), .Y(n381) );
  MXI4XL U660 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n745), .S1(n718), .Y(n552) );
  MXI4XL U661 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n745), .S1(n718), .Y(n553) );
  NAND3BXL U662 ( .AN(mem_ready), .B(proc_stall), .C(n1105), .Y(n1107) );
  INVX1 U663 ( .A(proc_addr[0]), .Y(n1111) );
  AND2XL U664 ( .A(proc_addr[0]), .B(proc_addr[1]), .Y(n376) );
  NAND2XL U665 ( .A(mem_rdata[0]), .B(n775), .Y(n1061) );
  MXI2XL U666 ( .A(n652), .B(n653), .S0(n694), .Y(blockdata[8]) );
  MXI4XL U667 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n746), .S1(n707), .Y(n662) );
  MXI4XL U668 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n734), .S1(n720), .Y(n663) );
  MXI4XL U669 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n742), .S1(n715), .Y(n660) );
  MXI4XL U670 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n743), .S1(n725), .Y(n661) );
  MXI4XL U671 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n747), .S1(n705), .Y(n656) );
  MXI4XL U672 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n739), .S1(n706), .Y(n657) );
  MXI4XL U673 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n739), .S1(n712), .Y(n654) );
  MXI4XL U674 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n750), .S1(n725), .Y(n655) );
  MXI2XL U675 ( .A(n424), .B(n425), .S0(n691), .Y(blockdata[104]) );
  MXI4XL U676 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n747), .S1(n721), .Y(n584) );
  MXI4XL U677 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n747), .S1(n721), .Y(n585) );
  MXI4XL U678 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n743), .S1(n716), .Y(n520) );
  MXI4XL U679 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n743), .S1(n716), .Y(n521) );
  MX4X1 U680 ( .A(n285), .B(n286), .C(n287), .D(n288), .S0(n746), .S1(n720), 
        .Y(n575) );
  MXI4XL U681 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n739), .S1(n711), .Y(n420) );
  MXI4XL U682 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n739), .S1(n711), .Y(n421) );
  MXI4XL U683 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n748), .S1(n722), .Y(n598) );
  MXI4XL U684 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n748), .S1(n722), .Y(n599) );
  MX4X1 U685 ( .A(n289), .B(n290), .C(n291), .D(n292), .S0(n738), .S1(n716), 
        .Y(n411) );
  MXI2XL U686 ( .A(n434), .B(n435), .S0(n693), .Y(blockdata[99]) );
  MXI4XL U687 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n740), .S1(n712), .Y(n434) );
  MXI4XL U688 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n740), .S1(n712), .Y(n435) );
  MXI4XL U689 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n746), .S1(n720), .Y(n576) );
  MXI4XL U690 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n746), .S1(n720), .Y(n577) );
  MXI2XL U691 ( .A(n534), .B(n535), .S0(n693), .Y(blockdata[67]) );
  MXI4XL U692 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n744), .S1(n717), .Y(n534) );
  MXI4XL U693 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n744), .S1(n717), .Y(n535) );
  MXI4XL U694 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n747), .S1(n721), .Y(n580) );
  MXI4XL U695 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n746), .S1(n721), .Y(n581) );
  MXI4XL U696 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n746), .S1(n720), .Y(n578) );
  MXI4XL U697 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n746), .S1(n720), .Y(n579) );
  MXI4XL U698 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n743), .S1(n715), .Y(n516) );
  MXI4XL U699 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n743), .S1(n715), .Y(n517) );
  MXI4XL U700 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n739), .S1(n711), .Y(n416) );
  MXI4XL U701 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n739), .S1(n711), .Y(n417) );
  MXI4XL U702 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n748), .S1(n722), .Y(n600) );
  MXI4XL U703 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n748), .S1(n722), .Y(n601) );
  MXI4XL U704 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n742), .S1(n715), .Y(n512) );
  MXI4XL U705 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n742), .S1(n715), .Y(n513) );
  MXI2XL U706 ( .A(n436), .B(n437), .S0(n693), .Y(blockdata[98]) );
  MXI4XL U707 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n740), .S1(n713), .Y(n436) );
  MXI4XL U708 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n740), .S1(n713), .Y(n437) );
  MXI2XL U709 ( .A(n536), .B(n537), .S0(n693), .Y(blockdata[66]) );
  MXI4XL U710 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n744), .S1(n717), .Y(n536) );
  MXI4XL U711 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n744), .S1(n717), .Y(n537) );
  MXI4XL U712 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n738), .S1(n711), .Y(n412) );
  MXI4XL U713 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n738), .S1(n711), .Y(n413) );
  MXI4XL U714 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n742), .S1(n715), .Y(n514) );
  MXI4XL U715 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n742), .S1(n715), .Y(n515) );
  MXI4XL U716 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n748), .S1(n722), .Y(n596) );
  MXI4XL U717 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n748), .S1(n722), .Y(n597) );
  MXI4XL U718 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n748), .S1(n722), .Y(n594) );
  MXI4XL U719 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n748), .S1(n722), .Y(n595) );
  MXI4XL U720 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n739), .S1(n711), .Y(n414) );
  MXI4XL U721 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n738), .S1(n711), .Y(n415) );
  MXI4XL U722 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n747), .S1(n719), .Y(n646) );
  MXI4XL U723 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n739), .S1(n725), .Y(n647) );
  MXI2XL U724 ( .A(n432), .B(n433), .S0(n695), .Y(blockdata[100]) );
  MXI4XL U725 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n740), .S1(n712), .Y(n432) );
  MXI4XL U726 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n740), .S1(n712), .Y(n433) );
  MXI2XL U727 ( .A(n604), .B(n605), .S0(n696), .Y(blockdata[32]) );
  MXI4XL U728 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n748), .S1(n723), .Y(n604) );
  MXI4XL U729 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n748), .S1(n723), .Y(n605) );
  MXI4XL U730 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n748), .S1(n722), .Y(n602) );
  MXI4XL U731 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n748), .S1(n722), .Y(n603) );
  MXI2XL U732 ( .A(n532), .B(n533), .S0(n693), .Y(blockdata[68]) );
  MXI4XL U733 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n744), .S1(n717), .Y(n532) );
  MXI4XL U734 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n744), .S1(n717), .Y(n533) );
  MXI2XL U735 ( .A(n430), .B(n431), .S0(n694), .Y(blockdata[101]) );
  MXI4XL U736 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n740), .S1(n712), .Y(n430) );
  MXI4XL U737 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n740), .S1(n712), .Y(n431) );
  MXI4XL U738 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n747), .S1(n722), .Y(n592) );
  MXI4XL U739 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n747), .S1(n722), .Y(n593) );
  MXI4XL U740 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n744), .S1(n716), .Y(n530) );
  MXI4XL U741 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n744), .S1(n716), .Y(n531) );
  MXI2XL U742 ( .A(n440), .B(n441), .S0(n693), .Y(blockdata[96]) );
  MXI4XL U743 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n741), .S1(n713), .Y(n440) );
  MXI4XL U744 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n740), .S1(n713), .Y(n441) );
  MXI2XL U745 ( .A(n438), .B(n439), .S0(n691), .Y(blockdata[97]) );
  MXI4XL U746 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n740), .S1(n713), .Y(n438) );
  MXI4XL U747 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n740), .S1(n713), .Y(n439) );
  MXI2XL U748 ( .A(n428), .B(n429), .S0(n693), .Y(blockdata[102]) );
  MXI4XL U749 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n740), .S1(n712), .Y(n428) );
  MXI4XL U750 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n740), .S1(n712), .Y(n429) );
  MXI2XL U751 ( .A(n540), .B(n541), .S0(n693), .Y(blockdata[64]) );
  MXI4XL U752 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n744), .S1(n717), .Y(n540) );
  MXI4XL U753 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n744), .S1(n717), .Y(n541) );
  MXI2XL U754 ( .A(n538), .B(n539), .S0(n693), .Y(blockdata[65]) );
  MXI4XL U755 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n744), .S1(n717), .Y(n538) );
  MXI4XL U756 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n744), .S1(n717), .Y(n539) );
  MXI4XL U757 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n744), .S1(n716), .Y(n528) );
  MXI4XL U758 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n743), .S1(n716), .Y(n529) );
  MXI4XL U759 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n747), .S1(n721), .Y(n590) );
  MXI4XL U760 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n747), .S1(n721), .Y(n591) );
  MXI4XL U761 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n750), .S1(n725), .Y(n648) );
  MXI4XL U762 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n747), .S1(n719), .Y(n649) );
  MXI2XL U763 ( .A(n426), .B(n427), .S0(n691), .Y(blockdata[103]) );
  MXI4XL U764 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n739), .S1(n712), .Y(n426) );
  MXI4XL U765 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n739), .S1(n712), .Y(n427) );
  MXI4XL U766 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n743), .S1(n716), .Y(n526) );
  MXI4XL U767 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n743), .S1(n716), .Y(n527) );
  MX4XL U768 ( .A(n293), .B(n294), .C(n295), .D(n296), .S0(n751), .S1(n725), 
        .Y(n644) );
  MX4XL U769 ( .A(n297), .B(n298), .C(n299), .D(n300), .S0(n751), .S1(n725), 
        .Y(n645) );
  MXI4XL U770 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n751), .S1(n712), .Y(n640) );
  MXI4XL U771 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n751), .S1(n712), .Y(n641) );
  MXI4XL U772 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n751), .S1(n725), .Y(n642) );
  MXI4XL U773 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n751), .S1(n725), .Y(n643) );
  INVXL U774 ( .A(proc_addr[17]), .Y(n1082) );
  MX2XL U775 ( .A(n223), .B(n227), .S0(n775), .Y(n1100) );
  INVXL U776 ( .A(proc_addr[6]), .Y(n1098) );
  INVXL U777 ( .A(proc_addr[9]), .Y(n1096) );
  INVXL U778 ( .A(proc_addr[11]), .Y(n1094) );
  INVXL U779 ( .A(proc_addr[12]), .Y(n1092) );
  INVXL U780 ( .A(proc_addr[13]), .Y(n1090) );
  INVXL U781 ( .A(proc_addr[14]), .Y(n1088) );
  INVXL U782 ( .A(proc_addr[15]), .Y(n1086) );
  INVXL U783 ( .A(proc_addr[16]), .Y(n1084) );
  MX2XL U784 ( .A(n15), .B(n210), .S0(n775), .Y(n1079) );
  INVXL U785 ( .A(proc_addr[21]), .Y(n1077) );
  INVXL U786 ( .A(proc_addr[22]), .Y(n1075) );
  INVXL U787 ( .A(proc_addr[24]), .Y(n1073) );
  INVXL U788 ( .A(proc_addr[27]), .Y(n1071) );
  INVXL U789 ( .A(proc_addr[28]), .Y(n1069) );
  INVXL U790 ( .A(proc_addr[29]), .Y(n1067) );
  OAI211XL U791 ( .A0(mem_ready), .A1(valid), .B0(n894), .C0(n1103), .Y(n895)
         );
  INVX3 U792 ( .A(n895), .Y(n930) );
  MXI4XL U793 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n746), .S1(n704), .Y(n664) );
  MXI4XL U794 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n740), .S1(n721), .Y(n665) );
  MXI2XL U795 ( .A(n668), .B(n669), .S0(N33), .Y(blockdata[0]) );
  MXI4XL U796 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n743), .S1(n720), .Y(n668) );
  MXI4XL U797 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n743), .S1(n711), .Y(n669) );
  MXI4XL U798 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n734), .S1(n722), .Y(n666) );
  MXI4XL U799 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n740), .S1(n720), .Y(n667) );
  MXI4XL U800 ( .A(\block[0][5] ), .B(\block[1][5] ), .C(\block[2][5] ), .D(
        \block[3][5] ), .S0(n740), .S1(n712), .Y(n658) );
  MXI4XL U801 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n750), .S1(n716), .Y(n659) );
  AND2XL U802 ( .A(mem_ready), .B(n1105), .Y(n377) );
  MXI2XL U803 ( .A(n508), .B(n509), .S0(n692), .Y(blockdata[80]) );
  MXI4XL U804 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n742), .S1(n715), .Y(n509) );
  MXI4XL U805 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n742), .S1(n715), .Y(n508) );
  MXI2XL U806 ( .A(n572), .B(n573), .S0(n694), .Y(blockdata[48]) );
  MXI4XL U807 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n746), .S1(n720), .Y(n573) );
  MXI4XL U808 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n746), .S1(n720), .Y(n572) );
  MXI2XL U809 ( .A(n506), .B(n507), .S0(n691), .Y(blockdata[81]) );
  MXI4XL U810 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n742), .S1(n705), .Y(n507) );
  MXI4XL U811 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n742), .S1(n712), .Y(n506) );
  MXI2XL U812 ( .A(n570), .B(n571), .S0(n694), .Y(blockdata[49]) );
  MXI4XL U813 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n746), .S1(n720), .Y(n571) );
  MXI4XL U814 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n746), .S1(n720), .Y(n570) );
  MXI2XL U815 ( .A(n504), .B(n505), .S0(n691), .Y(blockdata[82]) );
  MXI4XL U816 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n742), .S1(n712), .Y(n505) );
  MXI4XL U817 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n742), .S1(n715), .Y(n504) );
  MXI2XL U818 ( .A(n568), .B(n569), .S0(n694), .Y(blockdata[50]) );
  MXI4XL U819 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n746), .S1(n720), .Y(n569) );
  MXI4XL U820 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n746), .S1(n720), .Y(n568) );
  MXI2XL U821 ( .A(n566), .B(n567), .S0(n694), .Y(blockdata[51]) );
  MXI2XL U822 ( .A(n466), .B(n502), .S0(n691), .Y(blockdata[83]) );
  MXI4XL U823 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n742), .S1(n720), .Y(n466) );
  MXI2XL U824 ( .A(n564), .B(n565), .S0(n694), .Y(blockdata[52]) );
  MXI2XL U825 ( .A(n464), .B(n465), .S0(n691), .Y(blockdata[84]) );
  MXI2XL U826 ( .A(n562), .B(n563), .S0(n694), .Y(blockdata[53]) );
  MXI2XL U827 ( .A(n462), .B(n463), .S0(n691), .Y(blockdata[85]) );
  MXI2XL U828 ( .A(n560), .B(n561), .S0(n694), .Y(blockdata[54]) );
  MXI2XL U829 ( .A(n460), .B(n461), .S0(n691), .Y(blockdata[86]) );
  MXI2XL U830 ( .A(n558), .B(n559), .S0(n694), .Y(blockdata[55]) );
  MXI2XL U831 ( .A(n458), .B(n459), .S0(n691), .Y(blockdata[87]) );
  MXI4XL U832 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n747), .S1(n714), .Y(n459) );
  MXI4XL U833 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n752), .S1(n714), .Y(n458) );
  MXI2XL U834 ( .A(n556), .B(n557), .S0(n694), .Y(blockdata[56]) );
  MXI2XL U835 ( .A(n456), .B(n457), .S0(n691), .Y(blockdata[88]) );
  MXI4XL U836 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n735), .S1(n714), .Y(n457) );
  MXI4XL U837 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n752), .S1(n714), .Y(n456) );
  MXI2XL U838 ( .A(n554), .B(n555), .S0(n693), .Y(blockdata[57]) );
  MXI4XL U839 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n745), .S1(n718), .Y(n555) );
  MXI4XL U840 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n734), .S1(n718), .Y(n554) );
  MXI2XL U841 ( .A(n454), .B(n455), .S0(n691), .Y(blockdata[89]) );
  MXI4XL U842 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n734), .S1(n714), .Y(n455) );
  MXI4XL U843 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n751), .S1(n714), .Y(n454) );
  MXI2XL U844 ( .A(n408), .B(n409), .S0(n690), .Y(blockdata[112]) );
  MXI4XL U845 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n738), .S1(n719), .Y(n409) );
  MXI4XL U846 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n738), .S1(n719), .Y(n408) );
  MXI2XL U847 ( .A(n636), .B(n637), .S0(n692), .Y(blockdata[16]) );
  MXI4XL U848 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n751), .S1(n725), .Y(n637) );
  MXI4XL U849 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n751), .S1(n725), .Y(n636) );
  MXI2XL U850 ( .A(n406), .B(n407), .S0(n690), .Y(blockdata[113]) );
  MXI4XL U851 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n738), .S1(n707), .Y(n407) );
  MXI4XL U852 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n738), .S1(n707), .Y(n406) );
  MXI2XL U853 ( .A(n634), .B(n635), .S0(n689), .Y(blockdata[17]) );
  MXI4XL U854 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n751), .S1(n725), .Y(n635) );
  MXI4XL U855 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n751), .S1(n725), .Y(n634) );
  MXI2XL U856 ( .A(n404), .B(n405), .S0(n690), .Y(blockdata[114]) );
  MXI4XL U857 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n738), .S1(n719), .Y(n405) );
  MXI4XL U858 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n738), .S1(n707), .Y(n404) );
  MXI2XL U859 ( .A(n632), .B(n633), .S0(n695), .Y(blockdata[18]) );
  MXI4XL U860 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n750), .S1(n725), .Y(n633) );
  MXI4XL U861 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n751), .S1(n725), .Y(n632) );
  MXI2XL U862 ( .A(n402), .B(n403), .S0(n690), .Y(blockdata[115]) );
  MXI4XL U863 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n738), .S1(n706), .Y(n403) );
  MXI4XL U864 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n738), .S1(n719), .Y(n402) );
  MXI2XL U865 ( .A(n630), .B(n631), .S0(n694), .Y(blockdata[19]) );
  MXI4XL U866 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n750), .S1(n725), .Y(n631) );
  MXI4XL U867 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n750), .S1(n725), .Y(n630) );
  MXI2XL U868 ( .A(n400), .B(n401), .S0(n690), .Y(blockdata[116]) );
  MXI4XL U869 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n737), .S1(n711), .Y(n401) );
  MXI4XL U870 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n737), .S1(n707), .Y(n400) );
  MXI2XL U871 ( .A(n628), .B(n629), .S0(n694), .Y(blockdata[20]) );
  MXI4XL U872 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n750), .S1(n725), .Y(n629) );
  MXI4XL U873 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n750), .S1(n725), .Y(n628) );
  MXI2XL U874 ( .A(n626), .B(n627), .S0(n696), .Y(blockdata[21]) );
  MXI4XL U875 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n750), .S1(n724), .Y(n627) );
  MXI4XL U876 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n750), .S1(n724), .Y(n626) );
  MXI2XL U877 ( .A(n624), .B(n625), .S0(n696), .Y(blockdata[22]) );
  MXI4XL U878 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n750), .S1(n724), .Y(n625) );
  MXI4XL U879 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n750), .S1(n724), .Y(n624) );
  MXI2XL U880 ( .A(n622), .B(n623), .S0(n696), .Y(blockdata[23]) );
  MXI4XL U881 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n750), .S1(n724), .Y(n623) );
  MXI4XL U882 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n750), .S1(n724), .Y(n622) );
  MXI2XL U883 ( .A(n620), .B(n621), .S0(n696), .Y(blockdata[24]) );
  MXI4XL U884 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n750), .S1(n724), .Y(n621) );
  MXI4XL U885 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n750), .S1(n724), .Y(n620) );
  MXI2XL U886 ( .A(n618), .B(n619), .S0(n696), .Y(blockdata[25]) );
  MXI4XL U887 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n749), .S1(n724), .Y(n619) );
  MXI4XL U888 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n749), .S1(n724), .Y(n618) );
  MXI2XL U889 ( .A(n398), .B(n399), .S0(n690), .Y(blockdata[117]) );
  MXI4XL U890 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n737), .S1(n710), .Y(n399) );
  MXI4XL U891 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n737), .S1(n710), .Y(n398) );
  MXI2XL U892 ( .A(n396), .B(n397), .S0(n690), .Y(blockdata[118]) );
  MXI4XL U893 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n737), .S1(n710), .Y(n397) );
  MXI4XL U894 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n737), .S1(n710), .Y(n396) );
  MXI2XL U895 ( .A(n394), .B(n395), .S0(n690), .Y(blockdata[119]) );
  MXI4XL U896 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n737), .S1(n710), .Y(n395) );
  MXI4XL U897 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n737), .S1(n710), .Y(n394) );
  MXI2XL U898 ( .A(n392), .B(n393), .S0(n690), .Y(blockdata[120]) );
  MXI4XL U899 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n737), .S1(n710), .Y(n393) );
  MXI4XL U900 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n737), .S1(n710), .Y(n392) );
  MXI2XL U901 ( .A(n390), .B(n391), .S0(n690), .Y(blockdata[121]) );
  MXI4XL U902 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n737), .S1(n710), .Y(n391) );
  MXI4XL U903 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n737), .S1(n710), .Y(n390) );
  NAND3BXL U904 ( .AN(proc_addr[0]), .B(n896), .C(n1112), .Y(n1063) );
  OR2X1 U905 ( .A(n2), .B(n1258), .Y(n301) );
  CLKBUFX3 U906 ( .A(n700), .Y(n718) );
  CLKBUFX3 U907 ( .A(n700), .Y(n714) );
  CLKBUFX3 U908 ( .A(n700), .Y(n723) );
  CLKBUFX3 U909 ( .A(n729), .Y(n717) );
  CLKBUFX3 U910 ( .A(n730), .Y(n713) );
  CLKBUFX3 U911 ( .A(n701), .Y(n724) );
  CLKBUFX3 U912 ( .A(n704), .Y(n721) );
  CLKBUFX3 U913 ( .A(n706), .Y(n716) );
  CLKBUFX3 U914 ( .A(n704), .Y(n722) );
  CLKBUFX3 U915 ( .A(n706), .Y(n715) );
  CLKBUFX3 U916 ( .A(n705), .Y(n720) );
  CLKBUFX3 U917 ( .A(n707), .Y(n711) );
  CLKBUFX3 U918 ( .A(n706), .Y(n712) );
  CLKBUFX3 U919 ( .A(n304), .Y(n841) );
  CLKBUFX3 U920 ( .A(n304), .Y(n842) );
  CLKBUFX3 U921 ( .A(n304), .Y(n843) );
  CLKBUFX3 U922 ( .A(n304), .Y(n844) );
  CLKBUFX3 U923 ( .A(n304), .Y(n845) );
  CLKBUFX3 U924 ( .A(n304), .Y(n846) );
  CLKBUFX3 U925 ( .A(n305), .Y(n808) );
  CLKBUFX3 U926 ( .A(n305), .Y(n809) );
  CLKBUFX3 U927 ( .A(n305), .Y(n810) );
  CLKBUFX3 U928 ( .A(n305), .Y(n811) );
  CLKBUFX3 U929 ( .A(n305), .Y(n812) );
  CLKBUFX3 U930 ( .A(n305), .Y(n813) );
  CLKBUFX3 U931 ( .A(n305), .Y(n814) );
  CLKBUFX3 U932 ( .A(n304), .Y(n839) );
  CLKBUFX3 U933 ( .A(n304), .Y(n840) );
  CLKBUFX3 U934 ( .A(n305), .Y(n807) );
  CLKBUFX3 U935 ( .A(n705), .Y(n719) );
  CLKBUFX3 U936 ( .A(n306), .Y(n825) );
  CLKBUFX3 U937 ( .A(n306), .Y(n826) );
  CLKBUFX3 U938 ( .A(n306), .Y(n827) );
  CLKBUFX3 U939 ( .A(n306), .Y(n828) );
  CLKBUFX3 U940 ( .A(n306), .Y(n829) );
  CLKBUFX3 U941 ( .A(n306), .Y(n830) );
  CLKBUFX3 U942 ( .A(n307), .Y(n792) );
  CLKBUFX3 U943 ( .A(n307), .Y(n793) );
  CLKBUFX3 U944 ( .A(n307), .Y(n794) );
  CLKBUFX3 U945 ( .A(n307), .Y(n795) );
  CLKBUFX3 U946 ( .A(n307), .Y(n796) );
  CLKBUFX3 U947 ( .A(n307), .Y(n797) );
  CLKBUFX3 U948 ( .A(n307), .Y(n798) );
  CLKBUFX3 U949 ( .A(n306), .Y(n823) );
  CLKBUFX3 U950 ( .A(n306), .Y(n824) );
  CLKBUFX3 U951 ( .A(n307), .Y(n791) );
  CLKBUFX3 U952 ( .A(n733), .Y(n737) );
  CLKBUFX3 U953 ( .A(n200), .Y(n748) );
  CLKBUFX3 U954 ( .A(n688), .Y(n691) );
  CLKBUFX3 U955 ( .A(n688), .Y(n696) );
  CLKBUFX3 U956 ( .A(n687), .Y(n693) );
  CLKBUFX3 U957 ( .A(n734), .Y(n744) );
  CLKBUFX3 U958 ( .A(n733), .Y(n746) );
  CLKBUFX3 U959 ( .A(n734), .Y(n742) );
  CLKBUFX3 U960 ( .A(n755), .Y(n740) );
  CLKBUFX3 U961 ( .A(n735), .Y(n738) );
  CLKBUFX3 U962 ( .A(n708), .Y(n710) );
  CLKBUFX3 U963 ( .A(n689), .Y(n695) );
  CLKBUFX3 U964 ( .A(n690), .Y(n692) );
  CLKBUFX3 U965 ( .A(n689), .Y(n694) );
  CLKBUFX3 U966 ( .A(n741), .Y(n750) );
  CLKBUFX3 U967 ( .A(n310), .Y(n849) );
  CLKBUFX3 U968 ( .A(n310), .Y(n850) );
  CLKBUFX3 U969 ( .A(n310), .Y(n851) );
  CLKBUFX3 U970 ( .A(n310), .Y(n852) );
  CLKBUFX3 U971 ( .A(n310), .Y(n853) );
  CLKBUFX3 U972 ( .A(n310), .Y(n854) );
  CLKBUFX3 U973 ( .A(n311), .Y(n817) );
  CLKBUFX3 U974 ( .A(n311), .Y(n818) );
  CLKBUFX3 U975 ( .A(n311), .Y(n819) );
  CLKBUFX3 U976 ( .A(n311), .Y(n820) );
  CLKBUFX3 U977 ( .A(n311), .Y(n821) );
  CLKBUFX3 U978 ( .A(n311), .Y(n822) );
  CLKBUFX3 U979 ( .A(n310), .Y(n847) );
  CLKBUFX3 U980 ( .A(n310), .Y(n848) );
  CLKBUFX3 U981 ( .A(n311), .Y(n815) );
  CLKBUFX3 U982 ( .A(n311), .Y(n816) );
  CLKBUFX3 U983 ( .A(n315), .Y(n833) );
  CLKBUFX3 U984 ( .A(n315), .Y(n834) );
  CLKBUFX3 U985 ( .A(n315), .Y(n835) );
  CLKBUFX3 U986 ( .A(n315), .Y(n836) );
  CLKBUFX3 U987 ( .A(n315), .Y(n837) );
  CLKBUFX3 U988 ( .A(n315), .Y(n838) );
  CLKBUFX3 U989 ( .A(n316), .Y(n801) );
  CLKBUFX3 U990 ( .A(n316), .Y(n802) );
  CLKBUFX3 U991 ( .A(n316), .Y(n803) );
  CLKBUFX3 U992 ( .A(n316), .Y(n804) );
  CLKBUFX3 U993 ( .A(n316), .Y(n805) );
  CLKBUFX3 U994 ( .A(n316), .Y(n806) );
  CLKBUFX3 U995 ( .A(n315), .Y(n831) );
  CLKBUFX3 U996 ( .A(n315), .Y(n832) );
  CLKBUFX3 U997 ( .A(n316), .Y(n799) );
  CLKBUFX3 U998 ( .A(n316), .Y(n800) );
  CLKBUFX6 U999 ( .A(n1315), .Y(mem_write) );
  CLKBUFX3 U1000 ( .A(n729), .Y(n701) );
  CLKBUFX3 U1001 ( .A(n730), .Y(n700) );
  CLKBUFX3 U1002 ( .A(n699), .Y(n708) );
  CLKBUFX3 U1003 ( .A(n729), .Y(n699) );
  CLKBUFX3 U1004 ( .A(n303), .Y(n770) );
  CLKBUFX3 U1005 ( .A(n319), .Y(n775) );
  CLKBUFX3 U1006 ( .A(n783), .Y(n776) );
  CLKBUFX3 U1007 ( .A(n783), .Y(n777) );
  CLKBUFX3 U1008 ( .A(n783), .Y(n778) );
  CLKBUFX3 U1009 ( .A(n319), .Y(n779) );
  CLKBUFX3 U1010 ( .A(n783), .Y(n780) );
  CLKBUFX3 U1011 ( .A(n783), .Y(n781) );
  CLKBUFX3 U1012 ( .A(n783), .Y(n782) );
  CLKBUFX3 U1013 ( .A(n733), .Y(n735) );
  AND2X2 U1014 ( .A(n308), .B(n998), .Y(n303) );
  CLKBUFX3 U1015 ( .A(n309), .Y(n766) );
  CLKBUFX3 U1016 ( .A(n309), .Y(n765) );
  CLKBUFX3 U1017 ( .A(n964), .Y(n761) );
  CLKINVX1 U1018 ( .A(n863), .Y(n866) );
  AND2X2 U1019 ( .A(n312), .B(n864), .Y(n304) );
  AND2X2 U1020 ( .A(n313), .B(n864), .Y(n305) );
  AND2X2 U1021 ( .A(n317), .B(n864), .Y(n306) );
  AND2X2 U1022 ( .A(n314), .B(n864), .Y(n307) );
  CLKBUFX3 U1023 ( .A(n865), .Y(n864) );
  CLKBUFX3 U1024 ( .A(n929), .Y(n760) );
  CLKBUFX3 U1025 ( .A(n929), .Y(n759) );
  CLKBUFX3 U1026 ( .A(n965), .Y(n763) );
  CLKBUFX3 U1027 ( .A(n965), .Y(n764) );
  OAI221X1 U1028 ( .A0(n5), .A1(n1173), .B0(n790), .B1(n1172), .C0(n1171), .Y(
        proc_rdata[11]) );
  OA22X1 U1029 ( .A0(n788), .A1(n1170), .B0(n7), .B1(n1169), .Y(n1171) );
  OAI221X1 U1030 ( .A0(n5), .A1(n1188), .B0(n790), .B1(n1187), .C0(n1186), .Y(
        proc_rdata[14]) );
  OA22X1 U1031 ( .A0(n789), .A1(n1185), .B0(n7), .B1(n1184), .Y(n1186) );
  OAI221X1 U1032 ( .A0(n6), .A1(n1183), .B0(n790), .B1(n1182), .C0(n1181), .Y(
        proc_rdata[13]) );
  OA22X1 U1033 ( .A0(n789), .A1(n1180), .B0(n7), .B1(n1179), .Y(n1181) );
  OAI221X1 U1034 ( .A0(n5), .A1(n1168), .B0(n790), .B1(n1167), .C0(n1166), .Y(
        proc_rdata[10]) );
  OA22X1 U1035 ( .A0(n788), .A1(n1165), .B0(n8), .B1(n1164), .Y(n1166) );
  OAI221X1 U1036 ( .A0(n6), .A1(n1158), .B0(n790), .B1(n1157), .C0(n1156), .Y(
        proc_rdata[8]) );
  OA22X1 U1037 ( .A0(n788), .A1(n1155), .B0(n7), .B1(n1154), .Y(n1156) );
  OAI221X1 U1038 ( .A0(n5), .A1(n1148), .B0(n790), .B1(n1147), .C0(n1146), .Y(
        proc_rdata[6]) );
  OA22X1 U1039 ( .A0(n788), .A1(n1145), .B0(n8), .B1(n1144), .Y(n1146) );
  OAI221X1 U1040 ( .A0(n5), .A1(n1193), .B0(n790), .B1(n1192), .C0(n1191), .Y(
        proc_rdata[15]) );
  OAI221X1 U1041 ( .A0(n6), .A1(n1178), .B0(n790), .B1(n1177), .C0(n1176), .Y(
        proc_rdata[12]) );
  OA22X1 U1042 ( .A0(n789), .A1(n1175), .B0(n7), .B1(n1174), .Y(n1176) );
  OAI221X1 U1043 ( .A0(n5), .A1(n1123), .B0(n790), .B1(n1122), .C0(n1121), .Y(
        proc_rdata[1]) );
  OAI221X1 U1044 ( .A0(n6), .A1(n1153), .B0(n790), .B1(n1152), .C0(n1151), .Y(
        proc_rdata[7]) );
  OAI221X1 U1045 ( .A0(n6), .A1(n1133), .B0(n790), .B1(n1132), .C0(n1131), .Y(
        proc_rdata[3]) );
  OAI221X1 U1046 ( .A0(n5), .A1(n1143), .B0(n790), .B1(n1142), .C0(n1141), .Y(
        proc_rdata[5]) );
  OA22X1 U1047 ( .A0(n788), .A1(n1140), .B0(n8), .B1(n1139), .Y(n1141) );
  OAI221X1 U1048 ( .A0(n5), .A1(n1138), .B0(n790), .B1(n1137), .C0(n1136), .Y(
        proc_rdata[4]) );
  OAI221X1 U1049 ( .A0(n5), .A1(n1128), .B0(n790), .B1(n1127), .C0(n1126), .Y(
        proc_rdata[2]) );
  OA22X1 U1050 ( .A0(n788), .A1(n1125), .B0(n8), .B1(n1124), .Y(n1126) );
  OAI221X1 U1051 ( .A0(n5), .A1(n1118), .B0(n790), .B1(n1117), .C0(n1116), .Y(
        proc_rdata[0]) );
  CLKINVX1 U1052 ( .A(n1106), .Y(n1315) );
  AND2X2 U1053 ( .A(n308), .B(n774), .Y(n309) );
  CLKBUFX3 U1054 ( .A(n105), .Y(n758) );
  CLKBUFX3 U1055 ( .A(n105), .Y(n757) );
  OAI221XL U1056 ( .A0(n6), .A1(n1198), .B0(n790), .B1(n1197), .C0(n1196), .Y(
        proc_rdata[16]) );
  OAI221XL U1057 ( .A0(n6), .A1(n1203), .B0(n790), .B1(n1202), .C0(n1201), .Y(
        proc_rdata[17]) );
  OAI221XL U1058 ( .A0(n5), .A1(n1208), .B0(n790), .B1(n1207), .C0(n1206), .Y(
        proc_rdata[18]) );
  OAI221XL U1059 ( .A0(n5), .A1(n1213), .B0(n790), .B1(n1212), .C0(n1211), .Y(
        proc_rdata[19]) );
  OAI221XL U1060 ( .A0(n5), .A1(n1218), .B0(n790), .B1(n1217), .C0(n1216), .Y(
        proc_rdata[20]) );
  OAI221XL U1061 ( .A0(n5), .A1(n1223), .B0(n790), .B1(n1222), .C0(n1221), .Y(
        proc_rdata[21]) );
  OAI221XL U1062 ( .A0(n6), .A1(n1228), .B0(n790), .B1(n1227), .C0(n1226), .Y(
        proc_rdata[22]) );
  OAI221XL U1063 ( .A0(n5), .A1(n1233), .B0(n790), .B1(n1232), .C0(n1231), .Y(
        proc_rdata[23]) );
  CLKBUFX3 U1064 ( .A(n787), .Y(n788) );
  CLKBUFX3 U1065 ( .A(n787), .Y(n789) );
  AND2X2 U1066 ( .A(n321), .B(n864), .Y(n310) );
  AND2X2 U1067 ( .A(n322), .B(n864), .Y(n311) );
  AND2X2 U1068 ( .A(n1310), .B(N31), .Y(n312) );
  AND2X2 U1069 ( .A(n1312), .B(N31), .Y(n313) );
  AND2X2 U1070 ( .A(n1313), .B(N31), .Y(n314) );
  AND2X2 U1071 ( .A(n323), .B(n864), .Y(n315) );
  AND2X2 U1072 ( .A(n324), .B(n864), .Y(n316) );
  AND2X2 U1073 ( .A(n1311), .B(N31), .Y(n317) );
  CLKBUFX3 U1074 ( .A(n1063), .Y(n772) );
  CLKBUFX3 U1075 ( .A(n1063), .Y(n773) );
  INVX3 U1076 ( .A(n769), .Y(n767) );
  INVX3 U1077 ( .A(n769), .Y(n768) );
  NAND2X1 U1078 ( .A(dirty), .B(valid), .Y(n1105) );
  CLKINVX1 U1079 ( .A(blockdata[124]), .Y(n1257) );
  CLKINVX1 U1080 ( .A(blockdata[28]), .Y(n1258) );
  CLKINVX1 U1081 ( .A(blockdata[122]), .Y(n1247) );
  CLKINVX1 U1082 ( .A(blockdata[60]), .Y(n1254) );
  CLKINVX1 U1083 ( .A(blockdata[58]), .Y(n1244) );
  CLKINVX1 U1084 ( .A(blockdata[92]), .Y(n1255) );
  CLKINVX1 U1085 ( .A(blockdata[90]), .Y(n1245) );
  CLKINVX1 U1086 ( .A(n1107), .Y(n1314) );
  CLKINVX1 U1087 ( .A(blockdata[26]), .Y(n1248) );
  CLKINVX1 U1088 ( .A(blockdata[104]), .Y(n1157) );
  CLKINVX1 U1089 ( .A(blockdata[8]), .Y(n1158) );
  CLKINVX1 U1090 ( .A(blockdata[103]), .Y(n1152) );
  CLKINVX1 U1091 ( .A(blockdata[7]), .Y(n1153) );
  CLKINVX1 U1092 ( .A(blockdata[102]), .Y(n1147) );
  CLKINVX1 U1093 ( .A(blockdata[6]), .Y(n1148) );
  CLKINVX1 U1094 ( .A(blockdata[101]), .Y(n1142) );
  CLKINVX1 U1095 ( .A(blockdata[100]), .Y(n1137) );
  CLKINVX1 U1096 ( .A(blockdata[4]), .Y(n1138) );
  CLKINVX1 U1097 ( .A(blockdata[98]), .Y(n1127) );
  CLKINVX1 U1098 ( .A(blockdata[2]), .Y(n1128) );
  CLKINVX1 U1099 ( .A(blockdata[96]), .Y(n1117) );
  CLKINVX1 U1100 ( .A(blockdata[0]), .Y(n1118) );
  CLKINVX1 U1101 ( .A(blockdata[97]), .Y(n1122) );
  CLKINVX1 U1102 ( .A(blockdata[1]), .Y(n1123) );
  CLKINVX1 U1103 ( .A(blockdata[99]), .Y(n1132) );
  CLKINVX1 U1104 ( .A(blockdata[3]), .Y(n1133) );
  CLKINVX1 U1105 ( .A(blockdata[32]), .Y(n1114) );
  CLKINVX1 U1106 ( .A(blockdata[68]), .Y(n1135) );
  CLKINVX1 U1107 ( .A(blockdata[66]), .Y(n1125) );
  CLKINVX1 U1108 ( .A(blockdata[64]), .Y(n1115) );
  CLKINVX1 U1109 ( .A(blockdata[65]), .Y(n1120) );
  CLKINVX1 U1110 ( .A(blockdata[67]), .Y(n1130) );
  AND2X2 U1111 ( .A(n930), .B(n929), .Y(n320) );
  AND2X2 U1112 ( .A(n1066), .B(n1065), .Y(n1101) );
  OAI21XL U1113 ( .A0(n1102), .A1(n1064), .B0(dirty), .Y(n1066) );
  CLKINVX1 U1114 ( .A(blockdata[112]), .Y(n1197) );
  CLKINVX1 U1115 ( .A(blockdata[16]), .Y(n1198) );
  CLKINVX1 U1116 ( .A(blockdata[113]), .Y(n1202) );
  CLKINVX1 U1117 ( .A(blockdata[17]), .Y(n1203) );
  CLKINVX1 U1118 ( .A(blockdata[114]), .Y(n1207) );
  CLKINVX1 U1119 ( .A(blockdata[18]), .Y(n1208) );
  CLKINVX1 U1120 ( .A(blockdata[115]), .Y(n1212) );
  CLKINVX1 U1121 ( .A(blockdata[19]), .Y(n1213) );
  CLKINVX1 U1122 ( .A(blockdata[116]), .Y(n1217) );
  CLKINVX1 U1123 ( .A(blockdata[20]), .Y(n1218) );
  CLKINVX1 U1124 ( .A(blockdata[117]), .Y(n1222) );
  CLKINVX1 U1125 ( .A(blockdata[21]), .Y(n1223) );
  CLKINVX1 U1126 ( .A(blockdata[118]), .Y(n1227) );
  CLKINVX1 U1127 ( .A(blockdata[22]), .Y(n1228) );
  CLKINVX1 U1128 ( .A(blockdata[119]), .Y(n1232) );
  CLKINVX1 U1129 ( .A(blockdata[23]), .Y(n1233) );
  CLKINVX1 U1130 ( .A(blockdata[120]), .Y(n1237) );
  CLKINVX1 U1131 ( .A(blockdata[24]), .Y(n1238) );
  CLKINVX1 U1132 ( .A(blockdata[121]), .Y(n1242) );
  CLKINVX1 U1133 ( .A(blockdata[25]), .Y(n1243) );
  CLKINVX1 U1134 ( .A(blockdata[48]), .Y(n1194) );
  CLKINVX1 U1135 ( .A(blockdata[49]), .Y(n1199) );
  CLKINVX1 U1136 ( .A(blockdata[50]), .Y(n1204) );
  CLKINVX1 U1137 ( .A(blockdata[51]), .Y(n1209) );
  CLKINVX1 U1138 ( .A(blockdata[52]), .Y(n1214) );
  CLKINVX1 U1139 ( .A(blockdata[53]), .Y(n1219) );
  CLKINVX1 U1140 ( .A(blockdata[54]), .Y(n1224) );
  CLKINVX1 U1141 ( .A(blockdata[55]), .Y(n1229) );
  CLKINVX1 U1142 ( .A(blockdata[56]), .Y(n1234) );
  CLKINVX1 U1143 ( .A(blockdata[57]), .Y(n1239) );
  CLKINVX1 U1144 ( .A(blockdata[80]), .Y(n1195) );
  CLKINVX1 U1145 ( .A(blockdata[81]), .Y(n1200) );
  CLKINVX1 U1146 ( .A(blockdata[82]), .Y(n1205) );
  CLKINVX1 U1147 ( .A(blockdata[83]), .Y(n1210) );
  CLKINVX1 U1148 ( .A(blockdata[84]), .Y(n1215) );
  CLKINVX1 U1149 ( .A(blockdata[85]), .Y(n1220) );
  CLKINVX1 U1150 ( .A(blockdata[86]), .Y(n1225) );
  CLKINVX1 U1151 ( .A(blockdata[87]), .Y(n1230) );
  CLKINVX1 U1152 ( .A(blockdata[88]), .Y(n1235) );
  CLKINVX1 U1153 ( .A(blockdata[89]), .Y(n1240) );
  NAND3BX1 U1154 ( .AN(n1112), .B(n896), .C(n1111), .Y(n965) );
  CLKINVX1 U1155 ( .A(n1065), .Y(n896) );
  NAND2X1 U1156 ( .A(n896), .B(n376), .Y(n929) );
  CLKINVX1 U1157 ( .A(n998), .Y(n769) );
  NAND3BX1 U1158 ( .AN(n1111), .B(n896), .C(n1112), .Y(n998) );
  CLKBUFX3 U1159 ( .A(n1063), .Y(n774) );
  MX4X1 U1160 ( .A(\blocktag[0][19] ), .B(\blocktag[1][19] ), .C(
        \blocktag[2][19] ), .D(\blocktag[3][19] ), .S0(n199), .S1(n703), .Y(
        n347) );
  MXI2X1 U1161 ( .A(n542), .B(n543), .S0(n693), .Y(blockdata[63]) );
  MXI2X1 U1162 ( .A(n442), .B(n443), .S0(n691), .Y(blockdata[95]) );
  MXI2X1 U1163 ( .A(n546), .B(n547), .S0(n693), .Y(blockdata[61]) );
  MXI4X1 U1164 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n745), .S1(n718), .Y(n546) );
  MXI4X1 U1165 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n745), .S1(n718), .Y(n547) );
  MXI2X1 U1166 ( .A(n446), .B(n447), .S0(n690), .Y(blockdata[93]) );
  MXI2X1 U1167 ( .A(n544), .B(n545), .S0(n693), .Y(blockdata[62]) );
  MXI4X1 U1168 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n745), .S1(n718), .Y(n544) );
  MXI4X1 U1169 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n745), .S1(n718), .Y(n545) );
  MXI2X1 U1170 ( .A(n444), .B(n445), .S0(n693), .Y(blockdata[94]) );
  MXI4X1 U1171 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n745), .S1(n718), .Y(n548) );
  MXI4X1 U1172 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n741), .S1(n714), .Y(n448) );
  MXI4X1 U1173 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n741), .S1(n714), .Y(n449) );
  MXI2X1 U1174 ( .A(n378), .B(n379), .S0(n690), .Y(blockdata[127]) );
  MXI2X1 U1175 ( .A(n606), .B(n607), .S0(n696), .Y(blockdata[31]) );
  MXI4X1 U1176 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n749), .S1(n723), .Y(n606) );
  MXI4X1 U1177 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n748), .S1(n723), .Y(n607) );
  MXI2X1 U1178 ( .A(n382), .B(n383), .S0(n690), .Y(blockdata[125]) );
  MXI2X1 U1179 ( .A(n610), .B(n611), .S0(n696), .Y(blockdata[29]) );
  MXI4X1 U1180 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n749), .S1(n723), .Y(n610) );
  MXI4X1 U1181 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n749), .S1(n723), .Y(n611) );
  MXI2X1 U1182 ( .A(n380), .B(n381), .S0(n690), .Y(blockdata[126]) );
  MXI2X1 U1183 ( .A(n608), .B(n609), .S0(n696), .Y(blockdata[30]) );
  MXI4X1 U1184 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n736), .S1(n709), .Y(n384) );
  MXI4X1 U1185 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n749), .S1(n723), .Y(n612) );
  MXI2X1 U1186 ( .A(n550), .B(n551), .S0(n693), .Y(blockdata[59]) );
  MXI4X1 U1187 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n745), .S1(n718), .Y(n550) );
  MXI4X1 U1188 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n745), .S1(n718), .Y(n551) );
  MXI2X1 U1189 ( .A(n450), .B(n451), .S0(n691), .Y(blockdata[91]) );
  MXI4X1 U1190 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n741), .S1(n714), .Y(n450) );
  MXI4X1 U1191 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n741), .S1(n714), .Y(n451) );
  MXI2X1 U1192 ( .A(n386), .B(n387), .S0(n690), .Y(blockdata[123]) );
  MXI2X1 U1193 ( .A(n614), .B(n615), .S0(n696), .Y(blockdata[27]) );
  NAND2X1 U1194 ( .A(mem_rdata[1]), .B(n776), .Y(n1059) );
  NAND2X1 U1195 ( .A(mem_rdata[2]), .B(n776), .Y(n1057) );
  NAND2X1 U1196 ( .A(mem_rdata[3]), .B(n776), .Y(n1055) );
  NAND2X1 U1197 ( .A(mem_rdata[4]), .B(n776), .Y(n1053) );
  NAND2X1 U1198 ( .A(mem_rdata[5]), .B(n776), .Y(n1051) );
  NAND2X1 U1199 ( .A(mem_rdata[6]), .B(n776), .Y(n1049) );
  NAND2X1 U1200 ( .A(mem_rdata[7]), .B(n776), .Y(n1047) );
  NAND2X1 U1201 ( .A(mem_rdata[8]), .B(n776), .Y(n1045) );
  NAND2X1 U1202 ( .A(mem_rdata[9]), .B(n776), .Y(n1043) );
  NAND2X1 U1203 ( .A(mem_rdata[10]), .B(n776), .Y(n1041) );
  NAND2X1 U1204 ( .A(mem_rdata[11]), .B(n776), .Y(n1039) );
  NAND2X1 U1205 ( .A(mem_rdata[12]), .B(n776), .Y(n1037) );
  NAND2X1 U1206 ( .A(mem_rdata[13]), .B(n776), .Y(n1035) );
  NAND2X1 U1207 ( .A(mem_rdata[14]), .B(n777), .Y(n1033) );
  NAND2X1 U1208 ( .A(mem_rdata[15]), .B(n777), .Y(n1031) );
  NAND2X1 U1209 ( .A(mem_rdata[16]), .B(n777), .Y(n1029) );
  NAND2X1 U1210 ( .A(mem_rdata[17]), .B(n777), .Y(n1027) );
  NAND2X1 U1211 ( .A(mem_rdata[18]), .B(n777), .Y(n1025) );
  NAND2X1 U1212 ( .A(mem_rdata[19]), .B(n777), .Y(n1023) );
  NAND2X1 U1213 ( .A(mem_rdata[20]), .B(n777), .Y(n1021) );
  NAND2X1 U1214 ( .A(mem_rdata[21]), .B(n777), .Y(n1019) );
  NAND2X1 U1215 ( .A(mem_rdata[22]), .B(n777), .Y(n1017) );
  NAND2X1 U1216 ( .A(mem_rdata[23]), .B(n777), .Y(n1015) );
  NAND2X1 U1217 ( .A(mem_rdata[24]), .B(n777), .Y(n1013) );
  NAND2X1 U1218 ( .A(mem_rdata[25]), .B(n777), .Y(n1011) );
  NAND2X1 U1219 ( .A(mem_rdata[26]), .B(n777), .Y(n1009) );
  NAND2X1 U1220 ( .A(mem_rdata[27]), .B(n778), .Y(n1007) );
  NAND2X1 U1221 ( .A(mem_rdata[28]), .B(n778), .Y(n1005) );
  NAND2X1 U1222 ( .A(mem_rdata[29]), .B(n778), .Y(n1003) );
  NAND2X1 U1223 ( .A(mem_rdata[30]), .B(n778), .Y(n1001) );
  NAND2X1 U1224 ( .A(mem_rdata[31]), .B(n778), .Y(n999) );
  NAND2X1 U1225 ( .A(mem_rdata[32]), .B(n778), .Y(n997) );
  NAND2X1 U1226 ( .A(mem_rdata[33]), .B(n778), .Y(n996) );
  NAND2X1 U1227 ( .A(mem_rdata[34]), .B(n778), .Y(n995) );
  NAND2X1 U1228 ( .A(mem_rdata[35]), .B(n778), .Y(n994) );
  NAND2X1 U1229 ( .A(mem_rdata[36]), .B(n778), .Y(n993) );
  NAND2X1 U1230 ( .A(mem_rdata[37]), .B(n778), .Y(n992) );
  NAND2X1 U1231 ( .A(mem_rdata[38]), .B(n778), .Y(n991) );
  NAND2X1 U1232 ( .A(mem_rdata[39]), .B(n778), .Y(n990) );
  NAND2X1 U1233 ( .A(mem_rdata[40]), .B(n778), .Y(n989) );
  NAND2X1 U1234 ( .A(mem_rdata[41]), .B(n776), .Y(n988) );
  NAND2X1 U1235 ( .A(mem_rdata[42]), .B(n777), .Y(n987) );
  NAND2X1 U1236 ( .A(mem_rdata[43]), .B(n776), .Y(n986) );
  NAND2X1 U1237 ( .A(mem_rdata[44]), .B(n777), .Y(n985) );
  NAND2X1 U1238 ( .A(mem_rdata[45]), .B(n783), .Y(n984) );
  NAND2X1 U1239 ( .A(mem_rdata[46]), .B(n783), .Y(n983) );
  NAND2X1 U1240 ( .A(mem_rdata[47]), .B(n779), .Y(n982) );
  NAND2X1 U1241 ( .A(mem_rdata[48]), .B(n780), .Y(n981) );
  NAND2X1 U1242 ( .A(mem_rdata[49]), .B(n776), .Y(n980) );
  NAND2X1 U1243 ( .A(mem_rdata[50]), .B(n319), .Y(n979) );
  NAND2X1 U1244 ( .A(mem_rdata[51]), .B(n783), .Y(n978) );
  NAND2X1 U1245 ( .A(mem_rdata[52]), .B(n319), .Y(n977) );
  NAND2X1 U1246 ( .A(mem_rdata[53]), .B(n779), .Y(n976) );
  NAND2X1 U1247 ( .A(mem_rdata[54]), .B(n779), .Y(n975) );
  NAND2X1 U1248 ( .A(mem_rdata[55]), .B(n779), .Y(n974) );
  NAND2X1 U1249 ( .A(mem_rdata[56]), .B(n779), .Y(n973) );
  NAND2X1 U1250 ( .A(mem_rdata[57]), .B(n779), .Y(n972) );
  NAND2X1 U1251 ( .A(mem_rdata[58]), .B(n779), .Y(n971) );
  NAND2X1 U1252 ( .A(mem_rdata[59]), .B(n779), .Y(n970) );
  NAND2X1 U1253 ( .A(mem_rdata[60]), .B(n779), .Y(n969) );
  NAND2X1 U1254 ( .A(mem_rdata[61]), .B(n779), .Y(n968) );
  NAND2X1 U1255 ( .A(mem_rdata[62]), .B(n779), .Y(n967) );
  NAND2X1 U1256 ( .A(mem_rdata[63]), .B(n779), .Y(n966) );
  NAND2X1 U1257 ( .A(mem_rdata[64]), .B(n779), .Y(n963) );
  NAND2X1 U1258 ( .A(mem_rdata[65]), .B(n779), .Y(n962) );
  NAND2X1 U1259 ( .A(mem_rdata[66]), .B(n780), .Y(n961) );
  NAND2X1 U1260 ( .A(mem_rdata[67]), .B(n780), .Y(n960) );
  NAND2X1 U1261 ( .A(mem_rdata[68]), .B(n780), .Y(n959) );
  NAND2X1 U1262 ( .A(mem_rdata[69]), .B(n780), .Y(n958) );
  NAND2X1 U1263 ( .A(mem_rdata[70]), .B(n780), .Y(n957) );
  NAND2X1 U1264 ( .A(mem_rdata[71]), .B(n780), .Y(n956) );
  NAND2X1 U1265 ( .A(mem_rdata[72]), .B(n780), .Y(n955) );
  NAND2X1 U1266 ( .A(mem_rdata[73]), .B(n780), .Y(n954) );
  NAND2X1 U1267 ( .A(mem_rdata[74]), .B(n780), .Y(n953) );
  NAND2X1 U1268 ( .A(mem_rdata[75]), .B(n780), .Y(n952) );
  NAND2X1 U1269 ( .A(mem_rdata[76]), .B(n780), .Y(n951) );
  NAND2X1 U1270 ( .A(mem_rdata[77]), .B(n780), .Y(n950) );
  NAND2X1 U1271 ( .A(mem_rdata[78]), .B(n780), .Y(n949) );
  NAND2X1 U1272 ( .A(mem_rdata[79]), .B(n781), .Y(n948) );
  NAND2X1 U1273 ( .A(mem_rdata[80]), .B(n781), .Y(n947) );
  NAND2X1 U1274 ( .A(mem_rdata[81]), .B(n781), .Y(n946) );
  NAND2X1 U1275 ( .A(mem_rdata[82]), .B(n781), .Y(n945) );
  NAND2X1 U1276 ( .A(mem_rdata[83]), .B(n781), .Y(n944) );
  NAND2X1 U1277 ( .A(mem_rdata[84]), .B(n781), .Y(n943) );
  NAND2X1 U1278 ( .A(mem_rdata[85]), .B(n781), .Y(n942) );
  NAND2X1 U1279 ( .A(mem_rdata[86]), .B(n781), .Y(n941) );
  NAND2X1 U1280 ( .A(mem_rdata[87]), .B(n781), .Y(n940) );
  NAND2X1 U1281 ( .A(mem_rdata[88]), .B(n781), .Y(n939) );
  NAND2X1 U1282 ( .A(mem_rdata[89]), .B(n781), .Y(n938) );
  NAND2X1 U1283 ( .A(mem_rdata[90]), .B(n781), .Y(n937) );
  NAND2X1 U1284 ( .A(mem_rdata[91]), .B(n781), .Y(n936) );
  NAND2X1 U1285 ( .A(mem_rdata[92]), .B(n782), .Y(n935) );
  NAND2X1 U1286 ( .A(mem_rdata[93]), .B(n782), .Y(n934) );
  NAND2X1 U1287 ( .A(mem_rdata[94]), .B(n782), .Y(n933) );
  NAND2X1 U1288 ( .A(mem_rdata[95]), .B(n782), .Y(n932) );
  CLKINVX1 U1289 ( .A(proc_addr[19]), .Y(n1080) );
  CLKMX2X2 U1290 ( .A(tag[5]), .B(proc_addr[10]), .S0(n783), .Y(n374) );
  MXI2X1 U1291 ( .A(n510), .B(n511), .S0(n692), .Y(blockdata[79]) );
  MXI2X1 U1292 ( .A(n574), .B(n575), .S0(n694), .Y(blockdata[47]) );
  MXI4X1 U1293 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n746), .S1(n720), .Y(n574) );
  MXI2X1 U1294 ( .A(n512), .B(n513), .S0(n692), .Y(blockdata[78]) );
  MXI2X1 U1295 ( .A(n576), .B(n577), .S0(n694), .Y(blockdata[46]) );
  MXI2X1 U1296 ( .A(n514), .B(n515), .S0(n692), .Y(blockdata[77]) );
  MXI2X1 U1297 ( .A(n578), .B(n579), .S0(n694), .Y(blockdata[45]) );
  MXI2X1 U1298 ( .A(n516), .B(n517), .S0(n692), .Y(blockdata[76]) );
  MXI2X1 U1299 ( .A(n580), .B(n581), .S0(n695), .Y(blockdata[44]) );
  MXI2X1 U1300 ( .A(n518), .B(n519), .S0(n692), .Y(blockdata[75]) );
  MXI2X1 U1301 ( .A(n582), .B(n583), .S0(n695), .Y(blockdata[43]) );
  MXI2X1 U1302 ( .A(n520), .B(n521), .S0(n692), .Y(blockdata[74]) );
  MXI2X1 U1303 ( .A(n584), .B(n585), .S0(n695), .Y(blockdata[42]) );
  MXI2X1 U1304 ( .A(n522), .B(n523), .S0(n692), .Y(blockdata[73]) );
  MXI2X1 U1305 ( .A(n586), .B(n587), .S0(n695), .Y(blockdata[41]) );
  MXI2X1 U1306 ( .A(n524), .B(n525), .S0(n692), .Y(blockdata[72]) );
  MXI4X1 U1307 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n743), .S1(n716), .Y(n524) );
  MXI4X1 U1308 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n743), .S1(n716), .Y(n525) );
  MXI2X1 U1309 ( .A(n588), .B(n589), .S0(n695), .Y(blockdata[40]) );
  MXI4X1 U1310 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n747), .S1(n721), .Y(n588) );
  MXI4X1 U1311 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n747), .S1(n721), .Y(n589) );
  MXI2X1 U1312 ( .A(n526), .B(n527), .S0(n692), .Y(blockdata[71]) );
  MXI2X1 U1313 ( .A(n590), .B(n591), .S0(n695), .Y(blockdata[39]) );
  MXI2X1 U1314 ( .A(n528), .B(n529), .S0(n692), .Y(blockdata[70]) );
  MXI2X1 U1315 ( .A(n592), .B(n593), .S0(n695), .Y(blockdata[38]) );
  MXI2X1 U1316 ( .A(n530), .B(n531), .S0(n692), .Y(blockdata[69]) );
  MXI2X1 U1317 ( .A(n594), .B(n595), .S0(n695), .Y(blockdata[37]) );
  MXI2X1 U1318 ( .A(n596), .B(n597), .S0(n695), .Y(blockdata[36]) );
  MXI2X1 U1319 ( .A(n600), .B(n601), .S0(n695), .Y(blockdata[34]) );
  MXI2X1 U1320 ( .A(n602), .B(n603), .S0(n695), .Y(blockdata[33]) );
  MXI2X1 U1321 ( .A(n598), .B(n599), .S0(n695), .Y(blockdata[35]) );
  MXI4X1 U1322 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n738), .S1(n719), .Y(n567) );
  MXI4X1 U1323 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n735), .S1(n719), .Y(n566) );
  MXI4X1 U1324 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n735), .S1(n705), .Y(n502) );
  MXI4X1 U1325 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n742), .S1(n719), .Y(n565) );
  MXI4X1 U1326 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n739), .S1(n719), .Y(n564) );
  MXI4X1 U1327 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n747), .S1(n712), .Y(n465) );
  MXI4X1 U1328 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n747), .S1(n706), .Y(n464) );
  MXI4X1 U1329 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n739), .S1(n719), .Y(n563) );
  MXI4X1 U1330 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n739), .S1(n719), .Y(n562) );
  MXI4X1 U1331 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n751), .S1(n707), .Y(n463) );
  MXI4X1 U1332 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n751), .S1(n706), .Y(n462) );
  MXI4X1 U1333 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n752), .S1(n719), .Y(n561) );
  MXI4X1 U1334 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n742), .S1(n719), .Y(n560) );
  MXI4X1 U1335 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n739), .S1(n712), .Y(n461) );
  MXI4X1 U1336 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n738), .S1(n705), .Y(n460) );
  MXI4X1 U1337 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n750), .S1(n719), .Y(n559) );
  MXI4X1 U1338 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n740), .S1(n719), .Y(n558) );
  MXI4X1 U1339 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n742), .S1(n719), .Y(n557) );
  MXI4X1 U1340 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n752), .S1(n719), .Y(n556) );
  MXI2X1 U1341 ( .A(n410), .B(n411), .S0(n689), .Y(blockdata[111]) );
  MXI4X1 U1342 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n738), .S1(n719), .Y(n410) );
  MXI2X1 U1343 ( .A(n638), .B(n639), .S0(n692), .Y(blockdata[15]) );
  MXI4X1 U1344 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n751), .S1(n725), .Y(n638) );
  MXI4X1 U1345 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n751), .S1(n725), .Y(n639) );
  MXI2X1 U1346 ( .A(n412), .B(n413), .S0(n689), .Y(blockdata[110]) );
  MXI2X1 U1347 ( .A(n640), .B(n641), .S0(n692), .Y(blockdata[14]) );
  MXI2X1 U1348 ( .A(n414), .B(n415), .S0(n695), .Y(blockdata[109]) );
  MXI2X1 U1349 ( .A(n642), .B(n643), .S0(n692), .Y(blockdata[13]) );
  MXI2X1 U1350 ( .A(n416), .B(n417), .S0(n695), .Y(blockdata[108]) );
  MXI2X1 U1351 ( .A(n644), .B(n645), .S0(n692), .Y(blockdata[12]) );
  MXI2X1 U1352 ( .A(n418), .B(n419), .S0(n689), .Y(blockdata[107]) );
  MXI2X1 U1353 ( .A(n646), .B(n647), .S0(n692), .Y(blockdata[11]) );
  MXI2X1 U1354 ( .A(n420), .B(n421), .S0(n689), .Y(blockdata[106]) );
  MXI2X1 U1355 ( .A(n648), .B(n649), .S0(n694), .Y(blockdata[10]) );
  MXI2X1 U1356 ( .A(n422), .B(n423), .S0(n694), .Y(blockdata[105]) );
  MXI2X1 U1357 ( .A(n650), .B(n651), .S0(n694), .Y(blockdata[9]) );
  MXI4X1 U1358 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n747), .S1(n711), .Y(n650) );
  MXI4X1 U1359 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n739), .S1(n719), .Y(n651) );
  MXI4X1 U1360 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n739), .S1(n712), .Y(n424) );
  MXI4X1 U1361 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n739), .S1(n712), .Y(n425) );
  MXI4X1 U1362 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n747), .S1(n715), .Y(n652) );
  MXI4X1 U1363 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n747), .S1(n707), .Y(n653) );
  CLKINVX1 U1364 ( .A(mem_ready), .Y(n1102) );
  NAND2X1 U1365 ( .A(mem_rdata[96]), .B(n782), .Y(n928) );
  NAND2X1 U1366 ( .A(mem_rdata[97]), .B(n782), .Y(n927) );
  NAND2X1 U1367 ( .A(mem_rdata[98]), .B(n782), .Y(n926) );
  NAND2X1 U1368 ( .A(mem_rdata[99]), .B(n782), .Y(n925) );
  NAND2X1 U1369 ( .A(mem_rdata[100]), .B(n782), .Y(n924) );
  NAND2X1 U1370 ( .A(mem_rdata[101]), .B(n782), .Y(n923) );
  NAND2X1 U1371 ( .A(mem_rdata[102]), .B(n782), .Y(n922) );
  NAND2X1 U1372 ( .A(mem_rdata[103]), .B(n782), .Y(n921) );
  NAND2X1 U1373 ( .A(mem_rdata[104]), .B(n782), .Y(n920) );
  NAND2X1 U1374 ( .A(mem_rdata[105]), .B(n783), .Y(n919) );
  NAND2X1 U1375 ( .A(mem_rdata[106]), .B(n778), .Y(n918) );
  NAND2X1 U1376 ( .A(mem_rdata[107]), .B(n779), .Y(n917) );
  NAND2X1 U1377 ( .A(mem_rdata[108]), .B(n780), .Y(n916) );
  NAND2X1 U1378 ( .A(mem_rdata[109]), .B(n319), .Y(n915) );
  NAND2X1 U1379 ( .A(mem_rdata[110]), .B(n781), .Y(n914) );
  NAND2X1 U1380 ( .A(mem_rdata[111]), .B(n782), .Y(n913) );
  NAND2X1 U1381 ( .A(mem_rdata[112]), .B(n319), .Y(n912) );
  NAND2X1 U1382 ( .A(mem_rdata[113]), .B(n779), .Y(n911) );
  NAND2X1 U1383 ( .A(mem_rdata[114]), .B(n780), .Y(n910) );
  NAND2X1 U1384 ( .A(mem_rdata[115]), .B(n777), .Y(n909) );
  NAND2X1 U1385 ( .A(mem_rdata[116]), .B(n778), .Y(n908) );
  NAND2X1 U1386 ( .A(mem_rdata[117]), .B(n775), .Y(n907) );
  NAND2X1 U1387 ( .A(mem_rdata[118]), .B(n319), .Y(n906) );
  NAND2X1 U1388 ( .A(mem_rdata[119]), .B(n319), .Y(n905) );
  NAND2X1 U1389 ( .A(mem_rdata[120]), .B(n319), .Y(n904) );
  NAND2X1 U1390 ( .A(mem_rdata[121]), .B(n319), .Y(n903) );
  NAND2X1 U1391 ( .A(mem_rdata[122]), .B(n319), .Y(n902) );
  NAND2X1 U1392 ( .A(mem_rdata[123]), .B(n776), .Y(n901) );
  NAND2X1 U1393 ( .A(mem_rdata[124]), .B(n783), .Y(n900) );
  NAND2X1 U1394 ( .A(mem_rdata[125]), .B(n777), .Y(n899) );
  NAND2X1 U1395 ( .A(mem_rdata[126]), .B(n783), .Y(n898) );
  NAND2X1 U1396 ( .A(mem_rdata[127]), .B(n776), .Y(n897) );
  MXI2X1 U1397 ( .A(n1301), .B(n106), .S0(n321), .Y(n1285) );
  MXI2X1 U1398 ( .A(n1300), .B(n106), .S0(n312), .Y(n1284) );
  MXI2X1 U1399 ( .A(n1299), .B(n106), .S0(n323), .Y(n1283) );
  MXI2X1 U1400 ( .A(n1298), .B(n106), .S0(n317), .Y(n1282) );
  MXI2X1 U1401 ( .A(n1297), .B(n106), .S0(n322), .Y(n1281) );
  MXI2X1 U1402 ( .A(n1296), .B(n106), .S0(n313), .Y(n1280) );
  MXI2X1 U1403 ( .A(n1295), .B(n106), .S0(n324), .Y(n1279) );
  MXI2X1 U1404 ( .A(n1294), .B(n106), .S0(n314), .Y(n1278) );
  MXI2X1 U1405 ( .A(n1309), .B(n1101), .S0(n321), .Y(n1293) );
  MXI2X1 U1406 ( .A(n1308), .B(n1101), .S0(n312), .Y(n1292) );
  MXI2X1 U1407 ( .A(n1307), .B(n1101), .S0(n323), .Y(n1291) );
  MXI2X1 U1408 ( .A(n1306), .B(n1101), .S0(n317), .Y(n1290) );
  MXI2X1 U1409 ( .A(n1305), .B(n1101), .S0(n322), .Y(n1289) );
  MXI2X1 U1410 ( .A(n1304), .B(n1101), .S0(n313), .Y(n1288) );
  MXI2X1 U1411 ( .A(n1303), .B(n1101), .S0(n324), .Y(n1287) );
  MXI2X1 U1412 ( .A(n1302), .B(n1101), .S0(n314), .Y(n1286) );
  CLKINVX1 U1413 ( .A(proc_wdata[0]), .Y(n1062) );
  CLKINVX1 U1414 ( .A(proc_wdata[1]), .Y(n1060) );
  CLKINVX1 U1415 ( .A(proc_wdata[2]), .Y(n1058) );
  CLKINVX1 U1416 ( .A(proc_wdata[3]), .Y(n1056) );
  CLKINVX1 U1417 ( .A(proc_wdata[4]), .Y(n1054) );
  CLKINVX1 U1418 ( .A(proc_wdata[5]), .Y(n1052) );
  CLKINVX1 U1419 ( .A(proc_wdata[6]), .Y(n1050) );
  CLKINVX1 U1420 ( .A(proc_wdata[7]), .Y(n1048) );
  CLKINVX1 U1421 ( .A(proc_wdata[8]), .Y(n1046) );
  CLKINVX1 U1422 ( .A(proc_wdata[9]), .Y(n1044) );
  CLKINVX1 U1423 ( .A(proc_wdata[10]), .Y(n1042) );
  CLKINVX1 U1424 ( .A(proc_wdata[11]), .Y(n1040) );
  CLKINVX1 U1425 ( .A(proc_wdata[12]), .Y(n1038) );
  CLKINVX1 U1426 ( .A(proc_wdata[13]), .Y(n1036) );
  CLKINVX1 U1427 ( .A(proc_wdata[14]), .Y(n1034) );
  CLKINVX1 U1428 ( .A(proc_wdata[15]), .Y(n1032) );
  CLKINVX1 U1429 ( .A(proc_wdata[16]), .Y(n1030) );
  CLKINVX1 U1430 ( .A(proc_wdata[17]), .Y(n1028) );
  CLKINVX1 U1431 ( .A(proc_wdata[18]), .Y(n1026) );
  CLKINVX1 U1432 ( .A(proc_wdata[19]), .Y(n1024) );
  CLKINVX1 U1433 ( .A(proc_wdata[20]), .Y(n1022) );
  CLKINVX1 U1434 ( .A(proc_wdata[21]), .Y(n1020) );
  CLKINVX1 U1435 ( .A(proc_wdata[22]), .Y(n1018) );
  CLKINVX1 U1436 ( .A(proc_wdata[23]), .Y(n1016) );
  CLKINVX1 U1437 ( .A(proc_wdata[24]), .Y(n1014) );
  CLKINVX1 U1438 ( .A(proc_wdata[25]), .Y(n1012) );
  CLKINVX1 U1439 ( .A(proc_wdata[26]), .Y(n1010) );
  CLKINVX1 U1440 ( .A(proc_wdata[27]), .Y(n1008) );
  CLKINVX1 U1441 ( .A(proc_wdata[28]), .Y(n1006) );
  CLKINVX1 U1442 ( .A(proc_wdata[29]), .Y(n1004) );
  CLKINVX1 U1443 ( .A(proc_wdata[30]), .Y(n1002) );
  CLKINVX1 U1444 ( .A(proc_wdata[31]), .Y(n1000) );
  CLKINVX1 U1445 ( .A(proc_write), .Y(n1108) );
  MXI4XL U1446 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n752), .S1(n707), .Y(n670) );
  MXI4XL U1447 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n200), .S1(n701), .Y(n671) );
  MXI4X2 U1448 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n200), .S1(n726), .Y(
        n678) );
  NOR2XL U1449 ( .A(n857), .B(N32), .Y(n1312) );
  NOR2XL U1450 ( .A(N33), .B(N32), .Y(n1310) );
  NAND3BX4 U1451 ( .AN(proc_addr[0]), .B(n1110), .C(n1112), .Y(n1277) );
  NAND3BX4 U1452 ( .AN(n1113), .B(proc_addr[1]), .C(n1111), .Y(n1272) );
  NAND3BX4 U1453 ( .AN(n1113), .B(proc_addr[0]), .C(n1112), .Y(n1270) );
  NAND3BXL U1454 ( .AN(n1109), .B(proc_write), .C(n866), .Y(n1065) );
  OA22XL U1455 ( .A0(n1109), .A1(n866), .B0(n893), .B1(n377), .Y(n894) );
  OAI221X2 U1456 ( .A0(n757), .A1(n1274), .B0(n1000), .B1(n759), .C0(n897), 
        .Y(block_next[127]) );
  OAI221X2 U1457 ( .A0(n757), .A1(n1267), .B0(n1002), .B1(n759), .C0(n898), 
        .Y(block_next[126]) );
  OAI221X2 U1458 ( .A0(n757), .A1(n1262), .B0(n1004), .B1(n759), .C0(n899), 
        .Y(block_next[125]) );
  OAI221X2 U1459 ( .A0(n757), .A1(n1257), .B0(n1006), .B1(n759), .C0(n900), 
        .Y(block_next[124]) );
  OAI221X2 U1460 ( .A0(n757), .A1(n1252), .B0(n1008), .B1(n759), .C0(n901), 
        .Y(block_next[123]) );
  OAI221X2 U1461 ( .A0(n757), .A1(n1247), .B0(n1010), .B1(n759), .C0(n902), 
        .Y(block_next[122]) );
  OAI221X2 U1462 ( .A0(n757), .A1(n1242), .B0(n1012), .B1(n759), .C0(n903), 
        .Y(block_next[121]) );
  OAI221X2 U1463 ( .A0(n757), .A1(n1237), .B0(n1014), .B1(n759), .C0(n904), 
        .Y(block_next[120]) );
  OAI221X2 U1464 ( .A0(n757), .A1(n1232), .B0(n1016), .B1(n759), .C0(n905), 
        .Y(block_next[119]) );
  OAI221X2 U1465 ( .A0(n757), .A1(n1227), .B0(n1018), .B1(n759), .C0(n906), 
        .Y(block_next[118]) );
  OAI221X2 U1466 ( .A0(n757), .A1(n1222), .B0(n1020), .B1(n759), .C0(n907), 
        .Y(block_next[117]) );
  OAI221X2 U1467 ( .A0(n757), .A1(n1217), .B0(n1022), .B1(n759), .C0(n908), 
        .Y(block_next[116]) );
  OAI221X2 U1468 ( .A0(n758), .A1(n1212), .B0(n1024), .B1(n760), .C0(n909), 
        .Y(block_next[115]) );
  OAI221X2 U1469 ( .A0(n758), .A1(n1207), .B0(n1026), .B1(n760), .C0(n910), 
        .Y(block_next[114]) );
  OAI221X2 U1470 ( .A0(n758), .A1(n1202), .B0(n1028), .B1(n760), .C0(n911), 
        .Y(block_next[113]) );
  OAI221X2 U1471 ( .A0(n758), .A1(n1197), .B0(n1030), .B1(n760), .C0(n912), 
        .Y(block_next[112]) );
  OAI221X2 U1472 ( .A0(n758), .A1(n1192), .B0(n1032), .B1(n760), .C0(n913), 
        .Y(block_next[111]) );
  OAI221X2 U1473 ( .A0(n758), .A1(n1187), .B0(n1034), .B1(n760), .C0(n914), 
        .Y(block_next[110]) );
  OAI221X2 U1474 ( .A0(n758), .A1(n1182), .B0(n1036), .B1(n760), .C0(n915), 
        .Y(block_next[109]) );
  OAI221X2 U1475 ( .A0(n758), .A1(n1177), .B0(n1038), .B1(n760), .C0(n916), 
        .Y(block_next[108]) );
  OAI221X2 U1476 ( .A0(n758), .A1(n1172), .B0(n1040), .B1(n760), .C0(n917), 
        .Y(block_next[107]) );
  OAI221X2 U1477 ( .A0(n758), .A1(n1167), .B0(n1042), .B1(n760), .C0(n918), 
        .Y(block_next[106]) );
  OAI221X2 U1478 ( .A0(n758), .A1(n1162), .B0(n1044), .B1(n760), .C0(n919), 
        .Y(block_next[105]) );
  OAI221X2 U1479 ( .A0(n758), .A1(n1157), .B0(n1046), .B1(n760), .C0(n920), 
        .Y(block_next[104]) );
  OAI221X2 U1480 ( .A0(n105), .A1(n1152), .B0(n1048), .B1(n929), .C0(n921), 
        .Y(block_next[103]) );
  OAI221X2 U1481 ( .A0(n105), .A1(n1147), .B0(n1050), .B1(n929), .C0(n922), 
        .Y(block_next[102]) );
  OAI221X2 U1482 ( .A0(n757), .A1(n1142), .B0(n1052), .B1(n760), .C0(n923), 
        .Y(block_next[101]) );
  OAI221X2 U1483 ( .A0(n758), .A1(n1137), .B0(n1054), .B1(n759), .C0(n924), 
        .Y(block_next[100]) );
  OAI221X2 U1484 ( .A0(n757), .A1(n1132), .B0(n1056), .B1(n760), .C0(n925), 
        .Y(block_next[99]) );
  OAI221X2 U1485 ( .A0(n758), .A1(n1127), .B0(n1058), .B1(n759), .C0(n926), 
        .Y(block_next[98]) );
  OAI221X2 U1486 ( .A0(n757), .A1(n1122), .B0(n1060), .B1(n760), .C0(n927), 
        .Y(block_next[97]) );
  OAI221X2 U1487 ( .A0(n758), .A1(n1117), .B0(n1062), .B1(n759), .C0(n928), 
        .Y(block_next[96]) );
  CLKINVX3 U1488 ( .A(n931), .Y(n964) );
  OAI221X2 U1489 ( .A0(n761), .A1(n1271), .B0(n1000), .B1(n764), .C0(n932), 
        .Y(block_next[95]) );
  OAI221X2 U1490 ( .A0(n761), .A1(n1265), .B0(n1002), .B1(n763), .C0(n933), 
        .Y(block_next[94]) );
  OAI221X2 U1491 ( .A0(n761), .A1(n1260), .B0(n1004), .B1(n764), .C0(n934), 
        .Y(block_next[93]) );
  OAI221X2 U1492 ( .A0(n761), .A1(n1255), .B0(n1006), .B1(n763), .C0(n935), 
        .Y(block_next[92]) );
  OAI221X2 U1493 ( .A0(n761), .A1(n1250), .B0(n1008), .B1(n764), .C0(n936), 
        .Y(block_next[91]) );
  OAI221X2 U1494 ( .A0(n761), .A1(n1245), .B0(n1010), .B1(n763), .C0(n937), 
        .Y(block_next[90]) );
  OAI221X2 U1495 ( .A0(n761), .A1(n1240), .B0(n1012), .B1(n965), .C0(n938), 
        .Y(block_next[89]) );
  OAI221X2 U1496 ( .A0(n761), .A1(n1235), .B0(n1014), .B1(n965), .C0(n939), 
        .Y(block_next[88]) );
  OAI221X2 U1497 ( .A0(n761), .A1(n1230), .B0(n1016), .B1(n764), .C0(n940), 
        .Y(block_next[87]) );
  OAI221X2 U1498 ( .A0(n761), .A1(n1225), .B0(n1018), .B1(n764), .C0(n941), 
        .Y(block_next[86]) );
  OAI221X2 U1499 ( .A0(n761), .A1(n1220), .B0(n1020), .B1(n764), .C0(n942), 
        .Y(block_next[85]) );
  OAI221X2 U1500 ( .A0(n761), .A1(n1215), .B0(n1022), .B1(n764), .C0(n943), 
        .Y(block_next[84]) );
  OAI221X2 U1501 ( .A0(n964), .A1(n1210), .B0(n1024), .B1(n764), .C0(n944), 
        .Y(block_next[83]) );
  OAI221X2 U1502 ( .A0(n964), .A1(n1205), .B0(n1026), .B1(n764), .C0(n945), 
        .Y(block_next[82]) );
  OAI221X2 U1503 ( .A0(n964), .A1(n1200), .B0(n1028), .B1(n764), .C0(n946), 
        .Y(block_next[81]) );
  OAI221X2 U1504 ( .A0(n964), .A1(n1195), .B0(n1030), .B1(n764), .C0(n947), 
        .Y(block_next[80]) );
  OAI221X2 U1505 ( .A0(n964), .A1(n1190), .B0(n1032), .B1(n764), .C0(n948), 
        .Y(block_next[79]) );
  OAI221X2 U1506 ( .A0(n964), .A1(n1185), .B0(n1034), .B1(n764), .C0(n949), 
        .Y(block_next[78]) );
  OAI221X2 U1507 ( .A0(n964), .A1(n1180), .B0(n1036), .B1(n764), .C0(n950), 
        .Y(block_next[77]) );
  OAI221X2 U1508 ( .A0(n964), .A1(n1175), .B0(n1038), .B1(n763), .C0(n951), 
        .Y(block_next[76]) );
  OAI221X2 U1509 ( .A0(n964), .A1(n1170), .B0(n1040), .B1(n763), .C0(n952), 
        .Y(block_next[75]) );
  OAI221X2 U1510 ( .A0(n964), .A1(n1165), .B0(n1042), .B1(n763), .C0(n953), 
        .Y(block_next[74]) );
  OAI221X2 U1511 ( .A0(n964), .A1(n1160), .B0(n1044), .B1(n763), .C0(n954), 
        .Y(block_next[73]) );
  OAI221X2 U1512 ( .A0(n761), .A1(n1155), .B0(n1046), .B1(n763), .C0(n955), 
        .Y(block_next[72]) );
  OAI221X2 U1513 ( .A0(n762), .A1(n1150), .B0(n1048), .B1(n764), .C0(n956), 
        .Y(block_next[71]) );
  OAI221X2 U1514 ( .A0(n762), .A1(n1145), .B0(n1050), .B1(n763), .C0(n957), 
        .Y(block_next[70]) );
  OAI221X2 U1515 ( .A0(n762), .A1(n1140), .B0(n1052), .B1(n763), .C0(n958), 
        .Y(block_next[69]) );
  OAI221X2 U1516 ( .A0(n762), .A1(n1135), .B0(n1054), .B1(n763), .C0(n959), 
        .Y(block_next[68]) );
  OAI221X2 U1517 ( .A0(n762), .A1(n1130), .B0(n1056), .B1(n763), .C0(n960), 
        .Y(block_next[67]) );
  OAI221X2 U1518 ( .A0(n762), .A1(n1125), .B0(n1058), .B1(n763), .C0(n961), 
        .Y(block_next[66]) );
  OAI221X2 U1519 ( .A0(n762), .A1(n1120), .B0(n1060), .B1(n763), .C0(n962), 
        .Y(block_next[65]) );
  OAI221X2 U1520 ( .A0(n762), .A1(n1115), .B0(n1062), .B1(n763), .C0(n963), 
        .Y(block_next[64]) );
  OAI221X2 U1521 ( .A0(n765), .A1(n1269), .B0(n1000), .B1(n768), .C0(n966), 
        .Y(block_next[63]) );
  OAI221X2 U1522 ( .A0(n765), .A1(n1264), .B0(n1002), .B1(n767), .C0(n967), 
        .Y(block_next[62]) );
  OAI221X2 U1523 ( .A0(n765), .A1(n1259), .B0(n1004), .B1(n768), .C0(n968), 
        .Y(block_next[61]) );
  OAI221X2 U1524 ( .A0(n765), .A1(n1254), .B0(n1006), .B1(n767), .C0(n969), 
        .Y(block_next[60]) );
  OAI221X2 U1525 ( .A0(n765), .A1(n1249), .B0(n1008), .B1(n768), .C0(n970), 
        .Y(block_next[59]) );
  OAI221X2 U1526 ( .A0(n765), .A1(n1244), .B0(n1010), .B1(n767), .C0(n971), 
        .Y(block_next[58]) );
  OAI221X2 U1527 ( .A0(n765), .A1(n1239), .B0(n1012), .B1(n998), .C0(n972), 
        .Y(block_next[57]) );
  OAI221X2 U1528 ( .A0(n765), .A1(n1234), .B0(n1014), .B1(n998), .C0(n973), 
        .Y(block_next[56]) );
  OAI221X2 U1529 ( .A0(n765), .A1(n1229), .B0(n1016), .B1(n768), .C0(n974), 
        .Y(block_next[55]) );
  OAI221X2 U1530 ( .A0(n765), .A1(n1224), .B0(n1018), .B1(n768), .C0(n975), 
        .Y(block_next[54]) );
  OAI221X2 U1531 ( .A0(n765), .A1(n1219), .B0(n1020), .B1(n768), .C0(n976), 
        .Y(block_next[53]) );
  OAI221X2 U1532 ( .A0(n765), .A1(n1214), .B0(n1022), .B1(n768), .C0(n977), 
        .Y(block_next[52]) );
  OAI221X2 U1533 ( .A0(n766), .A1(n1209), .B0(n1024), .B1(n768), .C0(n978), 
        .Y(block_next[51]) );
  OAI221X2 U1534 ( .A0(n766), .A1(n1204), .B0(n1026), .B1(n768), .C0(n979), 
        .Y(block_next[50]) );
  OAI221X2 U1535 ( .A0(n766), .A1(n1199), .B0(n1028), .B1(n768), .C0(n980), 
        .Y(block_next[49]) );
  OAI221X2 U1536 ( .A0(n766), .A1(n1194), .B0(n1030), .B1(n768), .C0(n981), 
        .Y(block_next[48]) );
  OAI221X2 U1537 ( .A0(n766), .A1(n1189), .B0(n1032), .B1(n768), .C0(n982), 
        .Y(block_next[47]) );
  OAI221X2 U1538 ( .A0(n766), .A1(n1184), .B0(n1034), .B1(n768), .C0(n983), 
        .Y(block_next[46]) );
  OAI221X2 U1539 ( .A0(n766), .A1(n1179), .B0(n1036), .B1(n768), .C0(n984), 
        .Y(block_next[45]) );
  OAI221X2 U1540 ( .A0(n766), .A1(n1174), .B0(n1038), .B1(n767), .C0(n985), 
        .Y(block_next[44]) );
  OAI221X2 U1541 ( .A0(n766), .A1(n1169), .B0(n1040), .B1(n767), .C0(n986), 
        .Y(block_next[43]) );
  OAI221X2 U1542 ( .A0(n766), .A1(n1164), .B0(n1042), .B1(n767), .C0(n987), 
        .Y(block_next[42]) );
  OAI221X2 U1543 ( .A0(n766), .A1(n1159), .B0(n1044), .B1(n767), .C0(n988), 
        .Y(block_next[41]) );
  OAI221X2 U1544 ( .A0(n766), .A1(n1154), .B0(n1046), .B1(n767), .C0(n989), 
        .Y(block_next[40]) );
  OAI221X2 U1545 ( .A0(n309), .A1(n1149), .B0(n1048), .B1(n768), .C0(n990), 
        .Y(block_next[39]) );
  OAI221X2 U1546 ( .A0(n309), .A1(n1144), .B0(n1050), .B1(n767), .C0(n991), 
        .Y(block_next[38]) );
  OAI221X2 U1547 ( .A0(n309), .A1(n1139), .B0(n1052), .B1(n767), .C0(n992), 
        .Y(block_next[37]) );
  OAI221X2 U1548 ( .A0(n309), .A1(n1134), .B0(n1054), .B1(n767), .C0(n993), 
        .Y(block_next[36]) );
  OAI221X2 U1549 ( .A0(n309), .A1(n1129), .B0(n1056), .B1(n767), .C0(n994), 
        .Y(block_next[35]) );
  OAI221X2 U1550 ( .A0(n309), .A1(n1124), .B0(n1058), .B1(n767), .C0(n995), 
        .Y(block_next[34]) );
  OAI221X2 U1551 ( .A0(n309), .A1(n1119), .B0(n1060), .B1(n767), .C0(n996), 
        .Y(block_next[33]) );
  OAI221X2 U1552 ( .A0(n309), .A1(n1114), .B0(n1062), .B1(n767), .C0(n997), 
        .Y(block_next[32]) );
  OAI221X2 U1553 ( .A0(n774), .A1(n1000), .B0(n770), .B1(n1276), .C0(n999), 
        .Y(block_next[31]) );
  OAI221X2 U1554 ( .A0(n774), .A1(n1002), .B0(n770), .B1(n1268), .C0(n1001), 
        .Y(block_next[30]) );
  OAI221X2 U1555 ( .A0(n774), .A1(n1004), .B0(n770), .B1(n1263), .C0(n1003), 
        .Y(block_next[29]) );
  OAI221X2 U1556 ( .A0(n774), .A1(n1006), .B0(n770), .B1(n1258), .C0(n1005), 
        .Y(block_next[28]) );
  OAI221X2 U1557 ( .A0(n774), .A1(n1008), .B0(n770), .B1(n1253), .C0(n1007), 
        .Y(block_next[27]) );
  OAI221X2 U1558 ( .A0(n774), .A1(n1010), .B0(n770), .B1(n1248), .C0(n1009), 
        .Y(block_next[26]) );
  OAI221X2 U1559 ( .A0(n774), .A1(n1012), .B0(n770), .B1(n1243), .C0(n1011), 
        .Y(block_next[25]) );
  OAI221X2 U1560 ( .A0(n773), .A1(n1014), .B0(n770), .B1(n1238), .C0(n1013), 
        .Y(block_next[24]) );
  OAI221X2 U1561 ( .A0(n773), .A1(n1016), .B0(n770), .B1(n1233), .C0(n1015), 
        .Y(block_next[23]) );
  OAI221X2 U1562 ( .A0(n773), .A1(n1018), .B0(n770), .B1(n1228), .C0(n1017), 
        .Y(block_next[22]) );
  OAI221X2 U1563 ( .A0(n773), .A1(n1020), .B0(n770), .B1(n1223), .C0(n1019), 
        .Y(block_next[21]) );
  OAI221X2 U1564 ( .A0(n773), .A1(n1022), .B0(n770), .B1(n1218), .C0(n1021), 
        .Y(block_next[20]) );
  OAI221X2 U1565 ( .A0(n773), .A1(n1024), .B0(n771), .B1(n1213), .C0(n1023), 
        .Y(block_next[19]) );
  OAI221X2 U1566 ( .A0(n773), .A1(n1026), .B0(n770), .B1(n1208), .C0(n1025), 
        .Y(block_next[18]) );
  OAI221X2 U1567 ( .A0(n773), .A1(n1028), .B0(n770), .B1(n1203), .C0(n1027), 
        .Y(block_next[17]) );
  OAI221X2 U1568 ( .A0(n773), .A1(n1030), .B0(n303), .B1(n1198), .C0(n1029), 
        .Y(block_next[16]) );
  OAI221X2 U1569 ( .A0(n773), .A1(n1032), .B0(n303), .B1(n1193), .C0(n1031), 
        .Y(block_next[15]) );
  OAI221X2 U1570 ( .A0(n773), .A1(n1034), .B0(n303), .B1(n1188), .C0(n1033), 
        .Y(block_next[14]) );
  OAI221X2 U1571 ( .A0(n773), .A1(n1036), .B0(n303), .B1(n1183), .C0(n1035), 
        .Y(block_next[13]) );
  OAI221X2 U1572 ( .A0(n772), .A1(n1038), .B0(n303), .B1(n1178), .C0(n1037), 
        .Y(block_next[12]) );
  OAI221X2 U1573 ( .A0(n772), .A1(n1040), .B0(n303), .B1(n1173), .C0(n1039), 
        .Y(block_next[11]) );
  OAI221X2 U1574 ( .A0(n772), .A1(n1042), .B0(n303), .B1(n1168), .C0(n1041), 
        .Y(block_next[10]) );
  OAI221X2 U1575 ( .A0(n772), .A1(n1044), .B0(n303), .B1(n1163), .C0(n1043), 
        .Y(block_next[9]) );
  OAI221X2 U1576 ( .A0(n772), .A1(n1046), .B0(n771), .B1(n1158), .C0(n1045), 
        .Y(block_next[8]) );
  OAI221X2 U1577 ( .A0(n772), .A1(n1048), .B0(n771), .B1(n1153), .C0(n1047), 
        .Y(block_next[7]) );
  OAI221X2 U1578 ( .A0(n772), .A1(n1050), .B0(n771), .B1(n1148), .C0(n1049), 
        .Y(block_next[6]) );
  OAI221X2 U1579 ( .A0(n772), .A1(n1052), .B0(n771), .B1(n1143), .C0(n1051), 
        .Y(block_next[5]) );
  OAI221X2 U1580 ( .A0(n772), .A1(n1054), .B0(n771), .B1(n1138), .C0(n1053), 
        .Y(block_next[4]) );
  OAI221X2 U1581 ( .A0(n772), .A1(n1056), .B0(n771), .B1(n1133), .C0(n1055), 
        .Y(block_next[3]) );
  OAI221X2 U1582 ( .A0(n772), .A1(n1058), .B0(n771), .B1(n1128), .C0(n1057), 
        .Y(block_next[2]) );
  OAI221X2 U1583 ( .A0(n772), .A1(n1060), .B0(n771), .B1(n1123), .C0(n1059), 
        .Y(block_next[1]) );
  OAI221X2 U1584 ( .A0(n773), .A1(n1062), .B0(n771), .B1(n1118), .C0(n1061), 
        .Y(block_next[0]) );
  CLKINVX3 U1585 ( .A(n1079), .Y(blocktag_next[15]) );
  CLKINVX3 U1586 ( .A(n1100), .Y(blocktag_next[0]) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, ICACHE_ren, ICACHE_stall,
         DCACHE_ren, DCACHE_stall, n18, n19, n20, n28, n29;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n28), .ICACHE_ren(ICACHE_ren), 
        .ICACHE_addr(ICACHE_addr), .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(
        ICACHE_rdata), .DCACHE_ren(DCACHE_ren), .DCACHE_wen(DCACHE_wen), 
        .DCACHE_addr({DCACHE_addr[29:23], n49, DCACHE_addr[21:5], n50, n51, 
        n52, DCACHE_addr[1:0]}), .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(
        DCACHE_stall), .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n29), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:4], n51, n52, 
        DCACHE_addr[1:0]}), .proc_wdata(DCACHE_wdata), .proc_stall(
        DCACHE_stall), .proc_rdata(DCACHE_rdata), .mem_read(n30), .mem_write(
        n31), .mem_addr(mem_addr_D), .mem_rdata(mem_rdata_D), .mem_wdata({n32, 
        mem_wdata_D[126:94], n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
        mem_wdata_D[83:15], n43, n44, n45, n46, mem_wdata_D[10:0]}), 
        .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n29), .proc_read(ICACHE_ren), 
        .proc_write(1'b0), .proc_addr({ICACHE_addr[29:5], n20, n19, n18, 
        ICACHE_addr[1:0]}), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(ICACHE_rdata), 
        .mem_read(n47), .mem_write(n48), .mem_addr(mem_addr_I), .mem_rdata(
        mem_rdata_I), .mem_wdata(mem_wdata_I), .mem_ready(mem_ready_I) );
  CLKBUFX20 U2 ( .A(n50), .Y(DCACHE_addr[4]) );
  CLKBUFX3 U3 ( .A(rst_n), .Y(n28) );
  BUFX16 U4 ( .A(ICACHE_addr[3]), .Y(n19) );
  BUFX4 U5 ( .A(ICACHE_addr[4]), .Y(n20) );
  BUFX12 U6 ( .A(n46), .Y(mem_wdata_D[11]) );
  BUFX12 U7 ( .A(n45), .Y(mem_wdata_D[12]) );
  BUFX12 U8 ( .A(n44), .Y(mem_wdata_D[13]) );
  BUFX12 U9 ( .A(n43), .Y(mem_wdata_D[14]) );
  BUFX12 U10 ( .A(n42), .Y(mem_wdata_D[84]) );
  BUFX12 U11 ( .A(n41), .Y(mem_wdata_D[85]) );
  BUFX12 U12 ( .A(n40), .Y(mem_wdata_D[86]) );
  BUFX12 U13 ( .A(n39), .Y(mem_wdata_D[87]) );
  BUFX12 U14 ( .A(n38), .Y(mem_wdata_D[88]) );
  BUFX12 U15 ( .A(n37), .Y(mem_wdata_D[89]) );
  BUFX12 U16 ( .A(n36), .Y(mem_wdata_D[90]) );
  BUFX12 U17 ( .A(n35), .Y(mem_wdata_D[91]) );
  BUFX12 U18 ( .A(n34), .Y(mem_wdata_D[92]) );
  BUFX12 U19 ( .A(n33), .Y(mem_wdata_D[93]) );
  INVXL U20 ( .A(n28), .Y(n29) );
  BUFX20 U21 ( .A(ICACHE_addr[2]), .Y(n18) );
  BUFX12 U22 ( .A(n32), .Y(mem_wdata_D[127]) );
  BUFX12 U23 ( .A(n52), .Y(DCACHE_addr[2]) );
  BUFX12 U24 ( .A(n51), .Y(DCACHE_addr[3]) );
  BUFX12 U25 ( .A(n31), .Y(mem_write_D) );
  BUFX12 U26 ( .A(n48), .Y(mem_write_I) );
  BUFX12 U27 ( .A(n30), .Y(mem_read_D) );
  BUFX12 U28 ( .A(n47), .Y(mem_read_I) );
  BUFX16 U29 ( .A(n49), .Y(DCACHE_addr[22]) );
endmodule

