
module cache ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N85, N86, N87, valid, mem_ready_r, dirty, proc_stall_next,
         mem_read_next, proc_write_r, \blocktag[7][24] , \blocktag[7][20] ,
         \blocktag[7][19] , \blocktag[7][18] , \blocktag[7][15] ,
         \blocktag[7][14] , \blocktag[7][13] , \blocktag[7][12] ,
         \blocktag[7][11] , \blocktag[7][10] , \blocktag[7][9] ,
         \blocktag[7][8] , \blocktag[7][5] , \blocktag[7][3] ,
         \blocktag[7][1] , \blocktag[7][0] , \blocktag[6][24] ,
         \blocktag[6][20] , \blocktag[6][19] , \blocktag[6][18] ,
         \blocktag[6][15] , \blocktag[6][14] , \blocktag[6][13] ,
         \blocktag[6][12] , \blocktag[6][11] , \blocktag[6][10] ,
         \blocktag[6][9] , \blocktag[6][8] , \blocktag[6][5] ,
         \blocktag[6][3] , \blocktag[6][1] , \blocktag[6][0] ,
         \blocktag[5][24] , \blocktag[5][20] , \blocktag[5][19] ,
         \blocktag[5][18] , \blocktag[5][15] , \blocktag[5][14] ,
         \blocktag[5][13] , \blocktag[5][12] , \blocktag[5][11] ,
         \blocktag[5][10] , \blocktag[5][9] , \blocktag[5][8] ,
         \blocktag[5][5] , \blocktag[5][3] , \blocktag[5][1] ,
         \blocktag[5][0] , \blocktag[4][24] , \blocktag[4][20] ,
         \blocktag[4][19] , \blocktag[4][18] , \blocktag[4][15] ,
         \blocktag[4][14] , \blocktag[4][13] , \blocktag[4][12] ,
         \blocktag[4][11] , \blocktag[4][10] , \blocktag[4][9] ,
         \blocktag[4][8] , \blocktag[4][5] , \blocktag[4][3] ,
         \blocktag[4][1] , \blocktag[4][0] , \blocktag[3][24] ,
         \blocktag[3][20] , \blocktag[3][19] , \blocktag[3][18] ,
         \blocktag[3][15] , \blocktag[3][14] , \blocktag[3][13] ,
         \blocktag[3][12] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][9] , \blocktag[3][8] , \blocktag[3][5] ,
         \blocktag[3][3] , \blocktag[3][1] , \blocktag[3][0] ,
         \blocktag[2][24] , \blocktag[2][20] , \blocktag[2][19] ,
         \blocktag[2][18] , \blocktag[2][15] , \blocktag[2][14] ,
         \blocktag[2][13] , \blocktag[2][12] , \blocktag[2][11] ,
         \blocktag[2][10] , \blocktag[2][9] , \blocktag[2][8] ,
         \blocktag[2][5] , \blocktag[2][3] , \blocktag[2][1] ,
         \blocktag[2][0] , \blocktag[1][24] , \blocktag[1][20] ,
         \blocktag[1][19] , \blocktag[1][18] , \blocktag[1][15] ,
         \blocktag[1][14] , \blocktag[1][13] , \blocktag[1][12] ,
         \blocktag[1][11] , \blocktag[1][10] , \blocktag[1][9] ,
         \blocktag[1][8] , \blocktag[1][5] , \blocktag[1][3] ,
         \blocktag[1][1] , \blocktag[1][0] , \blocktag[0][24] ,
         \blocktag[0][20] , \blocktag[0][19] , \blocktag[0][18] ,
         \blocktag[0][15] , \blocktag[0][14] , \blocktag[0][13] ,
         \blocktag[0][12] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][9] , \blocktag[0][8] , \blocktag[0][5] ,
         \blocktag[0][3] , \blocktag[0][1] , \blocktag[0][0] , \block[7][127] ,
         \block[7][126] , \block[7][125] , \block[7][124] , \block[7][123] ,
         \block[7][122] , \block[7][121] , \block[7][120] , \block[7][119] ,
         \block[7][118] , \block[7][117] , \block[7][116] , \block[7][115] ,
         \block[7][114] , \block[7][113] , \block[7][112] , \block[7][111] ,
         \block[7][110] , \block[7][109] , \block[7][108] , \block[7][107] ,
         \block[7][106] , \block[7][105] , \block[7][104] , \block[7][103] ,
         \block[7][102] , \block[7][101] , \block[7][100] , \block[7][99] ,
         \block[7][98] , \block[7][97] , \block[7][96] , \block[7][95] ,
         \block[7][94] , \block[7][93] , \block[7][92] , \block[7][91] ,
         \block[7][90] , \block[7][89] , \block[7][88] , \block[7][87] ,
         \block[7][86] , \block[7][85] , \block[7][84] , \block[7][83] ,
         \block[7][82] , \block[7][81] , \block[7][80] , \block[7][79] ,
         \block[7][78] , \block[7][77] , \block[7][76] , \block[7][75] ,
         \block[7][74] , \block[7][73] , \block[7][72] , \block[7][71] ,
         \block[7][70] , \block[7][69] , \block[7][68] , \block[7][67] ,
         \block[7][66] , \block[7][65] , \block[7][64] , \block[7][63] ,
         \block[7][62] , \block[7][61] , \block[7][60] , \block[7][59] ,
         \block[7][58] , \block[7][57] , \block[7][56] , \block[7][55] ,
         \block[7][54] , \block[7][53] , \block[7][52] , \block[7][51] ,
         \block[7][50] , \block[7][49] , \block[7][48] , \block[7][47] ,
         \block[7][46] , \block[7][45] , \block[7][44] , \block[7][43] ,
         \block[7][42] , \block[7][41] , \block[7][40] , \block[7][39] ,
         \block[7][38] , \block[7][37] , \block[7][36] , \block[7][35] ,
         \block[7][34] , \block[7][33] , \block[7][32] , \block[7][31] ,
         \block[7][30] , \block[7][29] , \block[7][28] , \block[7][27] ,
         \block[7][26] , \block[7][25] , \block[7][24] , \block[7][23] ,
         \block[7][22] , \block[7][21] , \block[7][20] , \block[7][19] ,
         \block[7][18] , \block[7][17] , \block[7][16] , \block[7][15] ,
         \block[7][14] , \block[7][13] , \block[7][12] , \block[7][11] ,
         \block[7][10] , \block[7][9] , \block[7][8] , \block[7][7] ,
         \block[7][6] , \block[7][5] , \block[7][4] , \block[7][3] ,
         \block[7][2] , \block[7][1] , \block[7][0] , \block[6][127] ,
         \block[6][126] , \block[6][125] , \block[6][124] , \block[6][123] ,
         \block[6][122] , \block[6][121] , \block[6][120] , \block[6][119] ,
         \block[6][118] , \block[6][117] , \block[6][116] , \block[6][115] ,
         \block[6][114] , \block[6][113] , \block[6][112] , \block[6][111] ,
         \block[6][110] , \block[6][109] , \block[6][108] , \block[6][107] ,
         \block[6][106] , \block[6][105] , \block[6][104] , \block[6][103] ,
         \block[6][102] , \block[6][101] , \block[6][100] , \block[6][99] ,
         \block[6][98] , \block[6][97] , \block[6][96] , \block[6][95] ,
         \block[6][94] , \block[6][93] , \block[6][92] , \block[6][91] ,
         \block[6][90] , \block[6][89] , \block[6][88] , \block[6][87] ,
         \block[6][86] , \block[6][85] , \block[6][84] , \block[6][83] ,
         \block[6][82] , \block[6][81] , \block[6][80] , \block[6][79] ,
         \block[6][78] , \block[6][77] , \block[6][76] , \block[6][75] ,
         \block[6][74] , \block[6][73] , \block[6][72] , \block[6][71] ,
         \block[6][70] , \block[6][69] , \block[6][68] , \block[6][67] ,
         \block[6][66] , \block[6][65] , \block[6][64] , \block[6][63] ,
         \block[6][62] , \block[6][61] , \block[6][60] , \block[6][59] ,
         \block[6][58] , \block[6][57] , \block[6][56] , \block[6][55] ,
         \block[6][54] , \block[6][53] , \block[6][52] , \block[6][51] ,
         \block[6][50] , \block[6][49] , \block[6][48] , \block[6][47] ,
         \block[6][46] , \block[6][45] , \block[6][44] , \block[6][43] ,
         \block[6][42] , \block[6][41] , \block[6][40] , \block[6][39] ,
         \block[6][38] , \block[6][37] , \block[6][36] , \block[6][35] ,
         \block[6][34] , \block[6][33] , \block[6][32] , \block[6][31] ,
         \block[6][30] , \block[6][29] , \block[6][28] , \block[6][27] ,
         \block[6][26] , \block[6][25] , \block[6][24] , \block[6][23] ,
         \block[6][22] , \block[6][21] , \block[6][20] , \block[6][19] ,
         \block[6][18] , \block[6][17] , \block[6][16] , \block[6][15] ,
         \block[6][14] , \block[6][13] , \block[6][12] , \block[6][11] ,
         \block[6][10] , \block[6][9] , \block[6][8] , \block[6][7] ,
         \block[6][6] , \block[6][5] , \block[6][4] , \block[6][3] ,
         \block[6][2] , \block[6][1] , \block[6][0] , \block[5][127] ,
         \block[5][126] , \block[5][125] , \block[5][124] , \block[5][123] ,
         \block[5][122] , \block[5][121] , \block[5][120] , \block[5][119] ,
         \block[5][118] , \block[5][117] , \block[5][116] , \block[5][115] ,
         \block[5][114] , \block[5][113] , \block[5][112] , \block[5][111] ,
         \block[5][110] , \block[5][109] , \block[5][108] , \block[5][107] ,
         \block[5][106] , \block[5][105] , \block[5][104] , \block[5][103] ,
         \block[5][102] , \block[5][101] , \block[5][100] , \block[5][99] ,
         \block[5][98] , \block[5][97] , \block[5][96] , \block[5][95] ,
         \block[5][94] , \block[5][93] , \block[5][92] , \block[5][91] ,
         \block[5][90] , \block[5][89] , \block[5][88] , \block[5][87] ,
         \block[5][86] , \block[5][85] , \block[5][84] , \block[5][83] ,
         \block[5][82] , \block[5][81] , \block[5][80] , \block[5][79] ,
         \block[5][78] , \block[5][77] , \block[5][76] , \block[5][75] ,
         \block[5][74] , \block[5][73] , \block[5][72] , \block[5][71] ,
         \block[5][70] , \block[5][69] , \block[5][68] , \block[5][67] ,
         \block[5][66] , \block[5][65] , \block[5][64] , \block[5][63] ,
         \block[5][62] , \block[5][61] , \block[5][60] , \block[5][59] ,
         \block[5][58] , \block[5][57] , \block[5][56] , \block[5][55] ,
         \block[5][54] , \block[5][53] , \block[5][52] , \block[5][51] ,
         \block[5][50] , \block[5][49] , \block[5][48] , \block[5][47] ,
         \block[5][46] , \block[5][45] , \block[5][44] , \block[5][43] ,
         \block[5][42] , \block[5][41] , \block[5][40] , \block[5][39] ,
         \block[5][38] , \block[5][37] , \block[5][36] , \block[5][35] ,
         \block[5][34] , \block[5][33] , \block[5][32] , \block[5][31] ,
         \block[5][30] , \block[5][29] , \block[5][28] , \block[5][27] ,
         \block[5][26] , \block[5][25] , \block[5][24] , \block[5][23] ,
         \block[5][22] , \block[5][21] , \block[5][20] , \block[5][19] ,
         \block[5][18] , \block[5][17] , \block[5][16] , \block[5][15] ,
         \block[5][14] , \block[5][13] , \block[5][12] , \block[5][11] ,
         \block[5][10] , \block[5][9] , \block[5][8] , \block[5][7] ,
         \block[5][6] , \block[5][5] , \block[5][4] , \block[5][3] ,
         \block[5][2] , \block[5][1] , \block[5][0] , \block[4][127] ,
         \block[4][126] , \block[4][125] , \block[4][124] , \block[4][123] ,
         \block[4][122] , \block[4][121] , \block[4][120] , \block[4][119] ,
         \block[4][118] , \block[4][117] , \block[4][116] , \block[4][115] ,
         \block[4][114] , \block[4][113] , \block[4][112] , \block[4][111] ,
         \block[4][110] , \block[4][109] , \block[4][108] , \block[4][107] ,
         \block[4][106] , \block[4][105] , \block[4][104] , \block[4][103] ,
         \block[4][102] , \block[4][101] , \block[4][100] , \block[4][99] ,
         \block[4][98] , \block[4][97] , \block[4][96] , \block[4][95] ,
         \block[4][94] , \block[4][93] , \block[4][92] , \block[4][91] ,
         \block[4][90] , \block[4][89] , \block[4][88] , \block[4][87] ,
         \block[4][86] , \block[4][85] , \block[4][84] , \block[4][83] ,
         \block[4][82] , \block[4][81] , \block[4][80] , \block[4][79] ,
         \block[4][78] , \block[4][77] , \block[4][76] , \block[4][75] ,
         \block[4][74] , \block[4][73] , \block[4][72] , \block[4][71] ,
         \block[4][70] , \block[4][69] , \block[4][68] , \block[4][67] ,
         \block[4][66] , \block[4][65] , \block[4][64] , \block[4][63] ,
         \block[4][62] , \block[4][61] , \block[4][60] , \block[4][59] ,
         \block[4][58] , \block[4][57] , \block[4][56] , \block[4][55] ,
         \block[4][54] , \block[4][53] , \block[4][52] , \block[4][51] ,
         \block[4][50] , \block[4][49] , \block[4][48] , \block[4][47] ,
         \block[4][46] , \block[4][45] , \block[4][44] , \block[4][43] ,
         \block[4][42] , \block[4][41] , \block[4][40] , \block[4][39] ,
         \block[4][38] , \block[4][37] , \block[4][36] , \block[4][35] ,
         \block[4][34] , \block[4][33] , \block[4][32] , \block[4][31] ,
         \block[4][30] , \block[4][29] , \block[4][28] , \block[4][27] ,
         \block[4][26] , \block[4][25] , \block[4][24] , \block[4][23] ,
         \block[4][22] , \block[4][21] , \block[4][20] , \block[4][19] ,
         \block[4][18] , \block[4][17] , \block[4][16] , \block[4][15] ,
         \block[4][14] , \block[4][13] , \block[4][12] , \block[4][11] ,
         \block[4][10] , \block[4][9] , \block[4][8] , \block[4][7] ,
         \block[4][6] , \block[4][5] , \block[4][4] , \block[4][3] ,
         \block[4][2] , \block[4][1] , \block[4][0] , \block[3][127] ,
         \block[3][126] , \block[3][125] , \block[3][124] , \block[3][123] ,
         \block[3][122] , \block[3][121] , \block[3][120] , \block[3][119] ,
         \block[3][118] , \block[3][117] , \block[3][116] , \block[3][115] ,
         \block[3][114] , \block[3][113] , \block[3][112] , \block[3][111] ,
         \block[3][110] , \block[3][109] , \block[3][108] , \block[3][107] ,
         \block[3][106] , \block[3][105] , \block[3][104] , \block[3][103] ,
         \block[3][102] , \block[3][101] , \block[3][100] , \block[3][99] ,
         \block[3][98] , \block[3][97] , \block[3][96] , \block[3][95] ,
         \block[3][94] , \block[3][93] , \block[3][92] , \block[3][91] ,
         \block[3][90] , \block[3][89] , \block[3][88] , \block[3][87] ,
         \block[3][86] , \block[3][85] , \block[3][84] , \block[3][83] ,
         \block[3][82] , \block[3][81] , \block[3][80] , \block[3][79] ,
         \block[3][78] , \block[3][77] , \block[3][76] , \block[3][75] ,
         \block[3][74] , \block[3][73] , \block[3][72] , \block[3][71] ,
         \block[3][70] , \block[3][69] , \block[3][68] , \block[3][67] ,
         \block[3][66] , \block[3][65] , \block[3][64] , \block[3][63] ,
         \block[3][62] , \block[3][61] , \block[3][60] , \block[3][59] ,
         \block[3][58] , \block[3][57] , \block[3][56] , \block[3][55] ,
         \block[3][54] , \block[3][53] , \block[3][52] , \block[3][51] ,
         \block[3][50] , \block[3][49] , \block[3][48] , \block[3][47] ,
         \block[3][46] , \block[3][45] , \block[3][44] , \block[3][43] ,
         \block[3][42] , \block[3][41] , \block[3][40] , \block[3][39] ,
         \block[3][38] , \block[3][37] , \block[3][36] , \block[3][35] ,
         \block[3][34] , \block[3][33] , \block[3][32] , \block[3][31] ,
         \block[3][30] , \block[3][29] , \block[3][28] , \block[3][27] ,
         \block[3][26] , \block[3][25] , \block[3][24] , \block[3][23] ,
         \block[3][22] , \block[3][21] , \block[3][20] , \block[3][19] ,
         \block[3][18] , \block[3][17] , \block[3][16] , \block[3][15] ,
         \block[3][14] , \block[3][13] , \block[3][12] , \block[3][11] ,
         \block[3][10] , \block[3][9] , \block[3][8] , \block[3][7] ,
         \block[3][6] , \block[3][5] , \block[3][4] , \block[3][3] ,
         \block[3][2] , \block[3][1] , \block[3][0] , \block[2][127] ,
         \block[2][126] , \block[2][125] , \block[2][124] , \block[2][123] ,
         \block[2][122] , \block[2][121] , \block[2][120] , \block[2][119] ,
         \block[2][118] , \block[2][117] , \block[2][116] , \block[2][115] ,
         \block[2][114] , \block[2][113] , \block[2][112] , \block[2][111] ,
         \block[2][110] , \block[2][109] , \block[2][108] , \block[2][107] ,
         \block[2][106] , \block[2][105] , \block[2][104] , \block[2][103] ,
         \block[2][102] , \block[2][101] , \block[2][100] , \block[2][99] ,
         \block[2][98] , \block[2][97] , \block[2][96] , \block[2][95] ,
         \block[2][94] , \block[2][93] , \block[2][92] , \block[2][91] ,
         \block[2][90] , \block[2][89] , \block[2][88] , \block[2][87] ,
         \block[2][86] , \block[2][85] , \block[2][84] , \block[2][83] ,
         \block[2][82] , \block[2][81] , \block[2][80] , \block[2][79] ,
         \block[2][78] , \block[2][77] , \block[2][76] , \block[2][75] ,
         \block[2][74] , \block[2][73] , \block[2][72] , \block[2][71] ,
         \block[2][70] , \block[2][69] , \block[2][68] , \block[2][67] ,
         \block[2][66] , \block[2][65] , \block[2][64] , \block[2][63] ,
         \block[2][62] , \block[2][61] , \block[2][60] , \block[2][59] ,
         \block[2][58] , \block[2][57] , \block[2][56] , \block[2][55] ,
         \block[2][54] , \block[2][53] , \block[2][52] , \block[2][51] ,
         \block[2][50] , \block[2][49] , \block[2][48] , \block[2][47] ,
         \block[2][46] , \block[2][45] , \block[2][44] , \block[2][43] ,
         \block[2][42] , \block[2][41] , \block[2][40] , \block[2][39] ,
         \block[2][38] , \block[2][37] , \block[2][36] , \block[2][35] ,
         \block[2][34] , \block[2][33] , \block[2][32] , \block[2][31] ,
         \block[2][30] , \block[2][29] , \block[2][28] , \block[2][27] ,
         \block[2][26] , \block[2][25] , \block[2][24] , \block[2][23] ,
         \block[2][22] , \block[2][21] , \block[2][20] , \block[2][19] ,
         \block[2][18] , \block[2][17] , \block[2][16] , \block[2][15] ,
         \block[2][14] , \block[2][13] , \block[2][12] , \block[2][11] ,
         \block[2][10] , \block[2][9] , \block[2][8] , \block[2][7] ,
         \block[2][6] , \block[2][5] , \block[2][4] , \block[2][3] ,
         \block[2][2] , \block[2][1] , \block[2][0] , \block[1][127] ,
         \block[1][126] , \block[1][125] , \block[1][124] , \block[1][123] ,
         \block[1][122] , \block[1][121] , \block[1][120] , \block[1][119] ,
         \block[1][118] , \block[1][117] , \block[1][116] , \block[1][115] ,
         \block[1][114] , \block[1][113] , \block[1][112] , \block[1][111] ,
         \block[1][110] , \block[1][109] , \block[1][108] , \block[1][107] ,
         \block[1][106] , \block[1][105] , \block[1][104] , \block[1][103] ,
         \block[1][102] , \block[1][101] , \block[1][100] , \block[1][99] ,
         \block[1][98] , \block[1][97] , \block[1][96] , \block[1][95] ,
         \block[1][94] , \block[1][93] , \block[1][92] , \block[1][91] ,
         \block[1][90] , \block[1][89] , \block[1][88] , \block[1][87] ,
         \block[1][86] , \block[1][85] , \block[1][84] , \block[1][83] ,
         \block[1][82] , \block[1][81] , \block[1][80] , \block[1][79] ,
         \block[1][78] , \block[1][77] , \block[1][76] , \block[1][75] ,
         \block[1][74] , \block[1][73] , \block[1][72] , \block[1][71] ,
         \block[1][70] , \block[1][69] , \block[1][68] , \block[1][67] ,
         \block[1][66] , \block[1][65] , \block[1][64] , \block[1][63] ,
         \block[1][62] , \block[1][61] , \block[1][60] , \block[1][59] ,
         \block[1][58] , \block[1][57] , \block[1][56] , \block[1][55] ,
         \block[1][54] , \block[1][53] , \block[1][52] , \block[1][51] ,
         \block[1][50] , \block[1][49] , \block[1][48] , \block[1][47] ,
         \block[1][46] , \block[1][45] , \block[1][44] , \block[1][43] ,
         \block[1][42] , \block[1][41] , \block[1][40] , \block[1][39] ,
         \block[1][38] , \block[1][37] , \block[1][36] , \block[1][35] ,
         \block[1][34] , \block[1][33] , \block[1][32] , \block[1][31] ,
         \block[1][30] , \block[1][29] , \block[1][28] , \block[1][27] ,
         \block[1][26] , \block[1][25] , \block[1][24] , \block[1][23] ,
         \block[1][22] , \block[1][21] , \block[1][20] , \block[1][19] ,
         \block[1][18] , \block[1][17] , \block[1][16] , \block[1][15] ,
         \block[1][14] , \block[1][13] , \block[1][12] , \block[1][11] ,
         \block[1][10] , \block[1][9] , \block[1][8] , \block[1][7] ,
         \block[1][6] , \block[1][5] , \block[1][4] , \block[1][3] ,
         \block[1][2] , \block[1][1] , \block[1][0] , \block[0][127] ,
         \block[0][126] , \block[0][125] , \block[0][124] , \block[0][123] ,
         \block[0][122] , \block[0][121] , \block[0][120] , \block[0][119] ,
         \block[0][118] , \block[0][117] , \block[0][116] , \block[0][115] ,
         \block[0][114] , \block[0][113] , \block[0][112] , \block[0][111] ,
         \block[0][110] , \block[0][109] , \block[0][108] , \block[0][107] ,
         \block[0][106] , \block[0][105] , \block[0][104] , \block[0][103] ,
         \block[0][102] , \block[0][101] , \block[0][100] , \block[0][99] ,
         \block[0][98] , \block[0][97] , \block[0][96] , \block[0][95] ,
         \block[0][94] , \block[0][93] , \block[0][92] , \block[0][91] ,
         \block[0][90] , \block[0][89] , \block[0][88] , \block[0][87] ,
         \block[0][86] , \block[0][85] , \block[0][84] , \block[0][83] ,
         \block[0][82] , \block[0][81] , \block[0][80] , \block[0][79] ,
         \block[0][78] , \block[0][77] , \block[0][76] , \block[0][75] ,
         \block[0][74] , \block[0][73] , \block[0][72] , \block[0][71] ,
         \block[0][70] , \block[0][69] , \block[0][68] , \block[0][67] ,
         \block[0][66] , \block[0][65] , \block[0][64] , \block[0][63] ,
         \block[0][62] , \block[0][61] , \block[0][60] , \block[0][59] ,
         \block[0][58] , \block[0][57] , \block[0][56] , \block[0][55] ,
         \block[0][54] , \block[0][53] , \block[0][52] , \block[0][51] ,
         \block[0][50] , \block[0][49] , \block[0][48] , \block[0][47] ,
         \block[0][46] , \block[0][45] , \block[0][44] , \block[0][43] ,
         \block[0][42] , \block[0][41] , \block[0][40] , \block[0][39] ,
         \block[0][38] , \block[0][37] , \block[0][36] , \block[0][35] ,
         \block[0][34] , \block[0][33] , \block[0][32] , \block[0][31] ,
         \block[0][30] , \block[0][29] , \block[0][28] , \block[0][27] ,
         \block[0][26] , \block[0][25] , \block[0][24] , \block[0][23] ,
         \block[0][22] , \block[0][21] , \block[0][20] , \block[0][19] ,
         \block[0][18] , \block[0][17] , \block[0][16] , \block[0][15] ,
         \block[0][14] , \block[0][13] , \block[0][12] , \block[0][11] ,
         \block[0][10] , \block[0][9] , \block[0][8] , \block[0][7] ,
         \block[0][6] , \block[0][5] , \block[0][4] , \block[0][3] ,
         \block[0][2] , \block[0][1] , \block[0][0] , N957, N960, N962, N965,
         n5, n6, n7, n9, n10, n11, n13, n17, n18, n20, n22, n24, n26, n28, n30,
         n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n74, n76, n78,
         n80, n83, n85, n87, n88, n89, n90, n99, n100, n101, n102, n111, n112,
         n113, n114, n123, n124, n125, n126, n135, n136, n137, n138, n147,
         n148, n149, n150, n159, n160, n161, n162, n171, n172, n173, n174,
         n183, n184, n185, n186, n195, n196, n197, n198, n207, n208, n209,
         n210, n219, n220, n221, n222, n231, n232, n233, n234, n243, n244,
         n245, n246, n255, n256, n257, n258, n267, n268, n269, n270, n279,
         n280, n281, n282, n291, n292, n293, n294, n303, n304, n305, n306,
         n315, n316, n317, n318, n327, n328, n329, n330, n339, n340, n341,
         n342, n351, n352, n353, n354, n363, n364, n365, n366, n375, n376,
         n377, n378, n387, n388, n389, n390, n399, n400, n401, n402, n411,
         n412, n413, n414, n423, n424, n425, n426, n435, n436, n437, n438,
         n447, n448, n449, n450, n453, n454, n455, n456, n460, n461, n465,
         n466, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n507, n508, n513, n514, n543, n544, n545, n546,
         n550, n554, n555, n556, n589, n590, n591, n592, n593, n594, n595,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639;
  wire   [1:0] wordIndex;
  wire   [24:0] dataTag;
  wire   [24:0] tag;
  wire   [127:0] mem_rdata_r;
  wire   [2:0] state;
  wire   [127:0] blockdata;
  wire   [2:0] state_next;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;

  DFFQX1 \mem_rdata_r_reg[127]  ( .D(mem_rdata[127]), .CK(clk), .Q(
        mem_rdata_r[127]) );
  DFFQX1 \mem_rdata_r_reg[126]  ( .D(mem_rdata[126]), .CK(clk), .Q(
        mem_rdata_r[126]) );
  DFFQX1 \mem_rdata_r_reg[125]  ( .D(mem_rdata[125]), .CK(clk), .Q(
        mem_rdata_r[125]) );
  DFFQX1 \mem_rdata_r_reg[124]  ( .D(mem_rdata[124]), .CK(clk), .Q(
        mem_rdata_r[124]) );
  DFFQX1 \mem_rdata_r_reg[123]  ( .D(mem_rdata[123]), .CK(clk), .Q(
        mem_rdata_r[123]) );
  DFFQX1 \mem_rdata_r_reg[122]  ( .D(mem_rdata[122]), .CK(clk), .Q(
        mem_rdata_r[122]) );
  DFFQX1 \mem_rdata_r_reg[121]  ( .D(mem_rdata[121]), .CK(clk), .Q(
        mem_rdata_r[121]) );
  DFFQX1 \mem_rdata_r_reg[120]  ( .D(mem_rdata[120]), .CK(clk), .Q(
        mem_rdata_r[120]) );
  DFFQX1 \mem_rdata_r_reg[119]  ( .D(mem_rdata[119]), .CK(clk), .Q(
        mem_rdata_r[119]) );
  DFFQX1 \mem_rdata_r_reg[118]  ( .D(mem_rdata[118]), .CK(clk), .Q(
        mem_rdata_r[118]) );
  DFFQX1 \mem_rdata_r_reg[117]  ( .D(mem_rdata[117]), .CK(clk), .Q(
        mem_rdata_r[117]) );
  DFFQX1 \mem_rdata_r_reg[116]  ( .D(mem_rdata[116]), .CK(clk), .Q(
        mem_rdata_r[116]) );
  DFFQX1 \mem_rdata_r_reg[115]  ( .D(mem_rdata[115]), .CK(clk), .Q(
        mem_rdata_r[115]) );
  DFFQX1 \mem_rdata_r_reg[114]  ( .D(mem_rdata[114]), .CK(clk), .Q(
        mem_rdata_r[114]) );
  DFFQX1 \mem_rdata_r_reg[113]  ( .D(mem_rdata[113]), .CK(clk), .Q(
        mem_rdata_r[113]) );
  DFFQX1 \mem_rdata_r_reg[112]  ( .D(mem_rdata[112]), .CK(clk), .Q(
        mem_rdata_r[112]) );
  DFFQX1 \mem_rdata_r_reg[111]  ( .D(mem_rdata[111]), .CK(clk), .Q(
        mem_rdata_r[111]) );
  DFFQX1 \mem_rdata_r_reg[110]  ( .D(mem_rdata[110]), .CK(clk), .Q(
        mem_rdata_r[110]) );
  DFFQX1 \mem_rdata_r_reg[109]  ( .D(mem_rdata[109]), .CK(clk), .Q(
        mem_rdata_r[109]) );
  DFFQX1 \mem_rdata_r_reg[108]  ( .D(mem_rdata[108]), .CK(clk), .Q(
        mem_rdata_r[108]) );
  DFFQX1 \mem_rdata_r_reg[107]  ( .D(mem_rdata[107]), .CK(clk), .Q(
        mem_rdata_r[107]) );
  DFFQX1 \mem_rdata_r_reg[106]  ( .D(mem_rdata[106]), .CK(clk), .Q(
        mem_rdata_r[106]) );
  DFFQX1 \mem_rdata_r_reg[105]  ( .D(mem_rdata[105]), .CK(clk), .Q(
        mem_rdata_r[105]) );
  DFFQX1 \mem_rdata_r_reg[104]  ( .D(mem_rdata[104]), .CK(clk), .Q(
        mem_rdata_r[104]) );
  DFFQX1 \mem_rdata_r_reg[103]  ( .D(mem_rdata[103]), .CK(clk), .Q(
        mem_rdata_r[103]) );
  DFFQX1 \mem_rdata_r_reg[102]  ( .D(mem_rdata[102]), .CK(clk), .Q(
        mem_rdata_r[102]) );
  DFFQX1 \mem_rdata_r_reg[101]  ( .D(mem_rdata[101]), .CK(clk), .Q(
        mem_rdata_r[101]) );
  DFFQX1 \mem_rdata_r_reg[100]  ( .D(mem_rdata[100]), .CK(clk), .Q(
        mem_rdata_r[100]) );
  DFFQX1 \mem_rdata_r_reg[99]  ( .D(mem_rdata[99]), .CK(clk), .Q(
        mem_rdata_r[99]) );
  DFFQX1 \mem_rdata_r_reg[98]  ( .D(mem_rdata[98]), .CK(clk), .Q(
        mem_rdata_r[98]) );
  DFFQX1 \mem_rdata_r_reg[97]  ( .D(mem_rdata[97]), .CK(clk), .Q(
        mem_rdata_r[97]) );
  DFFQX1 \mem_rdata_r_reg[96]  ( .D(mem_rdata[96]), .CK(clk), .Q(
        mem_rdata_r[96]) );
  DFFQX1 \mem_rdata_r_reg[95]  ( .D(mem_rdata[95]), .CK(clk), .Q(
        mem_rdata_r[95]) );
  DFFQX1 \mem_rdata_r_reg[94]  ( .D(mem_rdata[94]), .CK(clk), .Q(
        mem_rdata_r[94]) );
  DFFQX1 \mem_rdata_r_reg[93]  ( .D(mem_rdata[93]), .CK(clk), .Q(
        mem_rdata_r[93]) );
  DFFQX1 \mem_rdata_r_reg[92]  ( .D(mem_rdata[92]), .CK(clk), .Q(
        mem_rdata_r[92]) );
  DFFQX1 \mem_rdata_r_reg[91]  ( .D(mem_rdata[91]), .CK(clk), .Q(
        mem_rdata_r[91]) );
  DFFQX1 \mem_rdata_r_reg[90]  ( .D(mem_rdata[90]), .CK(clk), .Q(
        mem_rdata_r[90]) );
  DFFQX1 \mem_rdata_r_reg[89]  ( .D(mem_rdata[89]), .CK(clk), .Q(
        mem_rdata_r[89]) );
  DFFQX1 \mem_rdata_r_reg[88]  ( .D(mem_rdata[88]), .CK(clk), .Q(
        mem_rdata_r[88]) );
  DFFQX1 \mem_rdata_r_reg[87]  ( .D(mem_rdata[87]), .CK(clk), .Q(
        mem_rdata_r[87]) );
  DFFQX1 \mem_rdata_r_reg[86]  ( .D(mem_rdata[86]), .CK(clk), .Q(
        mem_rdata_r[86]) );
  DFFQX1 \mem_rdata_r_reg[85]  ( .D(mem_rdata[85]), .CK(clk), .Q(
        mem_rdata_r[85]) );
  DFFQX1 \mem_rdata_r_reg[84]  ( .D(mem_rdata[84]), .CK(clk), .Q(
        mem_rdata_r[84]) );
  DFFQX1 \mem_rdata_r_reg[83]  ( .D(mem_rdata[83]), .CK(clk), .Q(
        mem_rdata_r[83]) );
  DFFQX1 \mem_rdata_r_reg[82]  ( .D(mem_rdata[82]), .CK(clk), .Q(
        mem_rdata_r[82]) );
  DFFQX1 \mem_rdata_r_reg[81]  ( .D(mem_rdata[81]), .CK(clk), .Q(
        mem_rdata_r[81]) );
  DFFQX1 \mem_rdata_r_reg[80]  ( .D(mem_rdata[80]), .CK(clk), .Q(
        mem_rdata_r[80]) );
  DFFQX1 \mem_rdata_r_reg[79]  ( .D(mem_rdata[79]), .CK(clk), .Q(
        mem_rdata_r[79]) );
  DFFQX1 \mem_rdata_r_reg[78]  ( .D(mem_rdata[78]), .CK(clk), .Q(
        mem_rdata_r[78]) );
  DFFQX1 \mem_rdata_r_reg[77]  ( .D(mem_rdata[77]), .CK(clk), .Q(
        mem_rdata_r[77]) );
  DFFQX1 \mem_rdata_r_reg[76]  ( .D(mem_rdata[76]), .CK(clk), .Q(
        mem_rdata_r[76]) );
  DFFQX1 \mem_rdata_r_reg[75]  ( .D(mem_rdata[75]), .CK(clk), .Q(
        mem_rdata_r[75]) );
  DFFQX1 \mem_rdata_r_reg[74]  ( .D(mem_rdata[74]), .CK(clk), .Q(
        mem_rdata_r[74]) );
  DFFQX1 \mem_rdata_r_reg[73]  ( .D(mem_rdata[73]), .CK(clk), .Q(
        mem_rdata_r[73]) );
  DFFQX1 \mem_rdata_r_reg[72]  ( .D(mem_rdata[72]), .CK(clk), .Q(
        mem_rdata_r[72]) );
  DFFQX1 \mem_rdata_r_reg[71]  ( .D(mem_rdata[71]), .CK(clk), .Q(
        mem_rdata_r[71]) );
  DFFQX1 \mem_rdata_r_reg[70]  ( .D(mem_rdata[70]), .CK(clk), .Q(
        mem_rdata_r[70]) );
  DFFQX1 \mem_rdata_r_reg[69]  ( .D(mem_rdata[69]), .CK(clk), .Q(
        mem_rdata_r[69]) );
  DFFQX1 \mem_rdata_r_reg[68]  ( .D(mem_rdata[68]), .CK(clk), .Q(
        mem_rdata_r[68]) );
  DFFQX1 \mem_rdata_r_reg[67]  ( .D(mem_rdata[67]), .CK(clk), .Q(
        mem_rdata_r[67]) );
  DFFQX1 \mem_rdata_r_reg[66]  ( .D(mem_rdata[66]), .CK(clk), .Q(
        mem_rdata_r[66]) );
  DFFQX1 \mem_rdata_r_reg[65]  ( .D(mem_rdata[65]), .CK(clk), .Q(
        mem_rdata_r[65]) );
  DFFQX1 \mem_rdata_r_reg[64]  ( .D(mem_rdata[64]), .CK(clk), .Q(
        mem_rdata_r[64]) );
  DFFQX1 \mem_rdata_r_reg[63]  ( .D(mem_rdata[63]), .CK(clk), .Q(
        mem_rdata_r[63]) );
  DFFQX1 \mem_rdata_r_reg[62]  ( .D(mem_rdata[62]), .CK(clk), .Q(
        mem_rdata_r[62]) );
  DFFQX1 \mem_rdata_r_reg[61]  ( .D(mem_rdata[61]), .CK(clk), .Q(
        mem_rdata_r[61]) );
  DFFQX1 \mem_rdata_r_reg[60]  ( .D(mem_rdata[60]), .CK(clk), .Q(
        mem_rdata_r[60]) );
  DFFQX1 \mem_rdata_r_reg[59]  ( .D(mem_rdata[59]), .CK(clk), .Q(
        mem_rdata_r[59]) );
  DFFQX1 \mem_rdata_r_reg[58]  ( .D(mem_rdata[58]), .CK(clk), .Q(
        mem_rdata_r[58]) );
  DFFQX1 \mem_rdata_r_reg[57]  ( .D(mem_rdata[57]), .CK(clk), .Q(
        mem_rdata_r[57]) );
  DFFQX1 \mem_rdata_r_reg[56]  ( .D(mem_rdata[56]), .CK(clk), .Q(
        mem_rdata_r[56]) );
  DFFQX1 \mem_rdata_r_reg[55]  ( .D(mem_rdata[55]), .CK(clk), .Q(
        mem_rdata_r[55]) );
  DFFQX1 \mem_rdata_r_reg[54]  ( .D(mem_rdata[54]), .CK(clk), .Q(
        mem_rdata_r[54]) );
  DFFQX1 \mem_rdata_r_reg[53]  ( .D(mem_rdata[53]), .CK(clk), .Q(
        mem_rdata_r[53]) );
  DFFQX1 \mem_rdata_r_reg[52]  ( .D(mem_rdata[52]), .CK(clk), .Q(
        mem_rdata_r[52]) );
  DFFQX1 \mem_rdata_r_reg[51]  ( .D(mem_rdata[51]), .CK(clk), .Q(
        mem_rdata_r[51]) );
  DFFQX1 \mem_rdata_r_reg[50]  ( .D(mem_rdata[50]), .CK(clk), .Q(
        mem_rdata_r[50]) );
  DFFQX1 \mem_rdata_r_reg[49]  ( .D(mem_rdata[49]), .CK(clk), .Q(
        mem_rdata_r[49]) );
  DFFQX1 \mem_rdata_r_reg[48]  ( .D(mem_rdata[48]), .CK(clk), .Q(
        mem_rdata_r[48]) );
  DFFQX1 \mem_rdata_r_reg[47]  ( .D(mem_rdata[47]), .CK(clk), .Q(
        mem_rdata_r[47]) );
  DFFQX1 \mem_rdata_r_reg[46]  ( .D(mem_rdata[46]), .CK(clk), .Q(
        mem_rdata_r[46]) );
  DFFQX1 \mem_rdata_r_reg[45]  ( .D(mem_rdata[45]), .CK(clk), .Q(
        mem_rdata_r[45]) );
  DFFQX1 \mem_rdata_r_reg[44]  ( .D(mem_rdata[44]), .CK(clk), .Q(
        mem_rdata_r[44]) );
  DFFQX1 \mem_rdata_r_reg[43]  ( .D(mem_rdata[43]), .CK(clk), .Q(
        mem_rdata_r[43]) );
  DFFQX1 \mem_rdata_r_reg[42]  ( .D(mem_rdata[42]), .CK(clk), .Q(
        mem_rdata_r[42]) );
  DFFQX1 \mem_rdata_r_reg[41]  ( .D(mem_rdata[41]), .CK(clk), .Q(
        mem_rdata_r[41]) );
  DFFQX1 \mem_rdata_r_reg[40]  ( .D(mem_rdata[40]), .CK(clk), .Q(
        mem_rdata_r[40]) );
  DFFQX1 \mem_rdata_r_reg[39]  ( .D(mem_rdata[39]), .CK(clk), .Q(
        mem_rdata_r[39]) );
  DFFQX1 \mem_rdata_r_reg[38]  ( .D(mem_rdata[38]), .CK(clk), .Q(
        mem_rdata_r[38]) );
  DFFQX1 \mem_rdata_r_reg[37]  ( .D(mem_rdata[37]), .CK(clk), .Q(
        mem_rdata_r[37]) );
  DFFQX1 \mem_rdata_r_reg[36]  ( .D(mem_rdata[36]), .CK(clk), .Q(
        mem_rdata_r[36]) );
  DFFQX1 \mem_rdata_r_reg[35]  ( .D(mem_rdata[35]), .CK(clk), .Q(
        mem_rdata_r[35]) );
  DFFQX1 \mem_rdata_r_reg[34]  ( .D(mem_rdata[34]), .CK(clk), .Q(
        mem_rdata_r[34]) );
  DFFQX1 \mem_rdata_r_reg[33]  ( .D(mem_rdata[33]), .CK(clk), .Q(
        mem_rdata_r[33]) );
  DFFQX1 \mem_rdata_r_reg[32]  ( .D(mem_rdata[32]), .CK(clk), .Q(
        mem_rdata_r[32]) );
  DFFQX1 \mem_rdata_r_reg[31]  ( .D(mem_rdata[31]), .CK(clk), .Q(
        mem_rdata_r[31]) );
  DFFQX1 \mem_rdata_r_reg[30]  ( .D(mem_rdata[30]), .CK(clk), .Q(
        mem_rdata_r[30]) );
  DFFQX1 \mem_rdata_r_reg[29]  ( .D(mem_rdata[29]), .CK(clk), .Q(
        mem_rdata_r[29]) );
  DFFQX1 \mem_rdata_r_reg[28]  ( .D(mem_rdata[28]), .CK(clk), .Q(
        mem_rdata_r[28]) );
  DFFQX1 \mem_rdata_r_reg[27]  ( .D(mem_rdata[27]), .CK(clk), .Q(
        mem_rdata_r[27]) );
  DFFQX1 \mem_rdata_r_reg[26]  ( .D(mem_rdata[26]), .CK(clk), .Q(
        mem_rdata_r[26]) );
  DFFQX1 \mem_rdata_r_reg[25]  ( .D(mem_rdata[25]), .CK(clk), .Q(
        mem_rdata_r[25]) );
  DFFQX1 \mem_rdata_r_reg[24]  ( .D(mem_rdata[24]), .CK(clk), .Q(
        mem_rdata_r[24]) );
  DFFQX1 \mem_rdata_r_reg[23]  ( .D(mem_rdata[23]), .CK(clk), .Q(
        mem_rdata_r[23]) );
  DFFQX1 \mem_rdata_r_reg[22]  ( .D(mem_rdata[22]), .CK(clk), .Q(
        mem_rdata_r[22]) );
  DFFQX1 \mem_rdata_r_reg[21]  ( .D(mem_rdata[21]), .CK(clk), .Q(
        mem_rdata_r[21]) );
  DFFQX1 \mem_rdata_r_reg[20]  ( .D(mem_rdata[20]), .CK(clk), .Q(
        mem_rdata_r[20]) );
  DFFQX1 \mem_rdata_r_reg[19]  ( .D(mem_rdata[19]), .CK(clk), .Q(
        mem_rdata_r[19]) );
  DFFQX1 \mem_rdata_r_reg[18]  ( .D(mem_rdata[18]), .CK(clk), .Q(
        mem_rdata_r[18]) );
  DFFQX1 \mem_rdata_r_reg[17]  ( .D(mem_rdata[17]), .CK(clk), .Q(
        mem_rdata_r[17]) );
  DFFQX1 \mem_rdata_r_reg[16]  ( .D(mem_rdata[16]), .CK(clk), .Q(
        mem_rdata_r[16]) );
  DFFQX1 \mem_rdata_r_reg[15]  ( .D(mem_rdata[15]), .CK(clk), .Q(
        mem_rdata_r[15]) );
  DFFQX1 \mem_rdata_r_reg[14]  ( .D(mem_rdata[14]), .CK(clk), .Q(
        mem_rdata_r[14]) );
  DFFQX1 \mem_rdata_r_reg[13]  ( .D(mem_rdata[13]), .CK(clk), .Q(
        mem_rdata_r[13]) );
  DFFQX1 \mem_rdata_r_reg[12]  ( .D(mem_rdata[12]), .CK(clk), .Q(
        mem_rdata_r[12]) );
  DFFQX1 \mem_rdata_r_reg[11]  ( .D(mem_rdata[11]), .CK(clk), .Q(
        mem_rdata_r[11]) );
  DFFQX1 \mem_rdata_r_reg[10]  ( .D(mem_rdata[10]), .CK(clk), .Q(
        mem_rdata_r[10]) );
  DFFQX1 \mem_rdata_r_reg[9]  ( .D(mem_rdata[9]), .CK(clk), .Q(mem_rdata_r[9])
         );
  DFFQX1 \mem_rdata_r_reg[8]  ( .D(mem_rdata[8]), .CK(clk), .Q(mem_rdata_r[8])
         );
  DFFQX1 \mem_rdata_r_reg[7]  ( .D(mem_rdata[7]), .CK(clk), .Q(mem_rdata_r[7])
         );
  DFFQX1 \mem_rdata_r_reg[6]  ( .D(mem_rdata[6]), .CK(clk), .Q(mem_rdata_r[6])
         );
  DFFQX1 \mem_rdata_r_reg[5]  ( .D(mem_rdata[5]), .CK(clk), .Q(mem_rdata_r[5])
         );
  DFFQX1 \mem_rdata_r_reg[4]  ( .D(mem_rdata[4]), .CK(clk), .Q(mem_rdata_r[4])
         );
  DFFQX1 \mem_rdata_r_reg[3]  ( .D(mem_rdata[3]), .CK(clk), .Q(mem_rdata_r[3])
         );
  DFFQX1 \mem_rdata_r_reg[2]  ( .D(mem_rdata[2]), .CK(clk), .Q(mem_rdata_r[2])
         );
  DFFQX1 \mem_rdata_r_reg[1]  ( .D(mem_rdata[1]), .CK(clk), .Q(mem_rdata_r[1])
         );
  DFFQX1 \mem_rdata_r_reg[0]  ( .D(mem_rdata[0]), .CK(clk), .Q(mem_rdata_r[0])
         );
  DFFX1 \proc_wdata_r_reg[31]  ( .D(proc_wdata[31]), .CK(clk), .QN(n1476) );
  DFFX1 \proc_wdata_r_reg[30]  ( .D(proc_wdata[30]), .CK(clk), .QN(n1477) );
  DFFX1 \proc_wdata_r_reg[29]  ( .D(proc_wdata[29]), .CK(clk), .QN(n1478) );
  DFFX1 \proc_wdata_r_reg[28]  ( .D(proc_wdata[28]), .CK(clk), .QN(n1479) );
  DFFX1 \proc_wdata_r_reg[27]  ( .D(proc_wdata[27]), .CK(clk), .QN(n1480) );
  DFFX1 \proc_wdata_r_reg[26]  ( .D(proc_wdata[26]), .CK(clk), .QN(n1481) );
  DFFX1 \proc_wdata_r_reg[25]  ( .D(proc_wdata[25]), .CK(clk), .QN(n1482) );
  DFFX1 \proc_wdata_r_reg[24]  ( .D(proc_wdata[24]), .CK(clk), .QN(n1483) );
  DFFX1 \proc_wdata_r_reg[23]  ( .D(proc_wdata[23]), .CK(clk), .QN(n1484) );
  DFFX1 \proc_wdata_r_reg[22]  ( .D(proc_wdata[22]), .CK(clk), .QN(n1485) );
  DFFX1 \proc_wdata_r_reg[21]  ( .D(proc_wdata[21]), .CK(clk), .QN(n1486) );
  DFFX1 \proc_wdata_r_reg[20]  ( .D(proc_wdata[20]), .CK(clk), .QN(n1487) );
  DFFX1 \proc_wdata_r_reg[19]  ( .D(proc_wdata[19]), .CK(clk), .QN(n1488) );
  DFFX1 \proc_wdata_r_reg[18]  ( .D(proc_wdata[18]), .CK(clk), .QN(n1489) );
  DFFX1 \proc_wdata_r_reg[17]  ( .D(proc_wdata[17]), .CK(clk), .QN(n1490) );
  DFFX1 \proc_wdata_r_reg[16]  ( .D(proc_wdata[16]), .CK(clk), .QN(n1491) );
  DFFX1 \proc_wdata_r_reg[15]  ( .D(proc_wdata[15]), .CK(clk), .QN(n1492) );
  DFFX1 \proc_wdata_r_reg[14]  ( .D(proc_wdata[14]), .CK(clk), .QN(n1493) );
  DFFX1 \proc_wdata_r_reg[13]  ( .D(proc_wdata[13]), .CK(clk), .QN(n1494) );
  DFFX1 \proc_wdata_r_reg[12]  ( .D(proc_wdata[12]), .CK(clk), .QN(n1495) );
  DFFX1 \proc_wdata_r_reg[11]  ( .D(proc_wdata[11]), .CK(clk), .QN(n1496) );
  DFFX1 \proc_wdata_r_reg[10]  ( .D(proc_wdata[10]), .CK(clk), .QN(n1497) );
  DFFX1 \proc_wdata_r_reg[9]  ( .D(proc_wdata[9]), .CK(clk), .QN(n1498) );
  DFFX1 \proc_wdata_r_reg[8]  ( .D(proc_wdata[8]), .CK(clk), .QN(n1499) );
  DFFX1 \proc_wdata_r_reg[7]  ( .D(proc_wdata[7]), .CK(clk), .QN(n1500) );
  DFFX1 \proc_wdata_r_reg[6]  ( .D(proc_wdata[6]), .CK(clk), .QN(n1501) );
  DFFX1 \proc_wdata_r_reg[5]  ( .D(proc_wdata[5]), .CK(clk), .QN(n1502) );
  DFFX1 \proc_wdata_r_reg[4]  ( .D(proc_wdata[4]), .CK(clk), .QN(n1503) );
  DFFX1 \proc_wdata_r_reg[3]  ( .D(proc_wdata[3]), .CK(clk), .QN(n1504) );
  DFFX1 \proc_wdata_r_reg[2]  ( .D(proc_wdata[2]), .CK(clk), .QN(n1505) );
  DFFX1 \proc_wdata_r_reg[1]  ( .D(proc_wdata[1]), .CK(clk), .QN(n1506) );
  DFFX1 \proc_wdata_r_reg[0]  ( .D(proc_wdata[0]), .CK(clk), .QN(n1507) );
  DFFQX1 \proc_rdata_reg[31]  ( .D(n682), .CK(clk), .Q(proc_rdata[31]) );
  DFFQX1 \proc_rdata_reg[30]  ( .D(n681), .CK(clk), .Q(proc_rdata[30]) );
  DFFQX1 \proc_rdata_reg[29]  ( .D(n680), .CK(clk), .Q(proc_rdata[29]) );
  DFFQX1 \proc_rdata_reg[28]  ( .D(n679), .CK(clk), .Q(proc_rdata[28]) );
  DFFQX1 \proc_rdata_reg[27]  ( .D(n678), .CK(clk), .Q(proc_rdata[27]) );
  DFFQX1 \proc_rdata_reg[26]  ( .D(n677), .CK(clk), .Q(proc_rdata[26]) );
  DFFQX1 \proc_rdata_reg[25]  ( .D(n676), .CK(clk), .Q(proc_rdata[25]) );
  DFFQX1 \proc_rdata_reg[24]  ( .D(n675), .CK(clk), .Q(proc_rdata[24]) );
  EDFFX1 \block_reg[3][127]  ( .D(block_next[127]), .E(n1271), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFX1 \block_reg[7][127]  ( .D(block_next[127]), .E(n1237), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFX1 \block_reg[3][126]  ( .D(block_next[126]), .E(n1271), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFX1 \block_reg[7][126]  ( .D(block_next[126]), .E(n1237), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFX1 \block_reg[3][125]  ( .D(block_next[125]), .E(n1271), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFX1 \block_reg[7][125]  ( .D(block_next[125]), .E(n1237), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFX1 \block_reg[3][124]  ( .D(block_next[124]), .E(n1275), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFX1 \block_reg[7][124]  ( .D(block_next[124]), .E(n1241), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFX1 \block_reg[3][123]  ( .D(block_next[123]), .E(n1273), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFX1 \block_reg[7][123]  ( .D(block_next[123]), .E(n1239), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFX1 \block_reg[3][122]  ( .D(block_next[122]), .E(n1272), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFX1 \block_reg[7][122]  ( .D(block_next[122]), .E(n1238), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFX1 \block_reg[3][121]  ( .D(block_next[121]), .E(n1274), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFX1 \block_reg[7][121]  ( .D(block_next[121]), .E(n1240), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFX1 \block_reg[3][120]  ( .D(block_next[120]), .E(n1274), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFX1 \block_reg[7][120]  ( .D(block_next[120]), .E(n1240), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFX1 \block_reg[3][119]  ( .D(block_next[119]), .E(n1276), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFX1 \block_reg[7][119]  ( .D(block_next[119]), .E(n1242), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFX1 \block_reg[3][118]  ( .D(block_next[118]), .E(n1277), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFX1 \block_reg[7][118]  ( .D(block_next[118]), .E(n1243), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFX1 \block_reg[3][117]  ( .D(block_next[117]), .E(n1279), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFX1 \block_reg[7][117]  ( .D(block_next[117]), .E(n1245), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFX1 \block_reg[3][116]  ( .D(block_next[116]), .E(n1277), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFX1 \block_reg[7][116]  ( .D(block_next[116]), .E(n1243), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFX1 \block_reg[3][115]  ( .D(block_next[115]), .E(n1279), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFX1 \block_reg[7][115]  ( .D(block_next[115]), .E(n1245), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFX1 \block_reg[3][114]  ( .D(block_next[114]), .E(n1278), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFX1 \block_reg[7][114]  ( .D(block_next[114]), .E(n1244), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFX1 \block_reg[3][113]  ( .D(block_next[113]), .E(n1271), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFX1 \block_reg[7][113]  ( .D(block_next[113]), .E(n1237), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFX1 \block_reg[3][112]  ( .D(block_next[112]), .E(n1271), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFX1 \block_reg[7][112]  ( .D(block_next[112]), .E(n1237), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFX1 \block_reg[3][111]  ( .D(block_next[111]), .E(n1275), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFX1 \block_reg[7][111]  ( .D(block_next[111]), .E(n1241), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFX1 \block_reg[3][110]  ( .D(block_next[110]), .E(n1273), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFX1 \block_reg[7][110]  ( .D(block_next[110]), .E(n1239), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFX1 \block_reg[3][109]  ( .D(block_next[109]), .E(n1272), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFX1 \block_reg[7][109]  ( .D(block_next[109]), .E(n1238), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFX1 \block_reg[3][108]  ( .D(block_next[108]), .E(n1274), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFX1 \block_reg[7][108]  ( .D(block_next[108]), .E(n1240), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFX1 \block_reg[3][107]  ( .D(block_next[107]), .E(n1276), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFX1 \block_reg[7][107]  ( .D(block_next[107]), .E(n1242), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFX1 \block_reg[3][106]  ( .D(block_next[106]), .E(n1276), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFX1 \block_reg[7][106]  ( .D(block_next[106]), .E(n1242), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFX1 \block_reg[3][105]  ( .D(block_next[105]), .E(n1277), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFX1 \block_reg[7][105]  ( .D(block_next[105]), .E(n1243), .CK(clk), .Q(
        \block[7][105] ) );
  EDFFX1 \block_reg[3][104]  ( .D(block_next[104]), .E(n1279), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFX1 \block_reg[7][104]  ( .D(block_next[104]), .E(n1245), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFX1 \block_reg[3][103]  ( .D(block_next[103]), .E(n1278), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFX1 \block_reg[7][103]  ( .D(block_next[103]), .E(n1244), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFX1 \block_reg[3][102]  ( .D(block_next[102]), .E(n1278), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFX1 \block_reg[7][102]  ( .D(block_next[102]), .E(n1244), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFX1 \block_reg[3][101]  ( .D(block_next[101]), .E(n1278), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFX1 \block_reg[7][101]  ( .D(block_next[101]), .E(n1244), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFX1 \block_reg[3][100]  ( .D(block_next[100]), .E(n1278), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFX1 \block_reg[7][100]  ( .D(block_next[100]), .E(n1244), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFX1 \block_reg[3][99]  ( .D(block_next[99]), .E(n1278), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFX1 \block_reg[7][99]  ( .D(block_next[99]), .E(n1244), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFX1 \block_reg[3][98]  ( .D(block_next[98]), .E(n1278), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFX1 \block_reg[7][98]  ( .D(block_next[98]), .E(n1244), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFX1 \block_reg[3][97]  ( .D(block_next[97]), .E(n1278), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFX1 \block_reg[7][97]  ( .D(block_next[97]), .E(n1244), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFX1 \block_reg[3][96]  ( .D(block_next[96]), .E(n1278), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFX1 \block_reg[7][96]  ( .D(block_next[96]), .E(n1244), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFX1 \block_reg[3][95]  ( .D(block_next[95]), .E(n1278), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFX1 \block_reg[7][95]  ( .D(block_next[95]), .E(n1244), .CK(clk), .Q(
        \block[7][95] ) );
  EDFFX1 \block_reg[3][94]  ( .D(block_next[94]), .E(n1278), .CK(clk), .Q(
        \block[3][94] ) );
  EDFFX1 \block_reg[7][94]  ( .D(block_next[94]), .E(n1244), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFX1 \block_reg[3][93]  ( .D(block_next[93]), .E(n1278), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFX1 \block_reg[7][93]  ( .D(block_next[93]), .E(n1244), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFX1 \block_reg[3][92]  ( .D(block_next[92]), .E(n1278), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFX1 \block_reg[7][92]  ( .D(block_next[92]), .E(n1244), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFX1 \block_reg[3][91]  ( .D(block_next[91]), .E(n1278), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFX1 \block_reg[7][91]  ( .D(block_next[91]), .E(n1244), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFX1 \block_reg[3][90]  ( .D(block_next[90]), .E(n1277), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFX1 \block_reg[7][90]  ( .D(block_next[90]), .E(n1243), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFX1 \block_reg[3][89]  ( .D(block_next[89]), .E(n1277), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFX1 \block_reg[7][89]  ( .D(block_next[89]), .E(n1243), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFX1 \block_reg[3][88]  ( .D(block_next[88]), .E(n1277), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFX1 \block_reg[7][88]  ( .D(block_next[88]), .E(n1243), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFX1 \block_reg[3][87]  ( .D(block_next[87]), .E(n1277), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFX1 \block_reg[7][87]  ( .D(block_next[87]), .E(n1243), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFX1 \block_reg[3][86]  ( .D(block_next[86]), .E(n1277), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFX1 \block_reg[7][86]  ( .D(block_next[86]), .E(n1243), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFX1 \block_reg[3][85]  ( .D(block_next[85]), .E(n1277), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFX1 \block_reg[7][85]  ( .D(block_next[85]), .E(n1243), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFX1 \block_reg[3][84]  ( .D(block_next[84]), .E(n1277), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFX1 \block_reg[7][84]  ( .D(block_next[84]), .E(n1243), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFX1 \block_reg[3][83]  ( .D(block_next[83]), .E(n1277), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFX1 \block_reg[7][83]  ( .D(block_next[83]), .E(n1243), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFX1 \block_reg[3][82]  ( .D(block_next[82]), .E(n1277), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFX1 \block_reg[7][82]  ( .D(block_next[82]), .E(n1243), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFX1 \block_reg[3][81]  ( .D(block_next[81]), .E(n1277), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFX1 \block_reg[7][81]  ( .D(block_next[81]), .E(n1243), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFX1 \block_reg[3][80]  ( .D(block_next[80]), .E(n1277), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFX1 \block_reg[7][80]  ( .D(block_next[80]), .E(n1243), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFX1 \block_reg[3][79]  ( .D(block_next[79]), .E(n1277), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFX1 \block_reg[7][79]  ( .D(block_next[79]), .E(n1243), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFX1 \block_reg[3][78]  ( .D(block_next[78]), .E(n1277), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFX1 \block_reg[7][78]  ( .D(block_next[78]), .E(n1243), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFX1 \block_reg[3][77]  ( .D(block_next[77]), .E(n1278), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFX1 \block_reg[7][77]  ( .D(block_next[77]), .E(n1244), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFX1 \block_reg[3][76]  ( .D(block_next[76]), .E(n1275), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFX1 \block_reg[7][76]  ( .D(block_next[76]), .E(n1241), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFX1 \block_reg[3][75]  ( .D(block_next[75]), .E(n1273), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFX1 \block_reg[7][75]  ( .D(block_next[75]), .E(n1239), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFX1 \block_reg[3][74]  ( .D(block_next[74]), .E(n1272), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFX1 \block_reg[7][74]  ( .D(block_next[74]), .E(n1238), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFX1 \block_reg[3][73]  ( .D(block_next[73]), .E(n1274), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFX1 \block_reg[7][73]  ( .D(block_next[73]), .E(n1240), .CK(clk), .Q(
        \block[7][73] ) );
  EDFFX1 \block_reg[3][72]  ( .D(block_next[72]), .E(n1276), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFX1 \block_reg[7][72]  ( .D(block_next[72]), .E(n1242), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFX1 \block_reg[3][71]  ( .D(block_next[71]), .E(n1277), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFX1 \block_reg[7][71]  ( .D(block_next[71]), .E(n1243), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFX1 \block_reg[3][70]  ( .D(block_next[70]), .E(n1279), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFX1 \block_reg[7][70]  ( .D(block_next[70]), .E(n1245), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFX1 \block_reg[3][69]  ( .D(block_next[69]), .E(n1278), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFX1 \block_reg[7][69]  ( .D(block_next[69]), .E(n1244), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFX1 \block_reg[3][68]  ( .D(block_next[68]), .E(n1271), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFX1 \block_reg[7][68]  ( .D(block_next[68]), .E(n1237), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFX1 \block_reg[3][67]  ( .D(block_next[67]), .E(n1275), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFX1 \block_reg[7][67]  ( .D(block_next[67]), .E(n1241), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFX1 \block_reg[3][66]  ( .D(block_next[66]), .E(n1273), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFX1 \block_reg[7][66]  ( .D(block_next[66]), .E(n1239), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFX1 \block_reg[3][65]  ( .D(block_next[65]), .E(n1272), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFX1 \block_reg[7][65]  ( .D(block_next[65]), .E(n1238), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFX1 \block_reg[3][64]  ( .D(block_next[64]), .E(n1276), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[7][64]  ( .D(block_next[64]), .E(n1242), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFX1 \block_reg[3][63]  ( .D(block_next[63]), .E(n1276), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFX1 \block_reg[7][63]  ( .D(block_next[63]), .E(n1242), .CK(clk), .Q(
        \block[7][63] ) );
  EDFFX1 \block_reg[3][62]  ( .D(block_next[62]), .E(n1276), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFX1 \block_reg[7][62]  ( .D(block_next[62]), .E(n1242), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFX1 \block_reg[3][61]  ( .D(block_next[61]), .E(n1276), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFX1 \block_reg[7][61]  ( .D(block_next[61]), .E(n1242), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFX1 \block_reg[3][60]  ( .D(block_next[60]), .E(n1276), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFX1 \block_reg[7][60]  ( .D(block_next[60]), .E(n1242), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFX1 \block_reg[3][59]  ( .D(block_next[59]), .E(n1276), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFX1 \block_reg[7][59]  ( .D(block_next[59]), .E(n1242), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFX1 \block_reg[3][58]  ( .D(block_next[58]), .E(n1276), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFX1 \block_reg[7][58]  ( .D(block_next[58]), .E(n1242), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFX1 \block_reg[3][57]  ( .D(block_next[57]), .E(n1276), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFX1 \block_reg[7][57]  ( .D(block_next[57]), .E(n1242), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFX1 \block_reg[3][56]  ( .D(block_next[56]), .E(n1276), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFX1 \block_reg[7][56]  ( .D(block_next[56]), .E(n1242), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFX1 \block_reg[3][55]  ( .D(block_next[55]), .E(n1276), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFX1 \block_reg[7][55]  ( .D(block_next[55]), .E(n1242), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFX1 \block_reg[3][54]  ( .D(block_next[54]), .E(n1276), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFX1 \block_reg[7][54]  ( .D(block_next[54]), .E(n1242), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n1276), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n1242), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n1276), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n1242), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[3][51]  ( .D(block_next[51]), .E(n1275), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFX1 \block_reg[7][51]  ( .D(block_next[51]), .E(n1241), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFX1 \block_reg[3][50]  ( .D(block_next[50]), .E(n1275), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFX1 \block_reg[7][50]  ( .D(block_next[50]), .E(n1241), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n1275), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n1241), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[3][48]  ( .D(block_next[48]), .E(n1275), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFX1 \block_reg[7][48]  ( .D(block_next[48]), .E(n1241), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFX1 \block_reg[3][47]  ( .D(block_next[47]), .E(n1275), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFX1 \block_reg[7][47]  ( .D(block_next[47]), .E(n1241), .CK(clk), .Q(
        \block[7][47] ) );
  EDFFX1 \block_reg[3][46]  ( .D(block_next[46]), .E(n1275), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFX1 \block_reg[7][46]  ( .D(block_next[46]), .E(n1241), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFX1 \block_reg[3][45]  ( .D(block_next[45]), .E(n1275), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFX1 \block_reg[7][45]  ( .D(block_next[45]), .E(n1241), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFX1 \block_reg[3][44]  ( .D(block_next[44]), .E(n1275), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFX1 \block_reg[7][44]  ( .D(block_next[44]), .E(n1241), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFX1 \block_reg[3][43]  ( .D(block_next[43]), .E(n1275), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFX1 \block_reg[7][43]  ( .D(block_next[43]), .E(n1241), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFX1 \block_reg[3][42]  ( .D(block_next[42]), .E(n1275), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFX1 \block_reg[7][42]  ( .D(block_next[42]), .E(n1241), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n1275), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n1241), .CK(clk), .Q(
        \block[7][41] ) );
  EDFFX1 \block_reg[3][40]  ( .D(block_next[40]), .E(n1275), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFX1 \block_reg[7][40]  ( .D(block_next[40]), .E(n1241), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFX1 \block_reg[3][39]  ( .D(block_next[39]), .E(n1275), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFX1 \block_reg[7][39]  ( .D(block_next[39]), .E(n1241), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n1274), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n1240), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n1274), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n1240), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n1274), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n1240), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n1274), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n1240), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n1274), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n1240), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFX1 \block_reg[3][33]  ( .D(block_next[33]), .E(n1274), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFX1 \block_reg[7][33]  ( .D(block_next[33]), .E(n1240), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n1274), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n1240), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[3][31]  ( .D(block_next[31]), .E(n1274), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFX1 \block_reg[7][31]  ( .D(block_next[31]), .E(n1240), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFX1 \block_reg[3][30]  ( .D(block_next[30]), .E(n1274), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFX1 \block_reg[7][30]  ( .D(block_next[30]), .E(n1240), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFX1 \block_reg[3][29]  ( .D(block_next[29]), .E(n1274), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFX1 \block_reg[7][29]  ( .D(block_next[29]), .E(n1240), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFX1 \block_reg[3][28]  ( .D(block_next[28]), .E(n1274), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFX1 \block_reg[7][28]  ( .D(block_next[28]), .E(n1240), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFX1 \block_reg[3][27]  ( .D(block_next[27]), .E(n1274), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFX1 \block_reg[7][27]  ( .D(block_next[27]), .E(n1240), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFX1 \block_reg[3][26]  ( .D(block_next[26]), .E(n1274), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFX1 \block_reg[7][26]  ( .D(block_next[26]), .E(n1240), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFX1 \block_reg[3][25]  ( .D(block_next[25]), .E(n1273), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFX1 \block_reg[7][25]  ( .D(block_next[25]), .E(n1239), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFX1 \block_reg[3][24]  ( .D(block_next[24]), .E(n1273), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFX1 \block_reg[7][24]  ( .D(block_next[24]), .E(n1239), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFX1 \block_reg[3][23]  ( .D(block_next[23]), .E(n1273), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFX1 \block_reg[7][23]  ( .D(block_next[23]), .E(n1239), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFX1 \block_reg[3][22]  ( .D(block_next[22]), .E(n1273), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFX1 \block_reg[7][22]  ( .D(block_next[22]), .E(n1239), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFX1 \block_reg[3][21]  ( .D(block_next[21]), .E(n1273), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFX1 \block_reg[7][21]  ( .D(block_next[21]), .E(n1239), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n1273), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFX1 \block_reg[7][20]  ( .D(block_next[20]), .E(n1239), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFX1 \block_reg[3][19]  ( .D(block_next[19]), .E(n1273), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFX1 \block_reg[7][19]  ( .D(block_next[19]), .E(n1239), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFX1 \block_reg[3][18]  ( .D(block_next[18]), .E(n1273), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFX1 \block_reg[7][18]  ( .D(block_next[18]), .E(n1239), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFX1 \block_reg[3][17]  ( .D(block_next[17]), .E(n1273), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFX1 \block_reg[7][17]  ( .D(block_next[17]), .E(n1239), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFX1 \block_reg[3][16]  ( .D(block_next[16]), .E(n1273), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFX1 \block_reg[7][16]  ( .D(block_next[16]), .E(n1239), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFX1 \block_reg[3][15]  ( .D(block_next[15]), .E(n1273), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFX1 \block_reg[7][15]  ( .D(block_next[15]), .E(n1239), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFX1 \block_reg[3][14]  ( .D(block_next[14]), .E(n1273), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFX1 \block_reg[7][14]  ( .D(block_next[14]), .E(n1239), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFX1 \block_reg[3][13]  ( .D(block_next[13]), .E(n1273), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFX1 \block_reg[7][13]  ( .D(block_next[13]), .E(n1239), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFX1 \block_reg[3][12]  ( .D(block_next[12]), .E(n1272), .CK(clk), .Q(
        \block[3][12] ) );
  EDFFX1 \block_reg[7][12]  ( .D(block_next[12]), .E(n1238), .CK(clk), .Q(
        \block[7][12] ) );
  EDFFX1 \block_reg[3][11]  ( .D(block_next[11]), .E(n1272), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFX1 \block_reg[7][11]  ( .D(block_next[11]), .E(n1238), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFX1 \block_reg[3][10]  ( .D(block_next[10]), .E(n1272), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFX1 \block_reg[7][10]  ( .D(block_next[10]), .E(n1238), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFX1 \block_reg[3][9]  ( .D(block_next[9]), .E(n1272), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFX1 \block_reg[7][9]  ( .D(block_next[9]), .E(n1238), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFX1 \block_reg[3][8]  ( .D(block_next[8]), .E(n1272), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFX1 \block_reg[7][8]  ( .D(block_next[8]), .E(n1238), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFX1 \block_reg[3][7]  ( .D(block_next[7]), .E(n1272), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFX1 \block_reg[7][7]  ( .D(block_next[7]), .E(n1238), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFX1 \block_reg[3][6]  ( .D(block_next[6]), .E(n1272), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFX1 \block_reg[7][6]  ( .D(block_next[6]), .E(n1238), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFX1 \block_reg[3][5]  ( .D(block_next[5]), .E(n1272), .CK(clk), .Q(
        \block[3][5] ) );
  EDFFX1 \block_reg[7][5]  ( .D(block_next[5]), .E(n1238), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFX1 \block_reg[3][4]  ( .D(block_next[4]), .E(n1272), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFX1 \block_reg[7][4]  ( .D(block_next[4]), .E(n1238), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFX1 \block_reg[3][3]  ( .D(block_next[3]), .E(n1272), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFX1 \block_reg[7][3]  ( .D(block_next[3]), .E(n1238), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFX1 \block_reg[3][2]  ( .D(block_next[2]), .E(n1272), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFX1 \block_reg[7][2]  ( .D(block_next[2]), .E(n1238), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFX1 \block_reg[3][1]  ( .D(block_next[1]), .E(n1272), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFX1 \block_reg[7][1]  ( .D(block_next[1]), .E(n1238), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFX1 \block_reg[3][0]  ( .D(block_next[0]), .E(n1272), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFX1 \block_reg[7][0]  ( .D(block_next[0]), .E(n1238), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFX1 \block_reg[1][127]  ( .D(block_next[127]), .E(n1288), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFX1 \block_reg[5][127]  ( .D(block_next[127]), .E(n1257), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFX1 \block_reg[1][126]  ( .D(block_next[126]), .E(n1288), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFX1 \block_reg[5][126]  ( .D(block_next[126]), .E(n1254), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFX1 \block_reg[1][125]  ( .D(block_next[125]), .E(n1288), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFX1 \block_reg[5][125]  ( .D(block_next[125]), .E(n1254), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFX1 \block_reg[1][124]  ( .D(block_next[124]), .E(n1292), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFX1 \block_reg[5][124]  ( .D(block_next[124]), .E(n1254), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFX1 \block_reg[1][123]  ( .D(block_next[123]), .E(n1290), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFX1 \block_reg[5][123]  ( .D(block_next[123]), .E(n1254), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFX1 \block_reg[1][122]  ( .D(block_next[122]), .E(n1289), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFX1 \block_reg[5][122]  ( .D(block_next[122]), .E(n1254), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFX1 \block_reg[1][121]  ( .D(block_next[121]), .E(n1291), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFX1 \block_reg[5][121]  ( .D(block_next[121]), .E(n1254), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFX1 \block_reg[1][120]  ( .D(block_next[120]), .E(n1291), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFX1 \block_reg[5][120]  ( .D(block_next[120]), .E(n1254), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFX1 \block_reg[1][119]  ( .D(block_next[119]), .E(n1293), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFX1 \block_reg[5][119]  ( .D(block_next[119]), .E(n1254), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFX1 \block_reg[1][118]  ( .D(block_next[118]), .E(n1294), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFX1 \block_reg[5][118]  ( .D(block_next[118]), .E(N962), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFX1 \block_reg[1][117]  ( .D(block_next[117]), .E(n1296), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFX1 \block_reg[5][117]  ( .D(block_next[117]), .E(N962), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFX1 \block_reg[1][116]  ( .D(block_next[116]), .E(n1294), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFX1 \block_reg[5][116]  ( .D(block_next[116]), .E(n1260), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFX1 \block_reg[1][115]  ( .D(block_next[115]), .E(n1296), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFX1 \block_reg[5][115]  ( .D(block_next[115]), .E(n1259), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFX1 \block_reg[1][114]  ( .D(block_next[114]), .E(n1295), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFX1 \block_reg[5][114]  ( .D(block_next[114]), .E(n1261), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFX1 \block_reg[1][113]  ( .D(block_next[113]), .E(n1288), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFX1 \block_reg[5][113]  ( .D(block_next[113]), .E(n1256), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFX1 \block_reg[1][112]  ( .D(block_next[112]), .E(n1288), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFX1 \block_reg[5][112]  ( .D(block_next[112]), .E(n1255), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFX1 \block_reg[1][111]  ( .D(block_next[111]), .E(n1292), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFX1 \block_reg[5][111]  ( .D(block_next[111]), .E(n1257), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFX1 \block_reg[1][110]  ( .D(block_next[110]), .E(n1290), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFX1 \block_reg[5][110]  ( .D(block_next[110]), .E(n1262), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFX1 \block_reg[1][109]  ( .D(block_next[109]), .E(n1289), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFX1 \block_reg[5][109]  ( .D(block_next[109]), .E(n1254), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFX1 \block_reg[1][108]  ( .D(block_next[108]), .E(n1291), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFX1 \block_reg[5][108]  ( .D(block_next[108]), .E(n1260), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFX1 \block_reg[1][107]  ( .D(block_next[107]), .E(n1293), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFX1 \block_reg[5][107]  ( .D(block_next[107]), .E(n1259), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFX1 \block_reg[1][106]  ( .D(block_next[106]), .E(n1293), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFX1 \block_reg[5][106]  ( .D(block_next[106]), .E(n1261), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFX1 \block_reg[1][105]  ( .D(block_next[105]), .E(n1294), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFX1 \block_reg[5][105]  ( .D(block_next[105]), .E(n1256), .CK(clk), .Q(
        \block[5][105] ) );
  EDFFX1 \block_reg[1][104]  ( .D(block_next[104]), .E(n1296), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFX1 \block_reg[5][104]  ( .D(block_next[104]), .E(n1255), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFX1 \block_reg[1][103]  ( .D(block_next[103]), .E(n1295), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFX1 \block_reg[5][103]  ( .D(block_next[103]), .E(n1262), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFX1 \block_reg[1][102]  ( .D(block_next[102]), .E(n1295), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFX1 \block_reg[5][102]  ( .D(block_next[102]), .E(n1262), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFX1 \block_reg[1][101]  ( .D(block_next[101]), .E(n1295), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFX1 \block_reg[5][101]  ( .D(block_next[101]), .E(n1262), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFX1 \block_reg[1][100]  ( .D(block_next[100]), .E(n1295), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFX1 \block_reg[5][100]  ( .D(block_next[100]), .E(n1262), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFX1 \block_reg[1][99]  ( .D(block_next[99]), .E(n1295), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFX1 \block_reg[5][99]  ( .D(block_next[99]), .E(n1262), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFX1 \block_reg[1][98]  ( .D(block_next[98]), .E(n1295), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFX1 \block_reg[5][98]  ( .D(block_next[98]), .E(n1262), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFX1 \block_reg[1][97]  ( .D(block_next[97]), .E(n1295), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFX1 \block_reg[5][97]  ( .D(block_next[97]), .E(n1262), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFX1 \block_reg[1][96]  ( .D(block_next[96]), .E(n1295), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFX1 \block_reg[5][96]  ( .D(block_next[96]), .E(n1262), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFX1 \block_reg[1][95]  ( .D(block_next[95]), .E(n1295), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFX1 \block_reg[5][95]  ( .D(block_next[95]), .E(n1262), .CK(clk), .Q(
        \block[5][95] ) );
  EDFFX1 \block_reg[1][94]  ( .D(block_next[94]), .E(n1295), .CK(clk), .Q(
        \block[1][94] ) );
  EDFFX1 \block_reg[5][94]  ( .D(block_next[94]), .E(n1262), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFX1 \block_reg[1][93]  ( .D(block_next[93]), .E(n1295), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFX1 \block_reg[5][93]  ( .D(block_next[93]), .E(n1262), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFX1 \block_reg[1][92]  ( .D(block_next[92]), .E(n1295), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFX1 \block_reg[5][92]  ( .D(block_next[92]), .E(n1262), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFX1 \block_reg[1][91]  ( .D(block_next[91]), .E(n1295), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFX1 \block_reg[5][91]  ( .D(block_next[91]), .E(n1262), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFX1 \block_reg[1][90]  ( .D(block_next[90]), .E(n1294), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFX1 \block_reg[5][90]  ( .D(block_next[90]), .E(n1261), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFX1 \block_reg[1][89]  ( .D(block_next[89]), .E(n1294), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFX1 \block_reg[5][89]  ( .D(block_next[89]), .E(n1261), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFX1 \block_reg[1][88]  ( .D(block_next[88]), .E(n1294), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFX1 \block_reg[5][88]  ( .D(block_next[88]), .E(n1261), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFX1 \block_reg[1][87]  ( .D(block_next[87]), .E(n1294), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFX1 \block_reg[5][87]  ( .D(block_next[87]), .E(n1261), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFX1 \block_reg[1][86]  ( .D(block_next[86]), .E(n1294), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFX1 \block_reg[5][86]  ( .D(block_next[86]), .E(n1261), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFX1 \block_reg[1][85]  ( .D(block_next[85]), .E(n1294), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFX1 \block_reg[5][85]  ( .D(block_next[85]), .E(n1261), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFX1 \block_reg[1][84]  ( .D(block_next[84]), .E(n1294), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFX1 \block_reg[5][84]  ( .D(block_next[84]), .E(n1261), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFX1 \block_reg[1][83]  ( .D(block_next[83]), .E(n1294), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFX1 \block_reg[5][83]  ( .D(block_next[83]), .E(n1261), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFX1 \block_reg[1][82]  ( .D(block_next[82]), .E(n1294), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFX1 \block_reg[5][82]  ( .D(block_next[82]), .E(n1261), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFX1 \block_reg[1][81]  ( .D(block_next[81]), .E(n1294), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFX1 \block_reg[5][81]  ( .D(block_next[81]), .E(n1261), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFX1 \block_reg[1][80]  ( .D(block_next[80]), .E(n1294), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFX1 \block_reg[5][80]  ( .D(block_next[80]), .E(n1261), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFX1 \block_reg[1][79]  ( .D(block_next[79]), .E(n1294), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFX1 \block_reg[5][79]  ( .D(block_next[79]), .E(n1261), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFX1 \block_reg[1][78]  ( .D(block_next[78]), .E(n1294), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFX1 \block_reg[5][78]  ( .D(block_next[78]), .E(n1261), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFX1 \block_reg[1][77]  ( .D(block_next[77]), .E(n1295), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFX1 \block_reg[5][77]  ( .D(block_next[77]), .E(n1260), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFX1 \block_reg[1][76]  ( .D(block_next[76]), .E(n1292), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFX1 \block_reg[5][76]  ( .D(block_next[76]), .E(n1260), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFX1 \block_reg[1][75]  ( .D(block_next[75]), .E(n1290), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFX1 \block_reg[5][75]  ( .D(block_next[75]), .E(n1260), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFX1 \block_reg[1][74]  ( .D(block_next[74]), .E(n1289), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFX1 \block_reg[5][74]  ( .D(block_next[74]), .E(n1260), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFX1 \block_reg[1][73]  ( .D(block_next[73]), .E(n1291), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFX1 \block_reg[5][73]  ( .D(block_next[73]), .E(n1260), .CK(clk), .Q(
        \block[5][73] ) );
  EDFFX1 \block_reg[1][72]  ( .D(block_next[72]), .E(n1293), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFX1 \block_reg[5][72]  ( .D(block_next[72]), .E(n1260), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFX1 \block_reg[1][71]  ( .D(block_next[71]), .E(n1294), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFX1 \block_reg[5][71]  ( .D(block_next[71]), .E(n1260), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFX1 \block_reg[1][70]  ( .D(block_next[70]), .E(n1296), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFX1 \block_reg[5][70]  ( .D(block_next[70]), .E(n1260), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFX1 \block_reg[1][69]  ( .D(block_next[69]), .E(n1295), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFX1 \block_reg[5][69]  ( .D(block_next[69]), .E(n1260), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFX1 \block_reg[1][68]  ( .D(block_next[68]), .E(n1288), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFX1 \block_reg[5][68]  ( .D(block_next[68]), .E(n1260), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFX1 \block_reg[1][67]  ( .D(block_next[67]), .E(n1292), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFX1 \block_reg[5][67]  ( .D(block_next[67]), .E(n1260), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFX1 \block_reg[1][66]  ( .D(block_next[66]), .E(n1290), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFX1 \block_reg[5][66]  ( .D(block_next[66]), .E(n1260), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFX1 \block_reg[1][65]  ( .D(block_next[65]), .E(n1289), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFX1 \block_reg[5][65]  ( .D(block_next[65]), .E(n1260), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFX1 \block_reg[1][64]  ( .D(block_next[64]), .E(n1293), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[5][64]  ( .D(block_next[64]), .E(n1259), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFX1 \block_reg[1][63]  ( .D(block_next[63]), .E(n1293), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFX1 \block_reg[5][63]  ( .D(block_next[63]), .E(n1259), .CK(clk), .Q(
        \block[5][63] ) );
  EDFFX1 \block_reg[1][62]  ( .D(block_next[62]), .E(n1293), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFX1 \block_reg[5][62]  ( .D(block_next[62]), .E(n1259), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFX1 \block_reg[1][61]  ( .D(block_next[61]), .E(n1293), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFX1 \block_reg[5][61]  ( .D(block_next[61]), .E(n1259), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFX1 \block_reg[1][60]  ( .D(block_next[60]), .E(n1293), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFX1 \block_reg[5][60]  ( .D(block_next[60]), .E(n1259), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFX1 \block_reg[1][59]  ( .D(block_next[59]), .E(n1293), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFX1 \block_reg[5][59]  ( .D(block_next[59]), .E(n1259), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFX1 \block_reg[1][58]  ( .D(block_next[58]), .E(n1293), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFX1 \block_reg[5][58]  ( .D(block_next[58]), .E(n1259), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFX1 \block_reg[1][57]  ( .D(block_next[57]), .E(n1293), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFX1 \block_reg[5][57]  ( .D(block_next[57]), .E(n1259), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFX1 \block_reg[1][56]  ( .D(block_next[56]), .E(n1293), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFX1 \block_reg[5][56]  ( .D(block_next[56]), .E(n1259), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFX1 \block_reg[1][55]  ( .D(block_next[55]), .E(n1293), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFX1 \block_reg[5][55]  ( .D(block_next[55]), .E(n1259), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFX1 \block_reg[1][54]  ( .D(block_next[54]), .E(n1293), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFX1 \block_reg[5][54]  ( .D(block_next[54]), .E(n1259), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n1293), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFX1 \block_reg[5][53]  ( .D(block_next[53]), .E(n1259), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n1293), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[5][52]  ( .D(block_next[52]), .E(n1259), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFX1 \block_reg[1][51]  ( .D(block_next[51]), .E(n1292), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFX1 \block_reg[5][51]  ( .D(block_next[51]), .E(n1258), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFX1 \block_reg[1][50]  ( .D(block_next[50]), .E(n1292), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFX1 \block_reg[5][50]  ( .D(block_next[50]), .E(n1258), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n1292), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[5][49]  ( .D(block_next[49]), .E(n1258), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFX1 \block_reg[1][48]  ( .D(block_next[48]), .E(n1292), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFX1 \block_reg[5][48]  ( .D(block_next[48]), .E(n1258), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFX1 \block_reg[1][47]  ( .D(block_next[47]), .E(n1292), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFX1 \block_reg[5][47]  ( .D(block_next[47]), .E(n1258), .CK(clk), .Q(
        \block[5][47] ) );
  EDFFX1 \block_reg[1][46]  ( .D(block_next[46]), .E(n1292), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFX1 \block_reg[5][46]  ( .D(block_next[46]), .E(n1258), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFX1 \block_reg[1][45]  ( .D(block_next[45]), .E(n1292), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFX1 \block_reg[5][45]  ( .D(block_next[45]), .E(n1258), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFX1 \block_reg[1][44]  ( .D(block_next[44]), .E(n1292), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFX1 \block_reg[5][44]  ( .D(block_next[44]), .E(n1258), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFX1 \block_reg[1][43]  ( .D(block_next[43]), .E(n1292), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFX1 \block_reg[5][43]  ( .D(block_next[43]), .E(n1258), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFX1 \block_reg[1][42]  ( .D(block_next[42]), .E(n1292), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFX1 \block_reg[5][42]  ( .D(block_next[42]), .E(n1258), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFX1 \block_reg[1][41]  ( .D(block_next[41]), .E(n1292), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n1258), .CK(clk), .Q(
        \block[5][41] ) );
  EDFFX1 \block_reg[1][40]  ( .D(block_next[40]), .E(n1292), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFX1 \block_reg[5][40]  ( .D(block_next[40]), .E(n1258), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFX1 \block_reg[1][39]  ( .D(block_next[39]), .E(n1292), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFX1 \block_reg[5][39]  ( .D(block_next[39]), .E(n1258), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFX1 \block_reg[1][38]  ( .D(block_next[38]), .E(n1291), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n1257), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFX1 \block_reg[1][37]  ( .D(block_next[37]), .E(n1291), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n1257), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFX1 \block_reg[1][36]  ( .D(block_next[36]), .E(n1291), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n1257), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(n1291), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFX1 \block_reg[5][35]  ( .D(block_next[35]), .E(n1257), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFX1 \block_reg[1][34]  ( .D(block_next[34]), .E(n1291), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFX1 \block_reg[5][34]  ( .D(block_next[34]), .E(n1257), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFX1 \block_reg[1][33]  ( .D(block_next[33]), .E(n1291), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFX1 \block_reg[5][33]  ( .D(block_next[33]), .E(n1257), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFX1 \block_reg[1][32]  ( .D(block_next[32]), .E(n1291), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n1257), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFX1 \block_reg[1][31]  ( .D(block_next[31]), .E(n1291), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFX1 \block_reg[5][31]  ( .D(block_next[31]), .E(n1257), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFX1 \block_reg[1][30]  ( .D(block_next[30]), .E(n1291), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFX1 \block_reg[5][30]  ( .D(block_next[30]), .E(n1257), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFX1 \block_reg[1][29]  ( .D(block_next[29]), .E(n1291), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFX1 \block_reg[5][29]  ( .D(block_next[29]), .E(n1257), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFX1 \block_reg[1][28]  ( .D(block_next[28]), .E(n1291), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFX1 \block_reg[5][28]  ( .D(block_next[28]), .E(n1257), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFX1 \block_reg[1][27]  ( .D(block_next[27]), .E(n1291), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFX1 \block_reg[5][27]  ( .D(block_next[27]), .E(n1257), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFX1 \block_reg[1][26]  ( .D(block_next[26]), .E(n1291), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFX1 \block_reg[5][26]  ( .D(block_next[26]), .E(n1257), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFX1 \block_reg[1][25]  ( .D(block_next[25]), .E(n1290), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFX1 \block_reg[5][25]  ( .D(block_next[25]), .E(n1256), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFX1 \block_reg[1][24]  ( .D(block_next[24]), .E(n1290), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFX1 \block_reg[5][24]  ( .D(block_next[24]), .E(n1256), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFX1 \block_reg[1][23]  ( .D(block_next[23]), .E(n1290), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFX1 \block_reg[5][23]  ( .D(block_next[23]), .E(n1256), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFX1 \block_reg[1][22]  ( .D(block_next[22]), .E(n1290), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFX1 \block_reg[5][22]  ( .D(block_next[22]), .E(n1256), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFX1 \block_reg[1][21]  ( .D(block_next[21]), .E(n1290), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFX1 \block_reg[5][21]  ( .D(block_next[21]), .E(n1256), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n1290), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFX1 \block_reg[5][20]  ( .D(block_next[20]), .E(n1256), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFX1 \block_reg[1][19]  ( .D(block_next[19]), .E(n1290), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFX1 \block_reg[5][19]  ( .D(block_next[19]), .E(n1256), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFX1 \block_reg[1][18]  ( .D(block_next[18]), .E(n1290), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFX1 \block_reg[5][18]  ( .D(block_next[18]), .E(n1256), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFX1 \block_reg[1][17]  ( .D(block_next[17]), .E(n1290), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFX1 \block_reg[5][17]  ( .D(block_next[17]), .E(n1256), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFX1 \block_reg[1][16]  ( .D(block_next[16]), .E(n1290), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFX1 \block_reg[5][16]  ( .D(block_next[16]), .E(n1256), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFX1 \block_reg[1][15]  ( .D(block_next[15]), .E(n1290), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFX1 \block_reg[5][15]  ( .D(block_next[15]), .E(n1256), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[1][14]  ( .D(block_next[14]), .E(n1290), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFX1 \block_reg[5][14]  ( .D(block_next[14]), .E(n1256), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFX1 \block_reg[1][13]  ( .D(block_next[13]), .E(n1290), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFX1 \block_reg[5][13]  ( .D(block_next[13]), .E(n1256), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFX1 \block_reg[1][12]  ( .D(block_next[12]), .E(n1289), .CK(clk), .Q(
        \block[1][12] ) );
  EDFFX1 \block_reg[5][12]  ( .D(block_next[12]), .E(n1255), .CK(clk), .Q(
        \block[5][12] ) );
  EDFFX1 \block_reg[1][11]  ( .D(block_next[11]), .E(n1289), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFX1 \block_reg[5][11]  ( .D(block_next[11]), .E(n1255), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFX1 \block_reg[1][10]  ( .D(block_next[10]), .E(n1289), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFX1 \block_reg[5][10]  ( .D(block_next[10]), .E(n1255), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFX1 \block_reg[1][9]  ( .D(block_next[9]), .E(n1289), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFX1 \block_reg[5][9]  ( .D(block_next[9]), .E(n1255), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFX1 \block_reg[1][8]  ( .D(block_next[8]), .E(n1289), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFX1 \block_reg[5][8]  ( .D(block_next[8]), .E(n1255), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFX1 \block_reg[1][7]  ( .D(block_next[7]), .E(n1289), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFX1 \block_reg[5][7]  ( .D(block_next[7]), .E(n1255), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFX1 \block_reg[1][6]  ( .D(block_next[6]), .E(n1289), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFX1 \block_reg[5][6]  ( .D(block_next[6]), .E(n1255), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFX1 \block_reg[1][5]  ( .D(block_next[5]), .E(n1289), .CK(clk), .Q(
        \block[1][5] ) );
  EDFFX1 \block_reg[5][5]  ( .D(block_next[5]), .E(n1255), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFX1 \block_reg[1][4]  ( .D(block_next[4]), .E(n1289), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFX1 \block_reg[5][4]  ( .D(block_next[4]), .E(n1255), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFX1 \block_reg[1][3]  ( .D(block_next[3]), .E(n1289), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFX1 \block_reg[5][3]  ( .D(block_next[3]), .E(n1255), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFX1 \block_reg[1][2]  ( .D(block_next[2]), .E(n1289), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFX1 \block_reg[5][2]  ( .D(block_next[2]), .E(n1255), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFX1 \block_reg[1][1]  ( .D(block_next[1]), .E(n1289), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFX1 \block_reg[5][1]  ( .D(block_next[1]), .E(n1255), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFX1 \block_reg[1][0]  ( .D(block_next[0]), .E(n1289), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFX1 \block_reg[5][0]  ( .D(block_next[0]), .E(n1255), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFX1 \block_reg[0][127]  ( .D(block_next[127]), .E(n1304), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFX1 \block_reg[4][127]  ( .D(block_next[127]), .E(n1270), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFX1 \block_reg[0][126]  ( .D(block_next[126]), .E(n1304), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFX1 \block_reg[4][126]  ( .D(block_next[126]), .E(n1270), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFX1 \block_reg[0][125]  ( .D(block_next[125]), .E(n1304), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFX1 \block_reg[4][125]  ( .D(block_next[125]), .E(n1270), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFX1 \block_reg[0][124]  ( .D(block_next[124]), .E(n1304), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFX1 \block_reg[4][124]  ( .D(block_next[124]), .E(n1270), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFX1 \block_reg[0][123]  ( .D(block_next[123]), .E(n1304), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFX1 \block_reg[4][123]  ( .D(block_next[123]), .E(n1270), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFX1 \block_reg[0][122]  ( .D(block_next[122]), .E(n1304), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFX1 \block_reg[4][122]  ( .D(block_next[122]), .E(n1270), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFX1 \block_reg[0][121]  ( .D(block_next[121]), .E(n1304), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFX1 \block_reg[4][121]  ( .D(block_next[121]), .E(n1270), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFX1 \block_reg[0][120]  ( .D(block_next[120]), .E(n1304), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFX1 \block_reg[4][120]  ( .D(block_next[120]), .E(n1270), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFX1 \block_reg[0][119]  ( .D(block_next[119]), .E(n1304), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFX1 \block_reg[4][119]  ( .D(block_next[119]), .E(n1270), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFX1 \block_reg[0][118]  ( .D(block_next[118]), .E(n1304), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFX1 \block_reg[4][118]  ( .D(block_next[118]), .E(n1270), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFX1 \block_reg[0][117]  ( .D(block_next[117]), .E(n1304), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFX1 \block_reg[4][117]  ( .D(block_next[117]), .E(n1270), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFX1 \block_reg[0][116]  ( .D(block_next[116]), .E(n1298), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFX1 \block_reg[4][116]  ( .D(block_next[116]), .E(n1268), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFX1 \block_reg[0][115]  ( .D(block_next[115]), .E(n1302), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFX1 \block_reg[4][115]  ( .D(block_next[115]), .E(n1267), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFX1 \block_reg[0][114]  ( .D(block_next[114]), .E(n1301), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFX1 \block_reg[4][114]  ( .D(block_next[114]), .E(n1266), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFX1 \block_reg[0][113]  ( .D(block_next[113]), .E(n1298), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFX1 \block_reg[4][113]  ( .D(block_next[113]), .E(n1268), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFX1 \block_reg[0][112]  ( .D(block_next[112]), .E(n1302), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFX1 \block_reg[4][112]  ( .D(block_next[112]), .E(n1267), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFX1 \block_reg[0][111]  ( .D(block_next[111]), .E(n1301), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFX1 \block_reg[4][111]  ( .D(block_next[111]), .E(n1266), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFX1 \block_reg[0][110]  ( .D(block_next[110]), .E(n1297), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFX1 \block_reg[4][110]  ( .D(block_next[110]), .E(n1268), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFX1 \block_reg[0][109]  ( .D(block_next[109]), .E(n1299), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFX1 \block_reg[4][109]  ( .D(block_next[109]), .E(n1263), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFX1 \block_reg[0][108]  ( .D(block_next[108]), .E(n1301), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFX1 \block_reg[4][108]  ( .D(block_next[108]), .E(n696), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFX1 \block_reg[0][107]  ( .D(block_next[107]), .E(n1300), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFX1 \block_reg[4][107]  ( .D(block_next[107]), .E(n696), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFX1 \block_reg[0][106]  ( .D(block_next[106]), .E(n1300), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFX1 \block_reg[4][106]  ( .D(block_next[106]), .E(n696), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFX1 \block_reg[0][105]  ( .D(block_next[105]), .E(n1300), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFX1 \block_reg[4][105]  ( .D(block_next[105]), .E(n696), .CK(clk), .Q(
        \block[4][105] ) );
  EDFFX1 \block_reg[0][104]  ( .D(block_next[104]), .E(n1300), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFX1 \block_reg[4][104]  ( .D(block_next[104]), .E(n696), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFX1 \block_reg[0][103]  ( .D(block_next[103]), .E(n1303), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFX1 \block_reg[4][103]  ( .D(block_next[103]), .E(n1269), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFX1 \block_reg[0][102]  ( .D(block_next[102]), .E(n1303), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFX1 \block_reg[4][102]  ( .D(block_next[102]), .E(n1269), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFX1 \block_reg[0][101]  ( .D(block_next[101]), .E(n1303), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFX1 \block_reg[4][101]  ( .D(block_next[101]), .E(n1269), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFX1 \block_reg[0][100]  ( .D(block_next[100]), .E(n1303), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFX1 \block_reg[4][100]  ( .D(block_next[100]), .E(n1269), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFX1 \block_reg[0][99]  ( .D(block_next[99]), .E(n1303), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFX1 \block_reg[4][99]  ( .D(block_next[99]), .E(n1269), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFX1 \block_reg[0][98]  ( .D(block_next[98]), .E(n1303), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFX1 \block_reg[4][98]  ( .D(block_next[98]), .E(n1269), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFX1 \block_reg[0][97]  ( .D(block_next[97]), .E(n1303), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFX1 \block_reg[4][97]  ( .D(block_next[97]), .E(n1269), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFX1 \block_reg[0][96]  ( .D(block_next[96]), .E(n1303), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFX1 \block_reg[4][96]  ( .D(block_next[96]), .E(n1269), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFX1 \block_reg[0][95]  ( .D(block_next[95]), .E(n1303), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFX1 \block_reg[4][95]  ( .D(block_next[95]), .E(n1269), .CK(clk), .Q(
        \block[4][95] ) );
  EDFFX1 \block_reg[0][94]  ( .D(block_next[94]), .E(n1303), .CK(clk), .Q(
        \block[0][94] ) );
  EDFFX1 \block_reg[4][94]  ( .D(block_next[94]), .E(n1269), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFX1 \block_reg[0][93]  ( .D(block_next[93]), .E(n1303), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFX1 \block_reg[4][93]  ( .D(block_next[93]), .E(n1269), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFX1 \block_reg[0][92]  ( .D(block_next[92]), .E(n1303), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFX1 \block_reg[4][92]  ( .D(block_next[92]), .E(n1269), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFX1 \block_reg[0][91]  ( .D(block_next[91]), .E(n1303), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFX1 \block_reg[4][91]  ( .D(block_next[91]), .E(n1269), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFX1 \block_reg[0][90]  ( .D(block_next[90]), .E(n1299), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFX1 \block_reg[4][90]  ( .D(block_next[90]), .E(n1268), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFX1 \block_reg[0][89]  ( .D(block_next[89]), .E(n1297), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFX1 \block_reg[4][89]  ( .D(block_next[89]), .E(n1268), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFX1 \block_reg[0][88]  ( .D(block_next[88]), .E(n1299), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFX1 \block_reg[4][88]  ( .D(block_next[88]), .E(n1268), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFX1 \block_reg[0][87]  ( .D(block_next[87]), .E(n698), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFX1 \block_reg[4][87]  ( .D(block_next[87]), .E(n1268), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFX1 \block_reg[0][86]  ( .D(block_next[86]), .E(n698), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFX1 \block_reg[4][86]  ( .D(block_next[86]), .E(n1268), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFX1 \block_reg[0][85]  ( .D(block_next[85]), .E(n698), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFX1 \block_reg[4][85]  ( .D(block_next[85]), .E(n1268), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFX1 \block_reg[0][84]  ( .D(block_next[84]), .E(n698), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFX1 \block_reg[4][84]  ( .D(block_next[84]), .E(n1268), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFX1 \block_reg[0][83]  ( .D(block_next[83]), .E(n698), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFX1 \block_reg[4][83]  ( .D(block_next[83]), .E(n1268), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFX1 \block_reg[0][82]  ( .D(block_next[82]), .E(n698), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFX1 \block_reg[4][82]  ( .D(block_next[82]), .E(n1268), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFX1 \block_reg[0][81]  ( .D(block_next[81]), .E(n1298), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFX1 \block_reg[4][81]  ( .D(block_next[81]), .E(n1268), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFX1 \block_reg[0][80]  ( .D(block_next[80]), .E(n1302), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFX1 \block_reg[4][80]  ( .D(block_next[80]), .E(n1268), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFX1 \block_reg[0][79]  ( .D(block_next[79]), .E(n1297), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFX1 \block_reg[4][79]  ( .D(block_next[79]), .E(n1268), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFX1 \block_reg[0][78]  ( .D(block_next[78]), .E(n1299), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFX1 \block_reg[4][78]  ( .D(block_next[78]), .E(n1268), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFX1 \block_reg[0][77]  ( .D(block_next[77]), .E(n1302), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFX1 \block_reg[4][77]  ( .D(block_next[77]), .E(n1267), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFX1 \block_reg[0][76]  ( .D(block_next[76]), .E(n1302), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFX1 \block_reg[4][76]  ( .D(block_next[76]), .E(n1267), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFX1 \block_reg[0][75]  ( .D(block_next[75]), .E(n1302), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFX1 \block_reg[4][75]  ( .D(block_next[75]), .E(n1267), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFX1 \block_reg[0][74]  ( .D(block_next[74]), .E(n1302), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFX1 \block_reg[4][74]  ( .D(block_next[74]), .E(n1267), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFX1 \block_reg[0][73]  ( .D(block_next[73]), .E(n1302), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFX1 \block_reg[4][73]  ( .D(block_next[73]), .E(n1267), .CK(clk), .Q(
        \block[4][73] ) );
  EDFFX1 \block_reg[0][72]  ( .D(block_next[72]), .E(n1302), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFX1 \block_reg[4][72]  ( .D(block_next[72]), .E(n1267), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFX1 \block_reg[0][71]  ( .D(block_next[71]), .E(n1302), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFX1 \block_reg[4][71]  ( .D(block_next[71]), .E(n1267), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFX1 \block_reg[0][70]  ( .D(block_next[70]), .E(n1302), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFX1 \block_reg[4][70]  ( .D(block_next[70]), .E(n1267), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFX1 \block_reg[0][69]  ( .D(block_next[69]), .E(n1302), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFX1 \block_reg[4][69]  ( .D(block_next[69]), .E(n1267), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFX1 \block_reg[0][68]  ( .D(block_next[68]), .E(n1302), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFX1 \block_reg[4][68]  ( .D(block_next[68]), .E(n1267), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFX1 \block_reg[0][67]  ( .D(block_next[67]), .E(n1302), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFX1 \block_reg[4][67]  ( .D(block_next[67]), .E(n1267), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFX1 \block_reg[0][66]  ( .D(block_next[66]), .E(n1302), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFX1 \block_reg[4][66]  ( .D(block_next[66]), .E(n1267), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFX1 \block_reg[0][65]  ( .D(block_next[65]), .E(n1302), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFX1 \block_reg[4][65]  ( .D(block_next[65]), .E(n1267), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFX1 \block_reg[0][64]  ( .D(block_next[64]), .E(n1301), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[4][64]  ( .D(block_next[64]), .E(n1266), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFX1 \block_reg[0][63]  ( .D(block_next[63]), .E(n1301), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFX1 \block_reg[4][63]  ( .D(block_next[63]), .E(n1266), .CK(clk), .Q(
        \block[4][63] ) );
  EDFFX1 \block_reg[0][62]  ( .D(block_next[62]), .E(n1301), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFX1 \block_reg[4][62]  ( .D(block_next[62]), .E(n1266), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFX1 \block_reg[0][61]  ( .D(block_next[61]), .E(n1301), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFX1 \block_reg[4][61]  ( .D(block_next[61]), .E(n1266), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFX1 \block_reg[0][60]  ( .D(block_next[60]), .E(n1301), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFX1 \block_reg[4][60]  ( .D(block_next[60]), .E(n1266), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFX1 \block_reg[0][59]  ( .D(block_next[59]), .E(n1301), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFX1 \block_reg[4][59]  ( .D(block_next[59]), .E(n1266), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFX1 \block_reg[0][58]  ( .D(block_next[58]), .E(n1301), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFX1 \block_reg[4][58]  ( .D(block_next[58]), .E(n1266), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFX1 \block_reg[0][57]  ( .D(block_next[57]), .E(n1301), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFX1 \block_reg[4][57]  ( .D(block_next[57]), .E(n1266), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFX1 \block_reg[0][56]  ( .D(block_next[56]), .E(n1301), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFX1 \block_reg[4][56]  ( .D(block_next[56]), .E(n1266), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFX1 \block_reg[0][55]  ( .D(block_next[55]), .E(n1301), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFX1 \block_reg[4][55]  ( .D(block_next[55]), .E(n1266), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFX1 \block_reg[0][54]  ( .D(block_next[54]), .E(n1301), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFX1 \block_reg[4][54]  ( .D(block_next[54]), .E(n1266), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n1301), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n1266), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n1301), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n1266), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[0][51]  ( .D(block_next[51]), .E(n1300), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFX1 \block_reg[4][51]  ( .D(block_next[51]), .E(n1265), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFX1 \block_reg[0][50]  ( .D(block_next[50]), .E(n1300), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFX1 \block_reg[4][50]  ( .D(block_next[50]), .E(n1265), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n1300), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n1265), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[0][48]  ( .D(block_next[48]), .E(n1300), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFX1 \block_reg[4][48]  ( .D(block_next[48]), .E(n1265), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFX1 \block_reg[0][47]  ( .D(block_next[47]), .E(n1300), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFX1 \block_reg[4][47]  ( .D(block_next[47]), .E(n1265), .CK(clk), .Q(
        \block[4][47] ) );
  EDFFX1 \block_reg[0][46]  ( .D(block_next[46]), .E(n1300), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFX1 \block_reg[4][46]  ( .D(block_next[46]), .E(n1265), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFX1 \block_reg[0][45]  ( .D(block_next[45]), .E(n1300), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFX1 \block_reg[4][45]  ( .D(block_next[45]), .E(n1265), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFX1 \block_reg[0][44]  ( .D(block_next[44]), .E(n1300), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFX1 \block_reg[4][44]  ( .D(block_next[44]), .E(n1265), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFX1 \block_reg[0][43]  ( .D(block_next[43]), .E(n1300), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFX1 \block_reg[4][43]  ( .D(block_next[43]), .E(n1265), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFX1 \block_reg[0][42]  ( .D(block_next[42]), .E(n1300), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFX1 \block_reg[4][42]  ( .D(block_next[42]), .E(n1265), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n1300), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n1265), .CK(clk), .Q(
        \block[4][41] ) );
  EDFFX1 \block_reg[0][40]  ( .D(block_next[40]), .E(n1300), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFX1 \block_reg[4][40]  ( .D(block_next[40]), .E(n1265), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFX1 \block_reg[0][39]  ( .D(block_next[39]), .E(n1300), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFX1 \block_reg[4][39]  ( .D(block_next[39]), .E(n1265), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n1299), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n1264), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n1299), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n1264), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n1299), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n1264), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n1299), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n1264), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFX1 \block_reg[0][34]  ( .D(block_next[34]), .E(n1299), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFX1 \block_reg[4][34]  ( .D(block_next[34]), .E(n1264), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFX1 \block_reg[0][33]  ( .D(block_next[33]), .E(n1299), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFX1 \block_reg[4][33]  ( .D(block_next[33]), .E(n1264), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n1299), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n1264), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[0][31]  ( .D(block_next[31]), .E(n1299), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFX1 \block_reg[4][31]  ( .D(block_next[31]), .E(n1264), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFX1 \block_reg[0][30]  ( .D(block_next[30]), .E(n1299), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFX1 \block_reg[4][30]  ( .D(block_next[30]), .E(n1264), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFX1 \block_reg[0][29]  ( .D(block_next[29]), .E(n1299), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFX1 \block_reg[4][29]  ( .D(block_next[29]), .E(n696), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFX1 \block_reg[0][28]  ( .D(block_next[28]), .E(n1299), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFX1 \block_reg[4][28]  ( .D(block_next[28]), .E(n696), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFX1 \block_reg[0][27]  ( .D(block_next[27]), .E(n1299), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFX1 \block_reg[4][27]  ( .D(block_next[27]), .E(n696), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFX1 \block_reg[0][26]  ( .D(block_next[26]), .E(n1299), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFX1 \block_reg[4][26]  ( .D(block_next[26]), .E(n696), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFX1 \block_reg[0][25]  ( .D(block_next[25]), .E(n1298), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFX1 \block_reg[4][25]  ( .D(block_next[25]), .E(n1264), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFX1 \block_reg[0][24]  ( .D(block_next[24]), .E(n1298), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFX1 \block_reg[4][24]  ( .D(block_next[24]), .E(n1264), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFX1 \block_reg[0][23]  ( .D(block_next[23]), .E(n1298), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFX1 \block_reg[4][23]  ( .D(block_next[23]), .E(n1267), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFX1 \block_reg[0][22]  ( .D(block_next[22]), .E(n1298), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFX1 \block_reg[4][22]  ( .D(block_next[22]), .E(n1266), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFX1 \block_reg[0][21]  ( .D(block_next[21]), .E(n1298), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFX1 \block_reg[4][21]  ( .D(block_next[21]), .E(n1268), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n1298), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n1263), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFX1 \block_reg[0][19]  ( .D(block_next[19]), .E(n1298), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFX1 \block_reg[4][19]  ( .D(block_next[19]), .E(n1269), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFX1 \block_reg[0][18]  ( .D(block_next[18]), .E(n1298), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFX1 \block_reg[4][18]  ( .D(block_next[18]), .E(n1270), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFX1 \block_reg[0][17]  ( .D(block_next[17]), .E(n1298), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFX1 \block_reg[4][17]  ( .D(block_next[17]), .E(n1265), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFX1 \block_reg[0][16]  ( .D(block_next[16]), .E(n1298), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFX1 \block_reg[4][16]  ( .D(block_next[16]), .E(n1269), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFX1 \block_reg[0][15]  ( .D(block_next[15]), .E(n1298), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFX1 \block_reg[4][15]  ( .D(block_next[15]), .E(n1270), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFX1 \block_reg[0][14]  ( .D(block_next[14]), .E(n1298), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFX1 \block_reg[4][14]  ( .D(block_next[14]), .E(n1265), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFX1 \block_reg[0][13]  ( .D(block_next[13]), .E(n1298), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFX1 \block_reg[4][13]  ( .D(block_next[13]), .E(n1269), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFX1 \block_reg[0][12]  ( .D(block_next[12]), .E(n1297), .CK(clk), .Q(
        \block[0][12] ) );
  EDFFX1 \block_reg[4][12]  ( .D(block_next[12]), .E(n1263), .CK(clk), .Q(
        \block[4][12] ) );
  EDFFX1 \block_reg[0][11]  ( .D(block_next[11]), .E(n1297), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFX1 \block_reg[4][11]  ( .D(block_next[11]), .E(n1263), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFX1 \block_reg[0][10]  ( .D(block_next[10]), .E(n1297), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFX1 \block_reg[4][10]  ( .D(block_next[10]), .E(n1263), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFX1 \block_reg[0][9]  ( .D(block_next[9]), .E(n1297), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFX1 \block_reg[4][9]  ( .D(block_next[9]), .E(n1263), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFX1 \block_reg[0][8]  ( .D(block_next[8]), .E(n1297), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFX1 \block_reg[4][8]  ( .D(block_next[8]), .E(n1263), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFX1 \block_reg[0][7]  ( .D(block_next[7]), .E(n1297), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFX1 \block_reg[4][7]  ( .D(block_next[7]), .E(n1263), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFX1 \block_reg[0][6]  ( .D(block_next[6]), .E(n1297), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFX1 \block_reg[4][6]  ( .D(block_next[6]), .E(n1263), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFX1 \block_reg[0][5]  ( .D(block_next[5]), .E(n1297), .CK(clk), .Q(
        \block[0][5] ) );
  EDFFX1 \block_reg[4][5]  ( .D(block_next[5]), .E(n1263), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFX1 \block_reg[0][4]  ( .D(block_next[4]), .E(n1297), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFX1 \block_reg[4][4]  ( .D(block_next[4]), .E(n1263), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFX1 \block_reg[0][3]  ( .D(block_next[3]), .E(n1297), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFX1 \block_reg[4][3]  ( .D(block_next[3]), .E(n1263), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFX1 \block_reg[0][2]  ( .D(block_next[2]), .E(n1297), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFX1 \block_reg[4][2]  ( .D(block_next[2]), .E(n1263), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFX1 \block_reg[0][1]  ( .D(block_next[1]), .E(n1297), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFX1 \block_reg[4][1]  ( .D(block_next[1]), .E(n1263), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFX1 \block_reg[0][0]  ( .D(block_next[0]), .E(n1297), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFX1 \block_reg[4][0]  ( .D(block_next[0]), .E(n1267), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFX1 \block_reg[2][127]  ( .D(block_next[127]), .E(n1287), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFX1 \block_reg[6][127]  ( .D(block_next[127]), .E(n1253), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFX1 \block_reg[2][126]  ( .D(block_next[126]), .E(n1287), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFX1 \block_reg[6][126]  ( .D(block_next[126]), .E(n1253), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFX1 \block_reg[2][125]  ( .D(block_next[125]), .E(n1287), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFX1 \block_reg[6][125]  ( .D(block_next[125]), .E(n1253), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFX1 \block_reg[2][124]  ( .D(block_next[124]), .E(n1287), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFX1 \block_reg[6][124]  ( .D(block_next[124]), .E(n1253), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFX1 \block_reg[2][123]  ( .D(block_next[123]), .E(n1287), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFX1 \block_reg[6][123]  ( .D(block_next[123]), .E(n1253), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFX1 \block_reg[2][122]  ( .D(block_next[122]), .E(n1287), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFX1 \block_reg[6][122]  ( .D(block_next[122]), .E(n1253), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFX1 \block_reg[2][121]  ( .D(block_next[121]), .E(n1287), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFX1 \block_reg[6][121]  ( .D(block_next[121]), .E(n1253), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFX1 \block_reg[2][120]  ( .D(block_next[120]), .E(n1287), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFX1 \block_reg[6][120]  ( .D(block_next[120]), .E(n1253), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFX1 \block_reg[2][119]  ( .D(block_next[119]), .E(n1287), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFX1 \block_reg[6][119]  ( .D(block_next[119]), .E(n1253), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFX1 \block_reg[2][118]  ( .D(block_next[118]), .E(n1287), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFX1 \block_reg[6][118]  ( .D(block_next[118]), .E(n1253), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFX1 \block_reg[2][117]  ( .D(block_next[117]), .E(n1287), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFX1 \block_reg[6][117]  ( .D(block_next[117]), .E(n1253), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFX1 \block_reg[2][116]  ( .D(block_next[116]), .E(n1282), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFX1 \block_reg[6][116]  ( .D(block_next[116]), .E(n1251), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFX1 \block_reg[2][115]  ( .D(block_next[115]), .E(n1280), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFX1 \block_reg[6][115]  ( .D(block_next[115]), .E(n1250), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFX1 \block_reg[2][114]  ( .D(block_next[114]), .E(n1282), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFX1 \block_reg[6][114]  ( .D(block_next[114]), .E(n1249), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFX1 \block_reg[2][113]  ( .D(block_next[113]), .E(n697), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFX1 \block_reg[6][113]  ( .D(block_next[113]), .E(n1251), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFX1 \block_reg[2][112]  ( .D(block_next[112]), .E(n697), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFX1 \block_reg[6][112]  ( .D(block_next[112]), .E(n1250), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFX1 \block_reg[2][111]  ( .D(block_next[111]), .E(n697), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFX1 \block_reg[6][111]  ( .D(block_next[111]), .E(n1249), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFX1 \block_reg[2][110]  ( .D(block_next[110]), .E(n697), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFX1 \block_reg[6][110]  ( .D(block_next[110]), .E(n1251), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFX1 \block_reg[2][109]  ( .D(block_next[109]), .E(n697), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFX1 \block_reg[6][109]  ( .D(block_next[109]), .E(n1246), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFX1 \block_reg[2][108]  ( .D(block_next[108]), .E(n697), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFX1 \block_reg[6][108]  ( .D(block_next[108]), .E(n695), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFX1 \block_reg[2][107]  ( .D(block_next[107]), .E(n1281), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFX1 \block_reg[6][107]  ( .D(block_next[107]), .E(n695), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFX1 \block_reg[2][106]  ( .D(block_next[106]), .E(n1285), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFX1 \block_reg[6][106]  ( .D(block_next[106]), .E(n695), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFX1 \block_reg[2][105]  ( .D(block_next[105]), .E(n1280), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFX1 \block_reg[6][105]  ( .D(block_next[105]), .E(n695), .CK(clk), .Q(
        \block[6][105] ) );
  EDFFX1 \block_reg[2][104]  ( .D(block_next[104]), .E(n1282), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFX1 \block_reg[6][104]  ( .D(block_next[104]), .E(n695), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFX1 \block_reg[2][103]  ( .D(block_next[103]), .E(n1286), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFX1 \block_reg[6][103]  ( .D(block_next[103]), .E(n1252), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFX1 \block_reg[2][102]  ( .D(block_next[102]), .E(n1286), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFX1 \block_reg[6][102]  ( .D(block_next[102]), .E(n1252), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFX1 \block_reg[2][101]  ( .D(block_next[101]), .E(n1286), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFX1 \block_reg[6][101]  ( .D(block_next[101]), .E(n1252), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFX1 \block_reg[2][100]  ( .D(block_next[100]), .E(n1286), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFX1 \block_reg[6][100]  ( .D(block_next[100]), .E(n1252), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFX1 \block_reg[2][99]  ( .D(block_next[99]), .E(n1286), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFX1 \block_reg[6][99]  ( .D(block_next[99]), .E(n1252), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFX1 \block_reg[2][98]  ( .D(block_next[98]), .E(n1286), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFX1 \block_reg[6][98]  ( .D(block_next[98]), .E(n1252), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFX1 \block_reg[2][97]  ( .D(block_next[97]), .E(n1286), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFX1 \block_reg[6][97]  ( .D(block_next[97]), .E(n1252), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFX1 \block_reg[2][96]  ( .D(block_next[96]), .E(n1286), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFX1 \block_reg[6][96]  ( .D(block_next[96]), .E(n1252), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFX1 \block_reg[2][95]  ( .D(block_next[95]), .E(n1286), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFX1 \block_reg[6][95]  ( .D(block_next[95]), .E(n1252), .CK(clk), .Q(
        \block[6][95] ) );
  EDFFX1 \block_reg[2][94]  ( .D(block_next[94]), .E(n1286), .CK(clk), .Q(
        \block[2][94] ) );
  EDFFX1 \block_reg[6][94]  ( .D(block_next[94]), .E(n1252), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFX1 \block_reg[2][93]  ( .D(block_next[93]), .E(n1286), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFX1 \block_reg[6][93]  ( .D(block_next[93]), .E(n1252), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFX1 \block_reg[2][92]  ( .D(block_next[92]), .E(n1286), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFX1 \block_reg[6][92]  ( .D(block_next[92]), .E(n1252), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFX1 \block_reg[2][91]  ( .D(block_next[91]), .E(n1286), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFX1 \block_reg[6][91]  ( .D(block_next[91]), .E(n1252), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFX1 \block_reg[2][90]  ( .D(block_next[90]), .E(n1283), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFX1 \block_reg[6][90]  ( .D(block_next[90]), .E(n1251), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFX1 \block_reg[2][89]  ( .D(block_next[89]), .E(n1281), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFX1 \block_reg[6][89]  ( .D(block_next[89]), .E(n1251), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFX1 \block_reg[2][88]  ( .D(block_next[88]), .E(n1285), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFX1 \block_reg[6][88]  ( .D(block_next[88]), .E(n1251), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFX1 \block_reg[2][87]  ( .D(block_next[87]), .E(n1286), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFX1 \block_reg[6][87]  ( .D(block_next[87]), .E(n1251), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFX1 \block_reg[2][86]  ( .D(block_next[86]), .E(n1283), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFX1 \block_reg[6][86]  ( .D(block_next[86]), .E(n1251), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFX1 \block_reg[2][85]  ( .D(block_next[85]), .E(n1280), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFX1 \block_reg[6][85]  ( .D(block_next[85]), .E(n1251), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFX1 \block_reg[2][84]  ( .D(block_next[84]), .E(n1282), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFX1 \block_reg[6][84]  ( .D(block_next[84]), .E(n1251), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFX1 \block_reg[2][83]  ( .D(block_next[83]), .E(n1284), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFX1 \block_reg[6][83]  ( .D(block_next[83]), .E(n1251), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFX1 \block_reg[2][82]  ( .D(block_next[82]), .E(n1284), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFX1 \block_reg[6][82]  ( .D(block_next[82]), .E(n1251), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFX1 \block_reg[2][81]  ( .D(block_next[81]), .E(n1284), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFX1 \block_reg[6][81]  ( .D(block_next[81]), .E(n1251), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFX1 \block_reg[2][80]  ( .D(block_next[80]), .E(n1284), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFX1 \block_reg[6][80]  ( .D(block_next[80]), .E(n1251), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFX1 \block_reg[2][79]  ( .D(block_next[79]), .E(n1284), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFX1 \block_reg[6][79]  ( .D(block_next[79]), .E(n1251), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFX1 \block_reg[2][78]  ( .D(block_next[78]), .E(n1284), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFX1 \block_reg[6][78]  ( .D(block_next[78]), .E(n1251), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFX1 \block_reg[2][77]  ( .D(block_next[77]), .E(n1285), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFX1 \block_reg[6][77]  ( .D(block_next[77]), .E(n1250), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFX1 \block_reg[2][76]  ( .D(block_next[76]), .E(n1285), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFX1 \block_reg[6][76]  ( .D(block_next[76]), .E(n1250), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFX1 \block_reg[2][75]  ( .D(block_next[75]), .E(n1285), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFX1 \block_reg[6][75]  ( .D(block_next[75]), .E(n1250), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFX1 \block_reg[2][74]  ( .D(block_next[74]), .E(n1285), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFX1 \block_reg[6][74]  ( .D(block_next[74]), .E(n1250), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFX1 \block_reg[2][73]  ( .D(block_next[73]), .E(n1285), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFX1 \block_reg[6][73]  ( .D(block_next[73]), .E(n1250), .CK(clk), .Q(
        \block[6][73] ) );
  EDFFX1 \block_reg[2][72]  ( .D(block_next[72]), .E(n1285), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFX1 \block_reg[6][72]  ( .D(block_next[72]), .E(n1250), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFX1 \block_reg[2][71]  ( .D(block_next[71]), .E(n1285), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFX1 \block_reg[6][71]  ( .D(block_next[71]), .E(n1250), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFX1 \block_reg[2][70]  ( .D(block_next[70]), .E(n1285), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFX1 \block_reg[6][70]  ( .D(block_next[70]), .E(n1250), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFX1 \block_reg[2][69]  ( .D(block_next[69]), .E(n1285), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFX1 \block_reg[6][69]  ( .D(block_next[69]), .E(n1250), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFX1 \block_reg[2][68]  ( .D(block_next[68]), .E(n1285), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFX1 \block_reg[6][68]  ( .D(block_next[68]), .E(n1250), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFX1 \block_reg[2][67]  ( .D(block_next[67]), .E(n1285), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFX1 \block_reg[6][67]  ( .D(block_next[67]), .E(n1250), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFX1 \block_reg[2][66]  ( .D(block_next[66]), .E(n1285), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFX1 \block_reg[6][66]  ( .D(block_next[66]), .E(n1250), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFX1 \block_reg[2][65]  ( .D(block_next[65]), .E(n1285), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFX1 \block_reg[6][65]  ( .D(block_next[65]), .E(n1250), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFX1 \block_reg[2][64]  ( .D(block_next[64]), .E(n1284), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFX1 \block_reg[6][64]  ( .D(block_next[64]), .E(n1249), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFX1 \block_reg[2][63]  ( .D(block_next[63]), .E(n1284), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFX1 \block_reg[6][63]  ( .D(block_next[63]), .E(n1249), .CK(clk), .Q(
        \block[6][63] ) );
  EDFFX1 \block_reg[2][62]  ( .D(block_next[62]), .E(n1284), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFX1 \block_reg[6][62]  ( .D(block_next[62]), .E(n1249), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFX1 \block_reg[2][61]  ( .D(block_next[61]), .E(n1284), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFX1 \block_reg[6][61]  ( .D(block_next[61]), .E(n1249), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFX1 \block_reg[2][60]  ( .D(block_next[60]), .E(n1284), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFX1 \block_reg[6][60]  ( .D(block_next[60]), .E(n1249), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFX1 \block_reg[2][59]  ( .D(block_next[59]), .E(n1284), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFX1 \block_reg[6][59]  ( .D(block_next[59]), .E(n1249), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFX1 \block_reg[2][58]  ( .D(block_next[58]), .E(n1284), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFX1 \block_reg[6][58]  ( .D(block_next[58]), .E(n1249), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFX1 \block_reg[2][57]  ( .D(block_next[57]), .E(n1284), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFX1 \block_reg[6][57]  ( .D(block_next[57]), .E(n1249), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFX1 \block_reg[2][56]  ( .D(block_next[56]), .E(n1284), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFX1 \block_reg[6][56]  ( .D(block_next[56]), .E(n1249), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFX1 \block_reg[2][55]  ( .D(block_next[55]), .E(n1284), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFX1 \block_reg[6][55]  ( .D(block_next[55]), .E(n1249), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFX1 \block_reg[2][54]  ( .D(block_next[54]), .E(n1284), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFX1 \block_reg[6][54]  ( .D(block_next[54]), .E(n1249), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFX1 \block_reg[2][53]  ( .D(block_next[53]), .E(n1284), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n1249), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFX1 \block_reg[2][52]  ( .D(block_next[52]), .E(n1284), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n1249), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[2][51]  ( .D(block_next[51]), .E(n1283), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFX1 \block_reg[6][51]  ( .D(block_next[51]), .E(n1248), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFX1 \block_reg[2][50]  ( .D(block_next[50]), .E(n1283), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFX1 \block_reg[6][50]  ( .D(block_next[50]), .E(n1248), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFX1 \block_reg[2][49]  ( .D(block_next[49]), .E(n1283), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFX1 \block_reg[6][49]  ( .D(block_next[49]), .E(n1248), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFX1 \block_reg[2][48]  ( .D(block_next[48]), .E(n1283), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFX1 \block_reg[6][48]  ( .D(block_next[48]), .E(n1248), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFX1 \block_reg[2][47]  ( .D(block_next[47]), .E(n1283), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFX1 \block_reg[6][47]  ( .D(block_next[47]), .E(n1248), .CK(clk), .Q(
        \block[6][47] ) );
  EDFFX1 \block_reg[2][46]  ( .D(block_next[46]), .E(n1283), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFX1 \block_reg[6][46]  ( .D(block_next[46]), .E(n1248), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFX1 \block_reg[2][45]  ( .D(block_next[45]), .E(n1283), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFX1 \block_reg[6][45]  ( .D(block_next[45]), .E(n1248), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFX1 \block_reg[2][44]  ( .D(block_next[44]), .E(n1283), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFX1 \block_reg[6][44]  ( .D(block_next[44]), .E(n1248), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFX1 \block_reg[2][43]  ( .D(block_next[43]), .E(n1283), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFX1 \block_reg[6][43]  ( .D(block_next[43]), .E(n1248), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFX1 \block_reg[2][42]  ( .D(block_next[42]), .E(n1283), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFX1 \block_reg[6][42]  ( .D(block_next[42]), .E(n1248), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFX1 \block_reg[2][41]  ( .D(block_next[41]), .E(n1283), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n1248), .CK(clk), .Q(
        \block[6][41] ) );
  EDFFX1 \block_reg[2][40]  ( .D(block_next[40]), .E(n1283), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFX1 \block_reg[6][40]  ( .D(block_next[40]), .E(n1248), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFX1 \block_reg[2][39]  ( .D(block_next[39]), .E(n1283), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFX1 \block_reg[6][39]  ( .D(block_next[39]), .E(n1248), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFX1 \block_reg[2][38]  ( .D(block_next[38]), .E(n1282), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n1247), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[2][37]  ( .D(block_next[37]), .E(n1282), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n1247), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[2][36]  ( .D(block_next[36]), .E(n1282), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n1247), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFX1 \block_reg[2][35]  ( .D(block_next[35]), .E(n1282), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n1247), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFX1 \block_reg[2][34]  ( .D(block_next[34]), .E(n1282), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFX1 \block_reg[6][34]  ( .D(block_next[34]), .E(n1247), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFX1 \block_reg[2][33]  ( .D(block_next[33]), .E(n1282), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFX1 \block_reg[6][33]  ( .D(block_next[33]), .E(n1247), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFX1 \block_reg[2][32]  ( .D(block_next[32]), .E(n1282), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n1247), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[2][31]  ( .D(block_next[31]), .E(n1282), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFX1 \block_reg[6][31]  ( .D(block_next[31]), .E(n1247), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFX1 \block_reg[2][30]  ( .D(block_next[30]), .E(n1282), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFX1 \block_reg[6][30]  ( .D(block_next[30]), .E(n1247), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFX1 \block_reg[2][29]  ( .D(block_next[29]), .E(n1282), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFX1 \block_reg[6][29]  ( .D(block_next[29]), .E(n695), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFX1 \block_reg[2][28]  ( .D(block_next[28]), .E(n1282), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFX1 \block_reg[6][28]  ( .D(block_next[28]), .E(n695), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFX1 \block_reg[2][27]  ( .D(block_next[27]), .E(n1282), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFX1 \block_reg[6][27]  ( .D(block_next[27]), .E(n695), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFX1 \block_reg[2][26]  ( .D(block_next[26]), .E(n1282), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFX1 \block_reg[6][26]  ( .D(block_next[26]), .E(n695), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFX1 \block_reg[2][25]  ( .D(block_next[25]), .E(n1281), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFX1 \block_reg[6][25]  ( .D(block_next[25]), .E(n1247), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFX1 \block_reg[2][24]  ( .D(block_next[24]), .E(n1281), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFX1 \block_reg[6][24]  ( .D(block_next[24]), .E(n1247), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFX1 \block_reg[2][23]  ( .D(block_next[23]), .E(n1281), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFX1 \block_reg[6][23]  ( .D(block_next[23]), .E(n1250), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFX1 \block_reg[2][22]  ( .D(block_next[22]), .E(n1281), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFX1 \block_reg[6][22]  ( .D(block_next[22]), .E(n1249), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFX1 \block_reg[2][21]  ( .D(block_next[21]), .E(n1281), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFX1 \block_reg[6][21]  ( .D(block_next[21]), .E(n1251), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFX1 \block_reg[2][20]  ( .D(block_next[20]), .E(n1281), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n1246), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFX1 \block_reg[2][19]  ( .D(block_next[19]), .E(n1281), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFX1 \block_reg[6][19]  ( .D(block_next[19]), .E(n1252), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFX1 \block_reg[2][18]  ( .D(block_next[18]), .E(n1281), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFX1 \block_reg[6][18]  ( .D(block_next[18]), .E(n1253), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFX1 \block_reg[2][17]  ( .D(block_next[17]), .E(n1281), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFX1 \block_reg[6][17]  ( .D(block_next[17]), .E(n1248), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFX1 \block_reg[2][16]  ( .D(block_next[16]), .E(n1281), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFX1 \block_reg[6][16]  ( .D(block_next[16]), .E(n1252), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFX1 \block_reg[2][15]  ( .D(block_next[15]), .E(n1281), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFX1 \block_reg[6][15]  ( .D(block_next[15]), .E(n1253), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFX1 \block_reg[2][14]  ( .D(block_next[14]), .E(n1281), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFX1 \block_reg[6][14]  ( .D(block_next[14]), .E(n1248), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFX1 \block_reg[2][13]  ( .D(block_next[13]), .E(n1281), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFX1 \block_reg[6][13]  ( .D(block_next[13]), .E(n1252), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFX1 \block_reg[2][12]  ( .D(block_next[12]), .E(n1280), .CK(clk), .Q(
        \block[2][12] ) );
  EDFFX1 \block_reg[6][12]  ( .D(block_next[12]), .E(n1246), .CK(clk), .Q(
        \block[6][12] ) );
  EDFFX1 \block_reg[2][11]  ( .D(block_next[11]), .E(n1280), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFX1 \block_reg[6][11]  ( .D(block_next[11]), .E(n1246), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFX1 \block_reg[2][10]  ( .D(block_next[10]), .E(n1280), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFX1 \block_reg[6][10]  ( .D(block_next[10]), .E(n1246), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFX1 \block_reg[2][9]  ( .D(block_next[9]), .E(n1280), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFX1 \block_reg[6][9]  ( .D(block_next[9]), .E(n1246), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFX1 \block_reg[2][8]  ( .D(block_next[8]), .E(n1280), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFX1 \block_reg[6][8]  ( .D(block_next[8]), .E(n1246), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFX1 \block_reg[2][7]  ( .D(block_next[7]), .E(n1280), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFX1 \block_reg[6][7]  ( .D(block_next[7]), .E(n1246), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFX1 \block_reg[2][6]  ( .D(block_next[6]), .E(n1280), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFX1 \block_reg[6][6]  ( .D(block_next[6]), .E(n1246), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFX1 \block_reg[2][5]  ( .D(block_next[5]), .E(n1280), .CK(clk), .Q(
        \block[2][5] ) );
  EDFFX1 \block_reg[6][5]  ( .D(block_next[5]), .E(n1246), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFX1 \block_reg[2][4]  ( .D(block_next[4]), .E(n1280), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFX1 \block_reg[6][4]  ( .D(block_next[4]), .E(n1246), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFX1 \block_reg[2][3]  ( .D(block_next[3]), .E(n1280), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFX1 \block_reg[6][3]  ( .D(block_next[3]), .E(n1246), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFX1 \block_reg[2][2]  ( .D(block_next[2]), .E(n1280), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFX1 \block_reg[6][2]  ( .D(block_next[2]), .E(n1246), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFX1 \block_reg[2][1]  ( .D(block_next[1]), .E(n1280), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFX1 \block_reg[6][1]  ( .D(block_next[1]), .E(n1246), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFX1 \block_reg[2][0]  ( .D(block_next[0]), .E(n1280), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFX1 \block_reg[6][0]  ( .D(block_next[0]), .E(n1250), .CK(clk), .Q(
        \block[6][0] ) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n612), .CK(clk), .RN(n1305), .Q(
        blockdirty[3]), .QN(n593) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n608), .CK(clk), .RN(n1305), .Q(
        blockdirty[7]), .QN(n589) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n614), .CK(clk), .RN(n1305), .Q(
        blockdirty[1]), .QN(n595) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n610), .CK(clk), .RN(n1305), .Q(
        blockdirty[5]), .QN(n591) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n615), .CK(clk), .RN(n1305), .Q(
        blockdirty[0]), .QN(n597) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n611), .CK(clk), .RN(n1305), .Q(
        blockdirty[4]), .QN(n592) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n613), .CK(clk), .RN(n1305), .Q(
        blockdirty[2]), .QN(n594) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n609), .CK(clk), .RN(n1305), .Q(
        blockdirty[6]), .QN(n590) );
  DFFX1 proc_read_r_reg ( .D(proc_read), .CK(clk), .QN(n1308) );
  DFFQX1 proc_write_r_reg ( .D(proc_write), .CK(clk), .Q(proc_write_r) );
  DFFQX1 \proc_addr_r_reg[25]  ( .D(proc_addr[25]), .CK(clk), .Q(dataTag[20])
         );
  DFFQX1 \proc_addr_r_reg[24]  ( .D(proc_addr[24]), .CK(clk), .Q(dataTag[19])
         );
  DFFQX1 \proc_addr_r_reg[20]  ( .D(proc_addr[20]), .CK(clk), .Q(dataTag[15])
         );
  DFFQX1 \proc_addr_r_reg[19]  ( .D(proc_addr[19]), .CK(clk), .Q(dataTag[14])
         );
  DFFQX1 \proc_addr_r_reg[18]  ( .D(proc_addr[18]), .CK(clk), .Q(dataTag[13])
         );
  DFFQX1 \proc_addr_r_reg[17]  ( .D(proc_addr[17]), .CK(clk), .Q(dataTag[12])
         );
  DFFQX1 \proc_addr_r_reg[16]  ( .D(proc_addr[16]), .CK(clk), .Q(dataTag[11])
         );
  DFFQX1 \proc_addr_r_reg[15]  ( .D(proc_addr[15]), .CK(clk), .Q(dataTag[10])
         );
  DFFQX1 \proc_addr_r_reg[14]  ( .D(proc_addr[14]), .CK(clk), .Q(dataTag[9])
         );
  DFFQX1 \proc_addr_r_reg[13]  ( .D(proc_addr[13]), .CK(clk), .Q(dataTag[8])
         );
  DFFQX1 \proc_addr_r_reg[8]  ( .D(proc_addr[8]), .CK(clk), .Q(dataTag[3]) );
  DFFQX1 \proc_addr_r_reg[6]  ( .D(proc_addr[6]), .CK(clk), .Q(dataTag[1]) );
  DFFQX1 \proc_addr_r_reg[5]  ( .D(proc_addr[5]), .CK(clk), .Q(dataTag[0]) );
  DFFQX1 \proc_addr_r_reg[29]  ( .D(proc_addr[29]), .CK(clk), .Q(dataTag[24])
         );
  DFFQX1 \proc_addr_r_reg[28]  ( .D(proc_addr[28]), .CK(clk), .Q(dataTag[23])
         );
  DFFQX1 \proc_addr_r_reg[27]  ( .D(proc_addr[27]), .CK(clk), .Q(dataTag[22])
         );
  DFFQX1 \proc_addr_r_reg[26]  ( .D(proc_addr[26]), .CK(clk), .Q(dataTag[21])
         );
  DFFQX1 \proc_addr_r_reg[23]  ( .D(proc_addr[23]), .CK(clk), .Q(dataTag[18])
         );
  DFFQX1 \proc_addr_r_reg[22]  ( .D(proc_addr[22]), .CK(clk), .Q(dataTag[17])
         );
  DFFQX1 \proc_addr_r_reg[21]  ( .D(proc_addr[21]), .CK(clk), .Q(dataTag[16])
         );
  DFFQX1 \proc_addr_r_reg[12]  ( .D(proc_addr[12]), .CK(clk), .Q(dataTag[7])
         );
  DFFQX1 \proc_addr_r_reg[11]  ( .D(proc_addr[11]), .CK(clk), .Q(dataTag[6])
         );
  DFFQX1 \proc_addr_r_reg[10]  ( .D(proc_addr[10]), .CK(clk), .Q(dataTag[5])
         );
  DFFQX1 \proc_addr_r_reg[9]  ( .D(proc_addr[9]), .CK(clk), .Q(dataTag[4]) );
  DFFQX1 \proc_addr_r_reg[7]  ( .D(proc_addr[7]), .CK(clk), .Q(dataTag[2]) );
  DFFQX1 \proc_addr_r_reg[0]  ( .D(proc_addr[0]), .CK(clk), .Q(wordIndex[0])
         );
  DFFQX1 \proc_addr_r_reg[1]  ( .D(proc_addr[1]), .CK(clk), .Q(wordIndex[1])
         );
  EDFFX1 \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n1271), .CK(clk), .Q(
        \blocktag[3][9] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n1237), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(N960), .CK(clk), .Q(
        \blocktag[3][8] ) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(N965), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(blocktag_next[7]), .E(N960), .CK(clk), .QN(
        n762) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(blocktag_next[7]), .E(N965), .CK(clk), .QN(
        n766) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(N960), .CK(clk), .QN(
        n754) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(N965), .CK(clk), .QN(
        n758) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(blocktag_next[5]), .E(n1271), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(blocktag_next[5]), .E(n1237), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(N960), .CK(clk), .QN(
        n778) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(N965), .CK(clk), .QN(
        n782) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n1271), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n1237), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n1271), .CK(clk), 
        .QN(n770) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n1237), .CK(clk), 
        .QN(n774) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n1271), .CK(clk), 
        .Q(\blocktag[3][24] ) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n1237), .CK(clk), 
        .Q(\blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(blocktag_next[23]), .E(n1271), .CK(clk), 
        .QN(n746) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(blocktag_next[23]), .E(n1237), .CK(clk), 
        .QN(n750) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n1279), .CK(clk), 
        .QN(n730) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n1245), .CK(clk), 
        .QN(n734) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n1279), .CK(clk), 
        .QN(n722) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n1245), .CK(clk), 
        .QN(n726) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][20] ) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n1279), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n1245), .CK(clk), .Q(
        \blocktag[7][1] ) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][19] ) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][19] ) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][18] ) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(blocktag_next[17]), .E(n1279), .CK(clk), 
        .QN(n714) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(blocktag_next[17]), .E(n1245), .CK(clk), 
        .QN(n718) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(n1279), .CK(clk), 
        .QN(n738) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(n1245), .CK(clk), 
        .QN(n742) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(blocktag_next[14]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][14] ) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(blocktag_next[14]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][14] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][13] ) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(blocktag_next[12]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][12] ) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(blocktag_next[12]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][12] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n1279), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n1245), .CK(clk), 
        .Q(\blocktag[7][11] ) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(blocktag_next[10]), .E(n1278), .CK(clk), 
        .Q(\blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(blocktag_next[10]), .E(n1244), .CK(clk), 
        .Q(\blocktag[7][10] ) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n1278), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n1244), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFX1 \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n1288), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n1262), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(N957), .CK(clk), .Q(
        \blocktag[1][8] ) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n1254), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(blocktag_next[7]), .E(N957), .CK(clk), .QN(
        n760) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(blocktag_next[7]), .E(n1262), .CK(clk), 
        .QN(n764) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(N957), .CK(clk), .QN(
        n752) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n1254), .CK(clk), 
        .QN(n756) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(blocktag_next[5]), .E(n1288), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(blocktag_next[5]), .E(n1258), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(N957), .CK(clk), .QN(
        n776) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n1258), .CK(clk), 
        .QN(n780) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n1288), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n1254), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n1288), .CK(clk), 
        .QN(n768) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n1262), .CK(clk), 
        .QN(n772) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n1288), .CK(clk), 
        .Q(\blocktag[1][24] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n1258), .CK(clk), 
        .Q(\blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(blocktag_next[23]), .E(n1288), .CK(clk), 
        .QN(n744) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(blocktag_next[23]), .E(n1258), .CK(clk), 
        .QN(n748) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n1296), .CK(clk), 
        .QN(n728) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n1257), .CK(clk), 
        .QN(n732) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n1296), .CK(clk), 
        .QN(n720) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n1255), .CK(clk), 
        .QN(n724) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][20] ) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n1260), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n1296), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n1259), .CK(clk), .Q(
        \blocktag[5][1] ) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][19] ) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n1261), .CK(clk), 
        .Q(\blocktag[5][19] ) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n1256), .CK(clk), 
        .Q(\blocktag[5][18] ) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(blocktag_next[17]), .E(n1296), .CK(clk), 
        .QN(n712) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(blocktag_next[17]), .E(n1256), .CK(clk), 
        .QN(n716) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n1296), .CK(clk), 
        .QN(n736) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(n1261), .CK(clk), 
        .QN(n740) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(n1255), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(blocktag_next[14]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][14] ) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(blocktag_next[14]), .E(n1257), .CK(clk), 
        .Q(\blocktag[5][14] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n1257), .CK(clk), 
        .Q(\blocktag[5][13] ) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(blocktag_next[12]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][12] ) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(blocktag_next[12]), .E(n1260), .CK(clk), 
        .Q(\blocktag[5][12] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n1296), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n1259), .CK(clk), 
        .Q(\blocktag[5][11] ) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(blocktag_next[10]), .E(n1295), .CK(clk), 
        .Q(\blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(blocktag_next[10]), .E(N962), .CK(clk), 
        .Q(\blocktag[5][10] ) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n1295), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(N962), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFX1 \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n1304), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n1265), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n1304), .CK(clk), .Q(
        \blocktag[0][8] ) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n1270), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(blocktag_next[7]), .E(n1304), .CK(clk), 
        .QN(n759) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(blocktag_next[7]), .E(n1269), .CK(clk), 
        .QN(n763) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n1301), .CK(clk), 
        .QN(n751) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n1270), .CK(clk), 
        .QN(n755) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(blocktag_next[5]), .E(n1304), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(blocktag_next[5]), .E(n1269), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n1302), .CK(clk), 
        .QN(n775) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n1265), .CK(clk), 
        .QN(n779) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n1304), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n1265), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n1298), .CK(clk), 
        .QN(n767) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n1269), .CK(clk), 
        .QN(n771) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n1304), .CK(clk), 
        .Q(\blocktag[0][24] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n1270), .CK(clk), 
        .Q(\blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(blocktag_next[23]), .E(n1300), .CK(clk), 
        .QN(n743) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(blocktag_next[23]), .E(n1265), .CK(clk), 
        .QN(n747) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n1300), .CK(clk), 
        .QN(n727) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n1264), .CK(clk), 
        .QN(n731) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n1297), .CK(clk), 
        .QN(n719) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n1270), .CK(clk), 
        .QN(n723) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][20] ) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n1266), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n1301), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n1264), .CK(clk), .Q(
        \blocktag[4][1] ) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][19] ) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n1264), .CK(clk), 
        .Q(\blocktag[4][19] ) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(n1268), .CK(clk), 
        .Q(\blocktag[4][18] ) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(blocktag_next[17]), .E(n1299), .CK(clk), 
        .QN(n711) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(blocktag_next[17]), .E(n1267), .CK(clk), 
        .QN(n715) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(n1301), .CK(clk), 
        .QN(n735) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(n1263), .CK(clk), 
        .QN(n739) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(n1298), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(n1263), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(blocktag_next[14]), .E(n1302), .CK(clk), 
        .Q(\blocktag[0][14] ) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(blocktag_next[14]), .E(n1266), .CK(clk), 
        .Q(\blocktag[4][14] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n1264), .CK(clk), 
        .Q(\blocktag[4][13] ) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(blocktag_next[12]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][12] ) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(blocktag_next[12]), .E(n696), .CK(clk), 
        .Q(\blocktag[4][12] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n1303), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n1268), .CK(clk), 
        .Q(\blocktag[4][11] ) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(blocktag_next[10]), .E(n1304), .CK(clk), 
        .Q(\blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(blocktag_next[10]), .E(n1270), .CK(clk), 
        .Q(\blocktag[4][10] ) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n1304), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n1270), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFX1 \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n1287), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n1248), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n1287), .CK(clk), .Q(
        \blocktag[2][8] ) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n1253), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(blocktag_next[7]), .E(n1287), .CK(clk), 
        .QN(n761) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(blocktag_next[7]), .E(n1252), .CK(clk), 
        .QN(n765) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n1285), .CK(clk), 
        .QN(n753) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n1253), .CK(clk), 
        .QN(n757) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(blocktag_next[5]), .E(n1287), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(blocktag_next[5]), .E(n1252), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n1281), .CK(clk), 
        .QN(n777) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n1248), .CK(clk), 
        .QN(n781) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n1287), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n1248), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n1283), .CK(clk), 
        .QN(n769) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n1252), .CK(clk), 
        .QN(n773) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n1287), .CK(clk), 
        .Q(\blocktag[2][24] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n1253), .CK(clk), 
        .Q(\blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(blocktag_next[23]), .E(n1286), .CK(clk), 
        .QN(n745) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(blocktag_next[23]), .E(n1248), .CK(clk), 
        .QN(n749) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n1283), .CK(clk), 
        .QN(n729) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n1247), .CK(clk), 
        .QN(n733) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n1281), .CK(clk), 
        .QN(n721) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n1253), .CK(clk), 
        .QN(n725) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n1286), .CK(clk), 
        .Q(\blocktag[2][20] ) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n1249), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n1283), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n1247), .CK(clk), .Q(
        \blocktag[6][1] ) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n1286), .CK(clk), 
        .Q(\blocktag[2][19] ) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n1247), .CK(clk), 
        .Q(\blocktag[6][19] ) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(n1280), .CK(clk), 
        .Q(\blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n1251), .CK(clk), 
        .Q(\blocktag[6][18] ) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(blocktag_next[17]), .E(n1285), .CK(clk), 
        .QN(n713) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(blocktag_next[17]), .E(n1250), .CK(clk), 
        .QN(n717) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(n1285), .CK(clk), 
        .QN(n737) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n1246), .CK(clk), 
        .QN(n741) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(n1283), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n1246), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(blocktag_next[14]), .E(n1281), .CK(clk), 
        .Q(\blocktag[2][14] ) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(blocktag_next[14]), .E(n1249), .CK(clk), 
        .Q(\blocktag[6][14] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n1286), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n1247), .CK(clk), 
        .Q(\blocktag[6][13] ) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(blocktag_next[12]), .E(n1286), .CK(clk), 
        .Q(\blocktag[2][12] ) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(blocktag_next[12]), .E(n695), .CK(clk), 
        .Q(\blocktag[6][12] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n1282), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n1251), .CK(clk), 
        .Q(\blocktag[6][11] ) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(blocktag_next[10]), .E(n1287), .CK(clk), 
        .Q(\blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(blocktag_next[10]), .E(n1253), .CK(clk), 
        .Q(\blocktag[6][10] ) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n1287), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n1253), .CK(clk), .Q(
        \blocktag[6][0] ) );
  DFFRX1 \blockvalid_reg[3]  ( .D(n620), .CK(clk), .RN(n1305), .Q(
        blockvalid[3]), .QN(n602) );
  DFFRX1 \blockvalid_reg[7]  ( .D(n616), .CK(clk), .RN(n1305), .Q(
        blockvalid[7]), .QN(n598) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n622), .CK(clk), .RN(n1305), .Q(
        blockvalid[1]), .QN(n604) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n618), .CK(clk), .RN(n1305), .Q(
        blockvalid[5]), .QN(n600) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n623), .CK(clk), .RN(n1305), .Q(
        blockvalid[0]), .QN(n605) );
  DFFRX1 \blockvalid_reg[4]  ( .D(n619), .CK(clk), .RN(n1305), .Q(
        blockvalid[4]), .QN(n601) );
  DFFRX1 \blockvalid_reg[2]  ( .D(n621), .CK(clk), .RN(n1305), .Q(
        blockvalid[2]), .QN(n603) );
  DFFRX1 \blockvalid_reg[6]  ( .D(n617), .CK(clk), .RN(n1305), .Q(
        blockvalid[6]), .QN(n599) );
  DFFRX1 \state_reg[1]  ( .D(state_next[1]), .CK(clk), .RN(n1305), .Q(state[1]), .QN(n1510) );
  DFFQX2 \proc_addr_r_reg[2]  ( .D(proc_addr[2]), .CK(clk), .Q(N85) );
  DFFQX1 mem_read_reg ( .D(mem_read_next), .CK(clk), .Q(mem_read) );
  EDFFX1 \mem_wdata_reg[127]  ( .D(blockdata[127]), .E(n1180), .CK(clk), .Q(
        mem_wdata[127]) );
  EDFFX1 \mem_wdata_reg[126]  ( .D(blockdata[126]), .E(n1179), .CK(clk), .Q(
        mem_wdata[126]) );
  EDFFX1 \mem_wdata_reg[125]  ( .D(blockdata[125]), .E(n1181), .CK(clk), .Q(
        mem_wdata[125]) );
  EDFFX1 \mem_wdata_reg[124]  ( .D(blockdata[124]), .E(n1180), .CK(clk), .Q(
        mem_wdata[124]) );
  EDFFX1 \mem_wdata_reg[123]  ( .D(blockdata[123]), .E(n1179), .CK(clk), .Q(
        mem_wdata[123]) );
  EDFFX1 \mem_wdata_reg[122]  ( .D(blockdata[122]), .E(n1181), .CK(clk), .Q(
        mem_wdata[122]) );
  EDFFX1 \mem_wdata_reg[121]  ( .D(blockdata[121]), .E(n1180), .CK(clk), .Q(
        mem_wdata[121]) );
  EDFFX1 \mem_wdata_reg[120]  ( .D(blockdata[120]), .E(n1179), .CK(clk), .Q(
        mem_wdata[120]) );
  EDFFX1 \mem_wdata_reg[119]  ( .D(blockdata[119]), .E(n1181), .CK(clk), .Q(
        mem_wdata[119]) );
  EDFFX1 \mem_wdata_reg[118]  ( .D(blockdata[118]), .E(n1180), .CK(clk), .Q(
        mem_wdata[118]) );
  EDFFX1 \mem_wdata_reg[117]  ( .D(blockdata[117]), .E(n1179), .CK(clk), .Q(
        mem_wdata[117]) );
  EDFFX1 \mem_wdata_reg[116]  ( .D(blockdata[116]), .E(n1181), .CK(clk), .Q(
        mem_wdata[116]) );
  EDFFX1 \mem_wdata_reg[115]  ( .D(blockdata[115]), .E(n1181), .CK(clk), .Q(
        mem_wdata[115]) );
  EDFFX1 \mem_wdata_reg[114]  ( .D(blockdata[114]), .E(n1181), .CK(clk), .Q(
        mem_wdata[114]) );
  EDFFX1 \mem_wdata_reg[113]  ( .D(blockdata[113]), .E(n1181), .CK(clk), .Q(
        mem_wdata[113]) );
  EDFFX1 \mem_wdata_reg[112]  ( .D(blockdata[112]), .E(n1181), .CK(clk), .Q(
        mem_wdata[112]) );
  EDFFX1 \mem_wdata_reg[111]  ( .D(blockdata[111]), .E(n1181), .CK(clk), .Q(
        mem_wdata[111]) );
  EDFFX1 \mem_wdata_reg[110]  ( .D(blockdata[110]), .E(n1181), .CK(clk), .Q(
        mem_wdata[110]) );
  EDFFX1 \mem_wdata_reg[109]  ( .D(blockdata[109]), .E(n1181), .CK(clk), .Q(
        mem_wdata[109]) );
  EDFFX1 \mem_wdata_reg[108]  ( .D(blockdata[108]), .E(n1181), .CK(clk), .Q(
        mem_wdata[108]) );
  EDFFX1 \mem_wdata_reg[107]  ( .D(blockdata[107]), .E(n1181), .CK(clk), .Q(
        mem_wdata[107]) );
  EDFFX1 \mem_wdata_reg[106]  ( .D(blockdata[106]), .E(n1181), .CK(clk), .Q(
        mem_wdata[106]) );
  EDFFX1 \mem_wdata_reg[105]  ( .D(blockdata[105]), .E(n1181), .CK(clk), .Q(
        mem_wdata[105]) );
  EDFFX1 \mem_wdata_reg[104]  ( .D(blockdata[104]), .E(n1181), .CK(clk), .Q(
        mem_wdata[104]) );
  EDFFX1 \mem_wdata_reg[103]  ( .D(blockdata[103]), .E(n1180), .CK(clk), .Q(
        mem_wdata[103]) );
  EDFFX1 \mem_wdata_reg[102]  ( .D(blockdata[102]), .E(n1180), .CK(clk), .Q(
        mem_wdata[102]) );
  EDFFX1 \mem_wdata_reg[101]  ( .D(blockdata[101]), .E(n1180), .CK(clk), .Q(
        mem_wdata[101]) );
  EDFFX1 \mem_wdata_reg[100]  ( .D(blockdata[100]), .E(n1180), .CK(clk), .Q(
        mem_wdata[100]) );
  EDFFX1 \mem_wdata_reg[99]  ( .D(blockdata[99]), .E(n1180), .CK(clk), .Q(
        mem_wdata[99]) );
  EDFFX1 \mem_wdata_reg[98]  ( .D(blockdata[98]), .E(n1180), .CK(clk), .Q(
        mem_wdata[98]) );
  EDFFX1 \mem_wdata_reg[97]  ( .D(blockdata[97]), .E(n1180), .CK(clk), .Q(
        mem_wdata[97]) );
  EDFFX1 \mem_wdata_reg[96]  ( .D(blockdata[96]), .E(n1180), .CK(clk), .Q(
        mem_wdata[96]) );
  EDFFX1 \mem_wdata_reg[95]  ( .D(blockdata[95]), .E(n1180), .CK(clk), .Q(
        mem_wdata[95]) );
  EDFFX1 \mem_wdata_reg[94]  ( .D(blockdata[94]), .E(n1180), .CK(clk), .Q(
        mem_wdata[94]) );
  EDFFX1 \mem_wdata_reg[93]  ( .D(blockdata[93]), .E(n1180), .CK(clk), .Q(
        mem_wdata[93]) );
  EDFFX1 \mem_wdata_reg[92]  ( .D(blockdata[92]), .E(n1180), .CK(clk), .Q(
        mem_wdata[92]) );
  EDFFX1 \mem_wdata_reg[91]  ( .D(blockdata[91]), .E(n1180), .CK(clk), .Q(
        mem_wdata[91]) );
  EDFFX1 \mem_wdata_reg[90]  ( .D(blockdata[90]), .E(n1179), .CK(clk), .Q(
        mem_wdata[90]) );
  EDFFX1 \mem_wdata_reg[89]  ( .D(blockdata[89]), .E(n1179), .CK(clk), .Q(
        mem_wdata[89]) );
  EDFFX1 \mem_wdata_reg[88]  ( .D(blockdata[88]), .E(n1179), .CK(clk), .Q(
        mem_wdata[88]) );
  EDFFX1 \mem_wdata_reg[87]  ( .D(blockdata[87]), .E(n1179), .CK(clk), .Q(
        mem_wdata[87]) );
  EDFFX1 \mem_wdata_reg[86]  ( .D(blockdata[86]), .E(n1179), .CK(clk), .Q(
        mem_wdata[86]) );
  EDFFX1 \mem_wdata_reg[85]  ( .D(blockdata[85]), .E(n1179), .CK(clk), .Q(
        mem_wdata[85]) );
  EDFFX1 \mem_wdata_reg[84]  ( .D(blockdata[84]), .E(n1179), .CK(clk), .Q(
        mem_wdata[84]) );
  EDFFX1 \mem_wdata_reg[83]  ( .D(blockdata[83]), .E(n1179), .CK(clk), .Q(
        mem_wdata[83]) );
  EDFFX1 \mem_wdata_reg[82]  ( .D(blockdata[82]), .E(n1179), .CK(clk), .Q(
        mem_wdata[82]) );
  EDFFX1 \mem_wdata_reg[81]  ( .D(blockdata[81]), .E(n1179), .CK(clk), .Q(
        mem_wdata[81]) );
  EDFFX1 \mem_wdata_reg[80]  ( .D(blockdata[80]), .E(n1179), .CK(clk), .Q(
        mem_wdata[80]) );
  EDFFX1 \mem_wdata_reg[79]  ( .D(blockdata[79]), .E(n1179), .CK(clk), .Q(
        mem_wdata[79]) );
  EDFFX1 \mem_wdata_reg[78]  ( .D(blockdata[78]), .E(n1179), .CK(clk), .Q(
        mem_wdata[78]) );
  EDFFX1 \mem_wdata_reg[77]  ( .D(blockdata[77]), .E(n1176), .CK(clk), .Q(
        mem_wdata[77]) );
  EDFFX1 \mem_wdata_reg[76]  ( .D(blockdata[76]), .E(n1176), .CK(clk), .Q(
        mem_wdata[76]) );
  EDFFX1 \mem_wdata_reg[75]  ( .D(blockdata[75]), .E(n1175), .CK(clk), .Q(
        mem_wdata[75]) );
  EDFFX1 \mem_wdata_reg[74]  ( .D(blockdata[74]), .E(n1177), .CK(clk), .Q(
        mem_wdata[74]) );
  EDFFX1 \mem_wdata_reg[73]  ( .D(blockdata[73]), .E(n1178), .CK(clk), .Q(
        mem_wdata[73]) );
  EDFFX1 \mem_wdata_reg[72]  ( .D(blockdata[72]), .E(n1177), .CK(clk), .Q(
        mem_wdata[72]) );
  EDFFX1 \mem_wdata_reg[71]  ( .D(blockdata[71]), .E(n1181), .CK(clk), .Q(
        mem_wdata[71]) );
  EDFFX1 \mem_wdata_reg[70]  ( .D(blockdata[70]), .E(n1180), .CK(clk), .Q(
        mem_wdata[70]) );
  EDFFX1 \mem_wdata_reg[69]  ( .D(blockdata[69]), .E(n1179), .CK(clk), .Q(
        mem_wdata[69]) );
  EDFFX1 \mem_wdata_reg[68]  ( .D(blockdata[68]), .E(n1181), .CK(clk), .Q(
        mem_wdata[68]) );
  EDFFX1 \mem_wdata_reg[67]  ( .D(blockdata[67]), .E(n1180), .CK(clk), .Q(
        mem_wdata[67]) );
  EDFFX1 \mem_wdata_reg[66]  ( .D(blockdata[66]), .E(n1179), .CK(clk), .Q(
        mem_wdata[66]) );
  EDFFX1 \mem_wdata_reg[65]  ( .D(blockdata[65]), .E(n1181), .CK(clk), .Q(
        mem_wdata[65]) );
  EDFFX1 \mem_wdata_reg[64]  ( .D(blockdata[64]), .E(n1177), .CK(clk), .Q(
        mem_wdata[64]) );
  EDFFX1 \mem_wdata_reg[63]  ( .D(blockdata[63]), .E(n1175), .CK(clk), .Q(
        mem_wdata[63]) );
  EDFFX1 \mem_wdata_reg[62]  ( .D(blockdata[62]), .E(n1178), .CK(clk), .Q(
        mem_wdata[62]) );
  EDFFX1 \mem_wdata_reg[61]  ( .D(blockdata[61]), .E(n1177), .CK(clk), .Q(
        mem_wdata[61]) );
  EDFFX1 \mem_wdata_reg[60]  ( .D(blockdata[60]), .E(n1175), .CK(clk), .Q(
        mem_wdata[60]) );
  EDFFX1 \mem_wdata_reg[59]  ( .D(blockdata[59]), .E(n1178), .CK(clk), .Q(
        mem_wdata[59]) );
  EDFFX1 \mem_wdata_reg[58]  ( .D(blockdata[58]), .E(n1177), .CK(clk), .Q(
        mem_wdata[58]) );
  EDFFX1 \mem_wdata_reg[57]  ( .D(blockdata[57]), .E(n1175), .CK(clk), .Q(
        mem_wdata[57]) );
  EDFFX1 \mem_wdata_reg[56]  ( .D(blockdata[56]), .E(n1178), .CK(clk), .Q(
        mem_wdata[56]) );
  EDFFX1 \mem_wdata_reg[55]  ( .D(blockdata[55]), .E(n1177), .CK(clk), .Q(
        mem_wdata[55]) );
  EDFFX1 \mem_wdata_reg[54]  ( .D(blockdata[54]), .E(n1176), .CK(clk), .Q(
        mem_wdata[54]) );
  EDFFX1 \mem_wdata_reg[53]  ( .D(blockdata[53]), .E(n1175), .CK(clk), .Q(
        mem_wdata[53]) );
  EDFFX1 \mem_wdata_reg[52]  ( .D(blockdata[52]), .E(n1178), .CK(clk), .Q(
        mem_wdata[52]) );
  EDFFX1 \mem_wdata_reg[51]  ( .D(blockdata[51]), .E(n1178), .CK(clk), .Q(
        mem_wdata[51]) );
  EDFFX1 \mem_wdata_reg[50]  ( .D(blockdata[50]), .E(n1178), .CK(clk), .Q(
        mem_wdata[50]) );
  EDFFX1 \mem_wdata_reg[49]  ( .D(blockdata[49]), .E(n1178), .CK(clk), .Q(
        mem_wdata[49]) );
  EDFFX1 \mem_wdata_reg[48]  ( .D(blockdata[48]), .E(n1178), .CK(clk), .Q(
        mem_wdata[48]) );
  EDFFX1 \mem_wdata_reg[47]  ( .D(blockdata[47]), .E(n1178), .CK(clk), .Q(
        mem_wdata[47]) );
  EDFFX1 \mem_wdata_reg[46]  ( .D(blockdata[46]), .E(n1178), .CK(clk), .Q(
        mem_wdata[46]) );
  EDFFX1 \mem_wdata_reg[45]  ( .D(blockdata[45]), .E(n1178), .CK(clk), .Q(
        mem_wdata[45]) );
  EDFFX1 \mem_wdata_reg[44]  ( .D(blockdata[44]), .E(n1178), .CK(clk), .Q(
        mem_wdata[44]) );
  EDFFX1 \mem_wdata_reg[43]  ( .D(blockdata[43]), .E(n1178), .CK(clk), .Q(
        mem_wdata[43]) );
  EDFFX1 \mem_wdata_reg[42]  ( .D(blockdata[42]), .E(n1178), .CK(clk), .Q(
        mem_wdata[42]) );
  EDFFX1 \mem_wdata_reg[41]  ( .D(blockdata[41]), .E(n1178), .CK(clk), .Q(
        mem_wdata[41]) );
  EDFFX1 \mem_wdata_reg[40]  ( .D(blockdata[40]), .E(n1178), .CK(clk), .Q(
        mem_wdata[40]) );
  EDFFX1 \mem_wdata_reg[39]  ( .D(blockdata[39]), .E(n1178), .CK(clk), .Q(
        mem_wdata[39]) );
  EDFFX1 \mem_wdata_reg[38]  ( .D(blockdata[38]), .E(n1177), .CK(clk), .Q(
        mem_wdata[38]) );
  EDFFX1 \mem_wdata_reg[37]  ( .D(blockdata[37]), .E(n1177), .CK(clk), .Q(
        mem_wdata[37]) );
  EDFFX1 \mem_wdata_reg[36]  ( .D(blockdata[36]), .E(n1177), .CK(clk), .Q(
        mem_wdata[36]) );
  EDFFX1 \mem_wdata_reg[35]  ( .D(blockdata[35]), .E(n1177), .CK(clk), .Q(
        mem_wdata[35]) );
  EDFFX1 \mem_wdata_reg[34]  ( .D(blockdata[34]), .E(n1177), .CK(clk), .Q(
        mem_wdata[34]) );
  EDFFX1 \mem_wdata_reg[33]  ( .D(blockdata[33]), .E(n1177), .CK(clk), .Q(
        mem_wdata[33]) );
  EDFFX1 \mem_wdata_reg[32]  ( .D(blockdata[32]), .E(n1177), .CK(clk), .Q(
        mem_wdata[32]) );
  EDFFX1 \mem_wdata_reg[31]  ( .D(blockdata[31]), .E(n1177), .CK(clk), .Q(
        mem_wdata[31]) );
  EDFFX1 \mem_wdata_reg[30]  ( .D(blockdata[30]), .E(n1177), .CK(clk), .Q(
        mem_wdata[30]) );
  EDFFX1 \mem_wdata_reg[29]  ( .D(blockdata[29]), .E(n1177), .CK(clk), .Q(
        mem_wdata[29]) );
  EDFFX1 \mem_wdata_reg[28]  ( .D(blockdata[28]), .E(n1177), .CK(clk), .Q(
        mem_wdata[28]) );
  EDFFX1 \mem_wdata_reg[27]  ( .D(blockdata[27]), .E(n1177), .CK(clk), .Q(
        mem_wdata[27]) );
  EDFFX1 \mem_wdata_reg[26]  ( .D(blockdata[26]), .E(n1177), .CK(clk), .Q(
        mem_wdata[26]) );
  EDFFX1 \mem_wdata_reg[25]  ( .D(blockdata[25]), .E(n1176), .CK(clk), .Q(
        mem_wdata[25]) );
  EDFFX1 \mem_wdata_reg[24]  ( .D(blockdata[24]), .E(n1176), .CK(clk), .Q(
        mem_wdata[24]) );
  EDFFX1 \mem_wdata_reg[23]  ( .D(blockdata[23]), .E(n1176), .CK(clk), .Q(
        mem_wdata[23]) );
  EDFFX1 \mem_wdata_reg[22]  ( .D(blockdata[22]), .E(n1176), .CK(clk), .Q(
        mem_wdata[22]) );
  EDFFX1 \mem_wdata_reg[21]  ( .D(blockdata[21]), .E(n1176), .CK(clk), .Q(
        mem_wdata[21]) );
  EDFFX1 \mem_wdata_reg[20]  ( .D(blockdata[20]), .E(n1176), .CK(clk), .Q(
        mem_wdata[20]) );
  EDFFX1 \mem_wdata_reg[19]  ( .D(blockdata[19]), .E(n1176), .CK(clk), .Q(
        mem_wdata[19]) );
  EDFFX1 \mem_wdata_reg[18]  ( .D(blockdata[18]), .E(n1176), .CK(clk), .Q(
        mem_wdata[18]) );
  EDFFX1 \mem_wdata_reg[17]  ( .D(blockdata[17]), .E(n1176), .CK(clk), .Q(
        mem_wdata[17]) );
  EDFFX1 \mem_wdata_reg[16]  ( .D(blockdata[16]), .E(n1176), .CK(clk), .Q(
        mem_wdata[16]) );
  EDFFX1 \mem_wdata_reg[15]  ( .D(blockdata[15]), .E(n1176), .CK(clk), .Q(
        mem_wdata[15]) );
  EDFFX1 \mem_wdata_reg[14]  ( .D(blockdata[14]), .E(n1176), .CK(clk), .Q(
        mem_wdata[14]) );
  EDFFX1 \mem_wdata_reg[13]  ( .D(blockdata[13]), .E(n1176), .CK(clk), .Q(
        mem_wdata[13]) );
  EDFFX1 \mem_wdata_reg[12]  ( .D(blockdata[12]), .E(n1175), .CK(clk), .Q(
        mem_wdata[12]) );
  EDFFX1 \mem_wdata_reg[11]  ( .D(blockdata[11]), .E(n1175), .CK(clk), .Q(
        mem_wdata[11]) );
  EDFFX1 \mem_wdata_reg[10]  ( .D(blockdata[10]), .E(n1175), .CK(clk), .Q(
        mem_wdata[10]) );
  EDFFX1 \mem_wdata_reg[9]  ( .D(blockdata[9]), .E(n1175), .CK(clk), .Q(
        mem_wdata[9]) );
  EDFFX1 \mem_wdata_reg[8]  ( .D(blockdata[8]), .E(n1175), .CK(clk), .Q(
        mem_wdata[8]) );
  EDFFX1 \mem_wdata_reg[7]  ( .D(blockdata[7]), .E(n1175), .CK(clk), .Q(
        mem_wdata[7]) );
  EDFFX1 \mem_wdata_reg[6]  ( .D(blockdata[6]), .E(n1175), .CK(clk), .Q(
        mem_wdata[6]) );
  EDFFX1 \mem_wdata_reg[5]  ( .D(blockdata[5]), .E(n1175), .CK(clk), .Q(
        mem_wdata[5]) );
  EDFFX1 \mem_wdata_reg[4]  ( .D(blockdata[4]), .E(n1175), .CK(clk), .Q(
        mem_wdata[4]) );
  EDFFX1 \mem_wdata_reg[3]  ( .D(blockdata[3]), .E(n1175), .CK(clk), .Q(
        mem_wdata[3]) );
  EDFFX1 \mem_wdata_reg[2]  ( .D(blockdata[2]), .E(n1175), .CK(clk), .Q(
        mem_wdata[2]) );
  EDFFX1 \mem_wdata_reg[1]  ( .D(blockdata[1]), .E(n1175), .CK(clk), .Q(
        mem_wdata[1]) );
  EDFFX1 \mem_wdata_reg[0]  ( .D(blockdata[0]), .E(n1175), .CK(clk), .Q(
        mem_wdata[0]) );
  DFFRX1 \state_reg[2]  ( .D(state_next[2]), .CK(clk), .RN(n1305), .Q(state[2]) );
  DFFRX1 \state_reg[0]  ( .D(state_next[0]), .CK(clk), .RN(n1305), .Q(state[0]) );
  DFFQX1 mem_write_reg ( .D(n1174), .CK(clk), .Q(mem_write) );
  DFFQX1 proc_stall_reg ( .D(proc_stall_next), .CK(clk), .Q(proc_stall) );
  EDFFX1 \mem_addr_reg[2]  ( .D(N87), .E(n1223), .CK(clk), .Q(mem_addr[2]) );
  EDFFX1 \mem_addr_reg[1]  ( .D(N86), .E(n1223), .CK(clk), .Q(mem_addr[1]) );
  EDFFX1 \mem_addr_reg[0]  ( .D(N85), .E(n1223), .CK(clk), .Q(mem_addr[0]) );
  DFFQX1 mem_ready_r_reg ( .D(mem_ready), .CK(clk), .Q(mem_ready_r) );
  DFFQXL \proc_rdata_reg[23]  ( .D(n674), .CK(clk), .Q(proc_rdata[23]) );
  DFFQXL \proc_rdata_reg[22]  ( .D(n673), .CK(clk), .Q(proc_rdata[22]) );
  DFFQXL \proc_rdata_reg[21]  ( .D(n672), .CK(clk), .Q(proc_rdata[21]) );
  DFFQXL \proc_rdata_reg[20]  ( .D(n671), .CK(clk), .Q(proc_rdata[20]) );
  DFFQXL \proc_rdata_reg[19]  ( .D(n670), .CK(clk), .Q(proc_rdata[19]) );
  DFFQXL \proc_rdata_reg[18]  ( .D(n669), .CK(clk), .Q(proc_rdata[18]) );
  DFFQXL \proc_rdata_reg[17]  ( .D(n668), .CK(clk), .Q(proc_rdata[17]) );
  DFFQXL \proc_rdata_reg[16]  ( .D(n667), .CK(clk), .Q(proc_rdata[16]) );
  DFFQXL \proc_rdata_reg[15]  ( .D(n666), .CK(clk), .Q(proc_rdata[15]) );
  DFFQXL \proc_rdata_reg[14]  ( .D(n665), .CK(clk), .Q(proc_rdata[14]) );
  DFFQXL \proc_rdata_reg[13]  ( .D(n664), .CK(clk), .Q(proc_rdata[13]) );
  DFFQXL \proc_rdata_reg[12]  ( .D(n663), .CK(clk), .Q(proc_rdata[12]) );
  DFFQXL \proc_rdata_reg[11]  ( .D(n662), .CK(clk), .Q(proc_rdata[11]) );
  DFFQXL \proc_rdata_reg[10]  ( .D(n661), .CK(clk), .Q(proc_rdata[10]) );
  DFFQXL \proc_rdata_reg[9]  ( .D(n660), .CK(clk), .Q(proc_rdata[9]) );
  DFFQXL \proc_rdata_reg[8]  ( .D(n659), .CK(clk), .Q(proc_rdata[8]) );
  DFFQXL \proc_rdata_reg[7]  ( .D(n658), .CK(clk), .Q(proc_rdata[7]) );
  DFFQXL \proc_rdata_reg[6]  ( .D(n657), .CK(clk), .Q(proc_rdata[6]) );
  DFFQXL \proc_rdata_reg[5]  ( .D(n656), .CK(clk), .Q(proc_rdata[5]) );
  DFFQXL \proc_rdata_reg[4]  ( .D(n655), .CK(clk), .Q(proc_rdata[4]) );
  DFFQXL \proc_rdata_reg[3]  ( .D(n654), .CK(clk), .Q(proc_rdata[3]) );
  DFFQXL \proc_rdata_reg[2]  ( .D(n653), .CK(clk), .Q(proc_rdata[2]) );
  DFFQXL \proc_rdata_reg[1]  ( .D(n652), .CK(clk), .Q(proc_rdata[1]) );
  DFFQXL \proc_rdata_reg[0]  ( .D(n651), .CK(clk), .Q(proc_rdata[0]) );
  DFFQXL \mem_addr_reg[25]  ( .D(n1310), .CK(clk), .Q(mem_addr[25]) );
  DFFQXL \mem_addr_reg[24]  ( .D(n1311), .CK(clk), .Q(mem_addr[24]) );
  DFFQXL \mem_addr_reg[23]  ( .D(n1312), .CK(clk), .Q(mem_addr[23]) );
  DFFQXL \mem_addr_reg[22]  ( .D(n1313), .CK(clk), .Q(mem_addr[22]) );
  DFFQXL \mem_addr_reg[21]  ( .D(n1314), .CK(clk), .Q(mem_addr[21]) );
  DFFQXL \mem_addr_reg[20]  ( .D(n1315), .CK(clk), .Q(mem_addr[20]) );
  DFFQXL \mem_addr_reg[19]  ( .D(n1316), .CK(clk), .Q(mem_addr[19]) );
  DFFQXL \mem_addr_reg[17]  ( .D(n1318), .CK(clk), .Q(mem_addr[17]) );
  DFFQXL \mem_addr_reg[16]  ( .D(n1319), .CK(clk), .Q(mem_addr[16]) );
  DFFQXL \mem_addr_reg[15]  ( .D(n1320), .CK(clk), .Q(mem_addr[15]) );
  DFFQXL \mem_addr_reg[14]  ( .D(n1321), .CK(clk), .Q(mem_addr[14]) );
  DFFQXL \mem_addr_reg[13]  ( .D(n1322), .CK(clk), .Q(mem_addr[13]) );
  DFFQXL \mem_addr_reg[12]  ( .D(n1323), .CK(clk), .Q(mem_addr[12]) );
  DFFQXL \mem_addr_reg[11]  ( .D(n1324), .CK(clk), .Q(mem_addr[11]) );
  DFFQXL \mem_addr_reg[10]  ( .D(n1325), .CK(clk), .Q(mem_addr[10]) );
  DFFQXL \mem_addr_reg[9]  ( .D(n1326), .CK(clk), .Q(mem_addr[9]) );
  DFFQXL \mem_addr_reg[8]  ( .D(n1327), .CK(clk), .Q(mem_addr[8]) );
  DFFQXL \mem_addr_reg[7]  ( .D(n1328), .CK(clk), .Q(mem_addr[7]) );
  DFFQXL \mem_addr_reg[6]  ( .D(n1329), .CK(clk), .Q(mem_addr[6]) );
  DFFQXL \mem_addr_reg[5]  ( .D(n1330), .CK(clk), .Q(mem_addr[5]) );
  DFFQXL \mem_addr_reg[4]  ( .D(n1331), .CK(clk), .Q(mem_addr[4]) );
  DFFQXL \mem_addr_reg[3]  ( .D(n1332), .CK(clk), .Q(mem_addr[3]) );
  DFFQXL \mem_addr_reg[27]  ( .D(n701), .CK(clk), .Q(mem_addr[27]) );
  DFFQXL \mem_addr_reg[18]  ( .D(n1317), .CK(clk), .Q(mem_addr[18]) );
  DFFQX1 \proc_addr_r_reg[4]  ( .D(proc_addr[4]), .CK(clk), .Q(N87) );
  DFFQXL \mem_addr_reg[26]  ( .D(n1309), .CK(clk), .Q(mem_addr[26]) );
  DFFX1 \proc_addr_r_reg[3]  ( .D(proc_addr[3]), .CK(clk), .Q(N86), .QN(n1472)
         );
  INVX1 U799 ( .A(n1169), .Y(n1306) );
  MX4X1 U800 ( .A(n759), .B(n760), .C(n761), .D(n762), .S0(n687), .S1(n1132), 
        .Y(n1079) );
  MXI2X2 U801 ( .A(n1057), .B(n1058), .S0(n1161), .Y(tag[18]) );
  MXI4X1 U802 ( .A(\blocktag[4][18] ), .B(\blocktag[5][18] ), .C(
        \blocktag[6][18] ), .D(\blocktag[7][18] ), .S0(n1106), .S1(n1134), .Y(
        n1058) );
  XOR2X4 U803 ( .A(tag[16]), .B(dataTag[16]), .Y(n482) );
  MXI2X2 U804 ( .A(n1047), .B(n1048), .S0(n1164), .Y(tag[23]) );
  CLKBUFX3 U805 ( .A(tag[0]), .Y(n683) );
  CLKBUFX3 U806 ( .A(tag[1]), .Y(n684) );
  CLKBUFX3 U807 ( .A(tag[3]), .Y(n685) );
  MXI2X2 U808 ( .A(n1049), .B(n1050), .S0(n1159), .Y(tag[22]) );
  MXI2X2 U809 ( .A(n1045), .B(n1046), .S0(n1164), .Y(tag[24]) );
  MXI2X2 U810 ( .A(n1059), .B(n1060), .S0(n1162), .Y(tag[17]) );
  CLKBUFX3 U811 ( .A(n1104), .Y(n686) );
  CLKBUFX3 U812 ( .A(n1104), .Y(n687) );
  CLKBUFX3 U813 ( .A(n1104), .Y(n688) );
  CLKBUFX2 U814 ( .A(n1102), .Y(n1104) );
  OAI222X1 U815 ( .A0(n1212), .A1(n1616), .B0(n1210), .B1(n1584), .C0(n1208), 
        .C1(n1520), .Y(n353) );
  OAI222X1 U816 ( .A0(n1211), .A1(n1628), .B0(n1210), .B1(n1596), .C0(n1207), 
        .C1(n1532), .Y(n209) );
  OAI222X4 U817 ( .A0(n1212), .A1(n1617), .B0(n1210), .B1(n1585), .C0(n1208), 
        .C1(n1521), .Y(n341) );
  OAI222X4 U818 ( .A0(n1211), .A1(n1629), .B0(n1210), .B1(n1597), .C0(n1207), 
        .C1(n1533), .Y(n197) );
  OAI222X4 U819 ( .A0(n1212), .A1(n1618), .B0(n1210), .B1(n1586), .C0(n1208), 
        .C1(n1522), .Y(n329) );
  OAI222X4 U820 ( .A0(n1211), .A1(n1630), .B0(n1210), .B1(n1598), .C0(n1207), 
        .C1(n1534), .Y(n185) );
  OAI222X4 U821 ( .A0(n1212), .A1(n1619), .B0(n1210), .B1(n1587), .C0(n1208), 
        .C1(n1523), .Y(n317) );
  OAI222X4 U822 ( .A0(n1211), .A1(n1631), .B0(n1210), .B1(n1599), .C0(n1207), 
        .C1(n1535), .Y(n173) );
  OAI222X4 U823 ( .A0(n1212), .A1(n1620), .B0(n1210), .B1(n1588), .C0(n1208), 
        .C1(n1524), .Y(n305) );
  OAI222X4 U824 ( .A0(n1211), .A1(n1632), .B0(n1210), .B1(n1600), .C0(n1207), 
        .C1(n1536), .Y(n161) );
  OAI222X4 U825 ( .A0(n1212), .A1(n1621), .B0(n1210), .B1(n1589), .C0(n1208), 
        .C1(n1525), .Y(n293) );
  OAI222X4 U826 ( .A0(n1211), .A1(n1633), .B0(n1210), .B1(n1601), .C0(n1207), 
        .C1(n1537), .Y(n149) );
  OAI222X4 U827 ( .A0(n1212), .A1(n1622), .B0(n1210), .B1(n1590), .C0(n1208), 
        .C1(n1526), .Y(n281) );
  OAI222X4 U828 ( .A0(n1211), .A1(n1634), .B0(n1210), .B1(n1602), .C0(n1207), 
        .C1(n1538), .Y(n137) );
  OAI222X4 U829 ( .A0(n1212), .A1(n1623), .B0(n1210), .B1(n1591), .C0(n1208), 
        .C1(n1527), .Y(n269) );
  OAI222X4 U830 ( .A0(n1211), .A1(n1635), .B0(n1210), .B1(n1603), .C0(n1207), 
        .C1(n1539), .Y(n125) );
  OAI222X4 U831 ( .A0(n1212), .A1(n1624), .B0(n1210), .B1(n1592), .C0(n1208), 
        .C1(n1528), .Y(n257) );
  OAI222X4 U832 ( .A0(n1211), .A1(n1636), .B0(n1210), .B1(n1604), .C0(n1207), 
        .C1(n1540), .Y(n113) );
  OAI222X4 U833 ( .A0(n1212), .A1(n1625), .B0(n1210), .B1(n1593), .C0(n1208), 
        .C1(n1529), .Y(n245) );
  OAI222X4 U834 ( .A0(n1211), .A1(n1637), .B0(n1210), .B1(n1605), .C0(n1207), 
        .C1(n1541), .Y(n101) );
  OAI222X4 U835 ( .A0(n1212), .A1(n1626), .B0(n1210), .B1(n1594), .C0(n1208), 
        .C1(n1530), .Y(n233) );
  OAI222X4 U836 ( .A0(n1211), .A1(n1638), .B0(n1210), .B1(n1606), .C0(n1207), 
        .C1(n1542), .Y(n89) );
  OAI222X4 U837 ( .A0(n1212), .A1(n1627), .B0(n1210), .B1(n1595), .C0(n1208), 
        .C1(n1531), .Y(n221) );
  OAI222X4 U838 ( .A0(n1211), .A1(n1639), .B0(n1210), .B1(n1607), .C0(n1207), 
        .C1(n1543), .Y(n68) );
  BUFX6 U839 ( .A(n76), .Y(n1210) );
  BUFX4 U840 ( .A(tag[21]), .Y(n689) );
  MXI2XL U841 ( .A(n1051), .B(n1052), .S0(n1162), .Y(tag[21]) );
  CLKBUFX3 U842 ( .A(tag[8]), .Y(n690) );
  CLKBUFX3 U843 ( .A(tag[5]), .Y(n691) );
  CLKBUFX3 U844 ( .A(tag[4]), .Y(n692) );
  MXI2X4 U845 ( .A(n1053), .B(n1054), .S0(n1159), .Y(tag[20]) );
  MXI4XL U846 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n1106), .S1(n1134), .Y(
        n1054) );
  MXI4XL U847 ( .A(\blocktag[0][20] ), .B(\blocktag[1][20] ), .C(
        \blocktag[2][20] ), .D(\blocktag[3][20] ), .S0(n1106), .S1(n1134), .Y(
        n1053) );
  CLKBUFX3 U848 ( .A(tag[12]), .Y(n693) );
  MXI2X2 U849 ( .A(n1089), .B(n1090), .S0(n1163), .Y(tag[2]) );
  CLKBUFX3 U850 ( .A(tag[19]), .Y(n694) );
  MXI2X2 U851 ( .A(n1075), .B(n1076), .S0(n1163), .Y(tag[9]) );
  MXI4XL U852 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(
        \blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n687), .S1(n1132), .Y(
        n1076) );
  MXI4XL U853 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(
        \blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n688), .S1(n1132), .Y(
        n1075) );
  MXI2X4 U854 ( .A(n1067), .B(n1068), .S0(n1160), .Y(tag[13]) );
  MXI4XL U855 ( .A(\blocktag[4][13] ), .B(\blocktag[5][13] ), .C(
        \blocktag[6][13] ), .D(\blocktag[7][13] ), .S0(n1105), .S1(n1133), .Y(
        n1068) );
  MXI4XL U856 ( .A(\blocktag[0][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[3][13] ), .S0(n1105), .S1(n1133), .Y(
        n1067) );
  MXI2X4 U857 ( .A(n1073), .B(n1074), .S0(n1163), .Y(tag[10]) );
  MXI4XL U858 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n687), .S1(n1132), .Y(
        n1074) );
  MXI4XL U859 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n687), .S1(n1132), .Y(
        n1073) );
  MXI2X4 U860 ( .A(n1081), .B(n1082), .S0(n1163), .Y(tag[6]) );
  MXI2X2 U861 ( .A(n1071), .B(n1072), .S0(n1160), .Y(tag[11]) );
  MXI4XL U862 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n686), .S1(n1133), .Y(
        n1072) );
  MXI4XL U863 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n688), .S1(n1133), .Y(
        n1071) );
  CLKAND2X12 U864 ( .A(n5), .B(n1223), .Y(n38) );
  CLKBUFX3 U865 ( .A(n1097), .Y(n1101) );
  CLKBUFX8 U866 ( .A(n453), .Y(n1169) );
  OR4X1 U867 ( .A(n496), .B(n497), .C(n498), .D(n499), .Y(n710) );
  CLKINVX1 U868 ( .A(n1124), .Y(n1096) );
  INVX3 U869 ( .A(N85), .Y(n1473) );
  NAND3X1 U870 ( .A(n6), .B(n1226), .C(n11), .Y(n37) );
  NOR3X2 U871 ( .A(state[0]), .B(state[2]), .C(n1510), .Y(n454) );
  NOR2X2 U872 ( .A(n703), .B(n20), .Y(n695) );
  NOR2X2 U873 ( .A(n703), .B(n24), .Y(n696) );
  NOR2X2 U874 ( .A(n703), .B(n28), .Y(n697) );
  NOR2X2 U875 ( .A(n703), .B(n32), .Y(n698) );
  NOR4BX1 U876 ( .AN(n11), .B(n1333), .C(n13), .D(n1334), .Y(n606) );
  AND2X2 U877 ( .A(n783), .B(n784), .Y(n699) );
  AND2X2 U878 ( .A(n708), .B(n709), .Y(n700) );
  NAND3X1 U879 ( .A(n704), .B(n705), .C(n706), .Y(n701) );
  OAI22XL U880 ( .A0(mem_ready_r), .A1(n9), .B0(n65), .B1(n1334), .Y(n650) );
  CLKINVX1 U881 ( .A(proc_reset), .Y(n702) );
  INVX3 U882 ( .A(n702), .Y(n703) );
  CLKINVX1 U883 ( .A(n1467), .Y(n1158) );
  CLKBUFX3 U884 ( .A(n1127), .Y(n1128) );
  OA22XL U885 ( .A0(n9), .A1(n1508), .B0(dirty), .B1(n65), .Y(n63) );
  CLKBUFX3 U886 ( .A(n1472), .Y(n1157) );
  NAND2X1 U887 ( .A(n1063), .B(n707), .Y(n708) );
  NAND2X1 U888 ( .A(n1064), .B(n1164), .Y(n709) );
  CLKBUFX3 U889 ( .A(n1130), .Y(n1132) );
  CLKBUFX3 U890 ( .A(n1127), .Y(n1129) );
  CLKBUFX3 U891 ( .A(n1158), .Y(n1163) );
  NAND2X1 U892 ( .A(n1065), .B(n707), .Y(n783) );
  NAND2X1 U893 ( .A(n1066), .B(n1160), .Y(n784) );
  XNOR2X1 U894 ( .A(dataTag[15]), .B(n700), .Y(n493) );
  AOI222XL U895 ( .A0(mem_addr[18]), .A1(n1220), .B0(n38), .B1(dataTag[15]), 
        .C0(n700), .C1(n1174), .Y(n54) );
  NAND2X1 U896 ( .A(mem_addr[27]), .B(n1220), .Y(n704) );
  NAND2XL U897 ( .A(n38), .B(dataTag[24]), .Y(n705) );
  NAND2XL U898 ( .A(tag[24]), .B(n1173), .Y(n706) );
  INVXL U899 ( .A(n1162), .Y(n707) );
  MXI4XL U900 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n1105), .S1(n1133), .Y(
        n1063) );
  MXI4XL U901 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n1105), .S1(n1133), .Y(
        n1064) );
  BUFX2 U902 ( .A(n1098), .Y(n1100) );
  CLKBUFX2 U903 ( .A(n1098), .Y(n1099) );
  CLKINVX1 U904 ( .A(n37), .Y(n1223) );
  CLKINVX1 U905 ( .A(n1157), .Y(n1125) );
  NAND2BXL U906 ( .AN(n5), .B(n6), .Y(state_next[1]) );
  CLKINVX1 U907 ( .A(n37), .Y(n1222) );
  INVXL U908 ( .A(n1124), .Y(n1095) );
  NAND2X1 U909 ( .A(n1307), .B(n460), .Y(n508) );
  NAND4BX2 U910 ( .AN(n710), .B(n471), .C(n472), .D(n473), .Y(n64) );
  NAND3X1 U911 ( .A(n1169), .B(n454), .C(n456), .Y(n76) );
  NAND3X1 U912 ( .A(n1169), .B(n454), .C(n461), .Y(n74) );
  NAND3X1 U913 ( .A(n1169), .B(n454), .C(n455), .Y(n72) );
  NAND3X1 U914 ( .A(n1169), .B(n10), .C(n461), .Y(n85) );
  NAND3X1 U915 ( .A(n1169), .B(n454), .C(n460), .Y(n78) );
  NAND3X1 U916 ( .A(n1169), .B(n10), .C(n456), .Y(n70) );
  NAND3X1 U917 ( .A(n1169), .B(n10), .C(n455), .Y(n80) );
  NAND3X1 U918 ( .A(n1169), .B(n10), .C(n460), .Y(n83) );
  NAND2X1 U919 ( .A(n1307), .B(n461), .Y(n505) );
  NAND2X1 U920 ( .A(n1307), .B(n456), .Y(n545) );
  NAND2X1 U921 ( .A(n1307), .B(n455), .Y(n514) );
  NAND2X1 U922 ( .A(n1226), .B(n546), .Y(n504) );
  NOR2XL U923 ( .A(n1467), .B(n1472), .Y(n550) );
  MX4XL U924 ( .A(n711), .B(n712), .C(n713), .D(n714), .S0(n1105), .S1(n1134), 
        .Y(n1059) );
  MX4XL U925 ( .A(n715), .B(n716), .C(n717), .D(n718), .S0(n1105), .S1(n1134), 
        .Y(n1060) );
  MX4XL U926 ( .A(n719), .B(n720), .C(n721), .D(n722), .S0(n1106), .S1(n1134), 
        .Y(n1051) );
  MX4XL U927 ( .A(n723), .B(n724), .C(n725), .D(n726), .S0(n1106), .S1(n1134), 
        .Y(n1052) );
  MX4XL U928 ( .A(n727), .B(n728), .C(n729), .D(n730), .S0(n1106), .S1(n1134), 
        .Y(n1049) );
  MX4XL U929 ( .A(n731), .B(n732), .C(n733), .D(n734), .S0(n1106), .S1(n1134), 
        .Y(n1050) );
  MX4XL U930 ( .A(n735), .B(n736), .C(n737), .D(n738), .S0(n1105), .S1(n1133), 
        .Y(n1061) );
  MX4XL U931 ( .A(n739), .B(n740), .C(n741), .D(n742), .S0(n1105), .S1(n1133), 
        .Y(n1062) );
  MX4XL U932 ( .A(n743), .B(n744), .C(n745), .D(n746), .S0(n1106), .S1(n1135), 
        .Y(n1047) );
  MX4XL U933 ( .A(n747), .B(n748), .C(n749), .D(n750), .S0(n1106), .S1(n1135), 
        .Y(n1048) );
  MXI4XL U934 ( .A(\blocktag[0][24] ), .B(\blocktag[1][24] ), .C(
        \blocktag[2][24] ), .D(\blocktag[3][24] ), .S0(n1106), .S1(n1135), .Y(
        n1045) );
  MXI4XL U935 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n1106), .S1(n1135), .Y(
        n1046) );
  MXI4XL U936 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n1105), .S1(n1134), .Y(
        n1057) );
  MX4XL U937 ( .A(n751), .B(n752), .C(n753), .D(n754), .S0(n687), .S1(n1132), 
        .Y(n1081) );
  MX4XL U938 ( .A(n755), .B(n756), .C(n757), .D(n758), .S0(n688), .S1(n1132), 
        .Y(n1082) );
  MX4XL U939 ( .A(n763), .B(n764), .C(n765), .D(n766), .S0(n686), .S1(n1132), 
        .Y(n1080) );
  MX4XL U940 ( .A(n767), .B(n768), .C(n769), .D(n770), .S0(n1103), .S1(n1131), 
        .Y(n1089) );
  MX4XL U941 ( .A(n771), .B(n772), .C(n773), .D(n774), .S0(n1103), .S1(n1131), 
        .Y(n1090) );
  MX4XL U942 ( .A(n775), .B(n776), .C(n777), .D(n778), .S0(n1103), .S1(n1131), 
        .Y(n1085) );
  MX4XL U943 ( .A(n779), .B(n780), .C(n781), .D(n782), .S0(n1103), .S1(n1131), 
        .Y(n1086) );
  MXI4XL U944 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(
        \blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n1103), .S1(n1132), .Y(
        n1083) );
  MXI4XL U945 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(
        \blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n688), .S1(n1132), .Y(
        n1084) );
  MXI4XL U946 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n1107), .S1(n1135), .Y(n1043) );
  MXI4XL U947 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n1107), .S1(n1135), .Y(n1044) );
  MXI4XL U948 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n1107), .S1(n1135), .Y(n1041) );
  MXI4XL U949 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n1107), .S1(n1135), .Y(n1042) );
  XNOR2X1 U950 ( .A(dataTag[14]), .B(n699), .Y(n492) );
  NOR2BX4 U951 ( .AN(n465), .B(proc_stall_next), .Y(n453) );
  INVX1 U952 ( .A(n50), .Y(n1321) );
  INVX1 U953 ( .A(n51), .Y(n1320) );
  INVX1 U954 ( .A(n52), .Y(n1319) );
  INVX1 U955 ( .A(n53), .Y(n1318) );
  AOI222XL U956 ( .A0(mem_addr[17]), .A1(n1220), .B0(n38), .B1(dataTag[14]), 
        .C0(n699), .C1(n1174), .Y(n53) );
  INVX1 U957 ( .A(n54), .Y(n1317) );
  INVX1 U958 ( .A(n55), .Y(n1316) );
  INVX1 U959 ( .A(n56), .Y(n1315) );
  INVX1 U960 ( .A(n57), .Y(n1314) );
  INVX1 U961 ( .A(n58), .Y(n1313) );
  INVX1 U962 ( .A(n59), .Y(n1312) );
  INVX1 U963 ( .A(n60), .Y(n1311) );
  INVX1 U964 ( .A(n61), .Y(n1310) );
  INVX1 U965 ( .A(n39), .Y(n1332) );
  INVX1 U966 ( .A(n40), .Y(n1331) );
  INVX1 U967 ( .A(n41), .Y(n1330) );
  INVX1 U968 ( .A(n42), .Y(n1329) );
  INVX1 U969 ( .A(n43), .Y(n1328) );
  INVX1 U970 ( .A(n44), .Y(n1327) );
  INVX1 U971 ( .A(n45), .Y(n1326) );
  INVX1 U972 ( .A(n46), .Y(n1325) );
  INVX1 U973 ( .A(n47), .Y(n1324) );
  INVX1 U974 ( .A(n48), .Y(n1323) );
  INVX1 U975 ( .A(n49), .Y(n1322) );
  INVX1 U976 ( .A(n62), .Y(n1309) );
  MXI4XL U977 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n1107), .S1(n1135), .Y(n1039) );
  MXI4XL U978 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n1107), .S1(n1135), .Y(n1040) );
  MXI4XL U979 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n1107), .S1(n1135), .Y(n1037) );
  MXI4XL U980 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n1107), .S1(n1135), .Y(n1038) );
  MXI4XL U981 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n1107), .S1(n1136), .Y(n1035) );
  MXI4XL U982 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n1107), .S1(n1136), .Y(n1036) );
  MXI4XL U983 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n1107), .S1(n1136), .Y(n1033) );
  MXI4XL U984 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n1107), .S1(n1136), .Y(n1034) );
  MXI4XL U985 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n1107), .S1(n1136), .Y(n1031) );
  NOR2X2 U986 ( .A(n1511), .B(state[0]), .Y(n10) );
  NAND2X1 U987 ( .A(n503), .B(state[0]), .Y(n9) );
  NAND3BXL U988 ( .AN(n7), .B(n1226), .C(n6), .Y(state_next[0]) );
  NOR2X1 U989 ( .A(wordIndex[0]), .B(wordIndex[1]), .Y(n461) );
  NOR2XL U990 ( .A(n1472), .B(N87), .Y(n555) );
  NOR2XL U991 ( .A(n1467), .B(N86), .Y(n554) );
  NOR2XL U992 ( .A(N87), .B(N86), .Y(n556) );
  MXI4XL U993 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n1105), .S1(n1133), .Y(
        n1065) );
  MXI4XL U994 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n1105), .S1(n1133), .Y(
        n1066) );
  INVX4 U995 ( .A(n1234), .Y(n1233) );
  INVX3 U996 ( .A(n1224), .Y(n1228) );
  INVX3 U997 ( .A(n1235), .Y(n1229) );
  INVX3 U998 ( .A(n1236), .Y(n1230) );
  INVX3 U999 ( .A(n1236), .Y(n1231) );
  INVX3 U1000 ( .A(n1225), .Y(n1227) );
  INVX3 U1001 ( .A(n1234), .Y(n1226) );
  INVX3 U1002 ( .A(n1235), .Y(n1232) );
  CLKBUFX3 U1003 ( .A(n1101), .Y(n1105) );
  CLKBUFX3 U1004 ( .A(n1100), .Y(n1107) );
  CLKBUFX3 U1005 ( .A(n1101), .Y(n1106) );
  CLKBUFX3 U1006 ( .A(n1102), .Y(n1103) );
  CLKBUFX3 U1007 ( .A(n1128), .Y(n1135) );
  CLKBUFX3 U1008 ( .A(n1129), .Y(n1134) );
  CLKBUFX3 U1009 ( .A(n1129), .Y(n1133) );
  CLKBUFX3 U1010 ( .A(n1099), .Y(n1108) );
  CLKBUFX3 U1011 ( .A(n1099), .Y(n1109) );
  CLKBUFX3 U1012 ( .A(n1099), .Y(n1110) );
  CLKBUFX3 U1013 ( .A(n1099), .Y(n1111) );
  CLKBUFX3 U1014 ( .A(n1120), .Y(n1112) );
  CLKBUFX3 U1015 ( .A(n1121), .Y(n1113) );
  CLKBUFX3 U1016 ( .A(n1099), .Y(n1114) );
  CLKBUFX3 U1017 ( .A(n1095), .Y(n1115) );
  CLKBUFX3 U1018 ( .A(n1110), .Y(n1116) );
  CLKBUFX3 U1019 ( .A(n1109), .Y(n1117) );
  CLKBUFX3 U1020 ( .A(n1121), .Y(n1118) );
  CLKBUFX3 U1021 ( .A(n1120), .Y(n1119) );
  CLKBUFX3 U1022 ( .A(n1095), .Y(n1120) );
  CLKBUFX3 U1023 ( .A(n1095), .Y(n1121) );
  CLKBUFX3 U1024 ( .A(n1099), .Y(n1122) );
  CLKBUFX3 U1025 ( .A(n1099), .Y(n1123) );
  CLKBUFX3 U1026 ( .A(n1128), .Y(n1136) );
  CLKBUFX3 U1027 ( .A(n1136), .Y(n1137) );
  CLKBUFX3 U1028 ( .A(n1136), .Y(n1138) );
  CLKBUFX3 U1029 ( .A(n1156), .Y(n1139) );
  CLKBUFX3 U1030 ( .A(n1155), .Y(n1140) );
  CLKBUFX3 U1031 ( .A(n1156), .Y(n1141) );
  CLKBUFX3 U1032 ( .A(n1156), .Y(n1142) );
  CLKBUFX3 U1033 ( .A(n1156), .Y(n1143) );
  CLKBUFX3 U1034 ( .A(n1156), .Y(n1144) );
  CLKBUFX3 U1035 ( .A(n1156), .Y(n1145) );
  CLKBUFX3 U1036 ( .A(n1156), .Y(n1146) );
  CLKBUFX3 U1037 ( .A(n1155), .Y(n1147) );
  CLKBUFX3 U1038 ( .A(n1155), .Y(n1148) );
  CLKBUFX3 U1039 ( .A(n1155), .Y(n1149) );
  CLKBUFX3 U1040 ( .A(n1156), .Y(n1150) );
  CLKBUFX3 U1041 ( .A(n1155), .Y(n1151) );
  CLKBUFX3 U1042 ( .A(n1155), .Y(n1152) );
  CLKBUFX3 U1043 ( .A(n1155), .Y(n1153) );
  CLKBUFX3 U1044 ( .A(n1155), .Y(n1154) );
  CLKBUFX3 U1045 ( .A(N86), .Y(n1155) );
  CLKBUFX3 U1046 ( .A(N86), .Y(n1156) );
  CLKBUFX3 U1047 ( .A(n1158), .Y(n1164) );
  CLKBUFX3 U1048 ( .A(n1224), .Y(n1235) );
  CLKBUFX3 U1049 ( .A(n1224), .Y(n1234) );
  CLKBUFX3 U1050 ( .A(n1176), .Y(n1177) );
  CLKBUFX3 U1051 ( .A(n1176), .Y(n1178) );
  CLKBUFX3 U1052 ( .A(n606), .Y(n1179) );
  CLKBUFX3 U1053 ( .A(n606), .Y(n1180) );
  CLKBUFX3 U1054 ( .A(n606), .Y(n1181) );
  CLKBUFX3 U1055 ( .A(n1130), .Y(n1131) );
  CLKBUFX3 U1056 ( .A(n1097), .Y(n1102) );
  CLKBUFX3 U1057 ( .A(n1166), .Y(n1165) );
  CLKBUFX3 U1058 ( .A(n1162), .Y(n1166) );
  CLKBUFX3 U1059 ( .A(n1165), .Y(n1167) );
  CLKBUFX3 U1060 ( .A(n1165), .Y(n1168) );
  CLKBUFX3 U1061 ( .A(n1234), .Y(n1236) );
  CLKBUFX3 U1062 ( .A(n1184), .Y(n1185) );
  CLKBUFX3 U1063 ( .A(n1188), .Y(n1189) );
  CLKBUFX3 U1064 ( .A(n1192), .Y(n1193) );
  INVX3 U1065 ( .A(n1222), .Y(n1220) );
  CLKBUFX3 U1066 ( .A(n1176), .Y(n1175) );
  CLKBUFX3 U1067 ( .A(n606), .Y(n1176) );
  CLKBUFX3 U1068 ( .A(n1225), .Y(n1224) );
  CLKBUFX3 U1069 ( .A(n1096), .Y(n1098) );
  CLKBUFX3 U1070 ( .A(n1125), .Y(n1127) );
  CLKBUFX3 U1071 ( .A(n1096), .Y(n1097) );
  CLKBUFX3 U1072 ( .A(n1126), .Y(n1130) );
  CLKBUFX3 U1073 ( .A(n1125), .Y(n1126) );
  CLKBUFX3 U1074 ( .A(n508), .Y(n1190) );
  CLKBUFX3 U1075 ( .A(n508), .Y(n1191) );
  CLKBUFX3 U1076 ( .A(n1237), .Y(n1238) );
  CLKBUFX3 U1077 ( .A(n1254), .Y(n1255) );
  CLKBUFX3 U1078 ( .A(n1271), .Y(n1272) );
  CLKBUFX3 U1079 ( .A(n1281), .Y(n1280) );
  CLKBUFX3 U1080 ( .A(n1288), .Y(n1289) );
  CLKBUFX3 U1081 ( .A(n1298), .Y(n1297) );
  CLKBUFX3 U1082 ( .A(n1237), .Y(n1239) );
  CLKBUFX3 U1083 ( .A(n1254), .Y(n1256) );
  CLKBUFX3 U1084 ( .A(n1271), .Y(n1273) );
  CLKBUFX3 U1085 ( .A(n697), .Y(n1281) );
  CLKBUFX3 U1086 ( .A(n1288), .Y(n1290) );
  CLKBUFX3 U1087 ( .A(n698), .Y(n1298) );
  CLKBUFX3 U1088 ( .A(n1237), .Y(n1240) );
  CLKBUFX3 U1089 ( .A(n1254), .Y(n1257) );
  CLKBUFX3 U1090 ( .A(n1271), .Y(n1274) );
  CLKBUFX3 U1091 ( .A(n1285), .Y(n1282) );
  CLKBUFX3 U1092 ( .A(n1288), .Y(n1291) );
  CLKBUFX3 U1093 ( .A(n1302), .Y(n1299) );
  CLKBUFX3 U1094 ( .A(n1237), .Y(n1241) );
  CLKBUFX3 U1095 ( .A(n1247), .Y(n1248) );
  CLKBUFX3 U1096 ( .A(n1254), .Y(n1258) );
  CLKBUFX3 U1097 ( .A(n1264), .Y(n1265) );
  CLKBUFX3 U1098 ( .A(n1271), .Y(n1275) );
  CLKBUFX3 U1099 ( .A(n697), .Y(n1283) );
  CLKBUFX3 U1100 ( .A(n1288), .Y(n1292) );
  CLKBUFX3 U1101 ( .A(n698), .Y(n1300) );
  CLKBUFX3 U1102 ( .A(n1237), .Y(n1242) );
  CLKBUFX3 U1103 ( .A(n1246), .Y(n1249) );
  CLKBUFX3 U1104 ( .A(n1254), .Y(n1259) );
  CLKBUFX3 U1105 ( .A(n1263), .Y(n1266) );
  CLKBUFX3 U1106 ( .A(n1271), .Y(n1276) );
  CLKBUFX3 U1107 ( .A(n697), .Y(n1284) );
  CLKBUFX3 U1108 ( .A(n1288), .Y(n1293) );
  CLKBUFX3 U1109 ( .A(n698), .Y(n1301) );
  CLKBUFX3 U1110 ( .A(n1246), .Y(n1250) );
  CLKBUFX3 U1111 ( .A(n1254), .Y(n1260) );
  CLKBUFX3 U1112 ( .A(n1263), .Y(n1267) );
  CLKBUFX3 U1113 ( .A(n697), .Y(n1285) );
  CLKBUFX3 U1114 ( .A(n698), .Y(n1302) );
  CLKBUFX3 U1115 ( .A(n1237), .Y(n1243) );
  CLKBUFX3 U1116 ( .A(n1246), .Y(n1251) );
  CLKBUFX3 U1117 ( .A(n1254), .Y(n1261) );
  CLKBUFX3 U1118 ( .A(n1263), .Y(n1268) );
  CLKBUFX3 U1119 ( .A(n1271), .Y(n1277) );
  CLKBUFX3 U1120 ( .A(n1288), .Y(n1294) );
  CLKBUFX3 U1121 ( .A(n1237), .Y(n1244) );
  CLKBUFX3 U1122 ( .A(n1247), .Y(n1252) );
  CLKBUFX3 U1123 ( .A(n1254), .Y(n1262) );
  CLKBUFX3 U1124 ( .A(n1264), .Y(n1269) );
  CLKBUFX3 U1125 ( .A(n1271), .Y(n1278) );
  CLKBUFX3 U1126 ( .A(n697), .Y(n1286) );
  CLKBUFX3 U1127 ( .A(n1288), .Y(n1295) );
  CLKBUFX3 U1128 ( .A(n698), .Y(n1303) );
  CLKBUFX3 U1129 ( .A(n1247), .Y(n1253) );
  CLKBUFX3 U1130 ( .A(n1264), .Y(n1270) );
  CLKBUFX3 U1131 ( .A(n697), .Y(n1287) );
  CLKBUFX3 U1132 ( .A(n698), .Y(n1304) );
  CLKBUFX3 U1133 ( .A(n1237), .Y(n1245) );
  CLKBUFX3 U1134 ( .A(n1271), .Y(n1279) );
  CLKBUFX3 U1135 ( .A(n1288), .Y(n1296) );
  CLKBUFX3 U1136 ( .A(n1158), .Y(n1162) );
  CLKBUFX3 U1137 ( .A(n1159), .Y(n1161) );
  NAND2X1 U1138 ( .A(n63), .B(n1509), .Y(n5) );
  CLKINVX1 U1139 ( .A(n64), .Y(n1333) );
  CLKBUFX3 U1140 ( .A(n80), .Y(n1204) );
  CLKBUFX3 U1141 ( .A(n80), .Y(n1205) );
  CLKBUFX3 U1142 ( .A(n70), .Y(n1217) );
  CLKBUFX3 U1143 ( .A(n83), .Y(n1201) );
  CLKBUFX3 U1144 ( .A(n70), .Y(n1218) );
  CLKBUFX3 U1145 ( .A(n83), .Y(n1202) );
  CLKBUFX3 U1146 ( .A(n72), .Y(n1214) );
  CLKBUFX3 U1147 ( .A(n72), .Y(n1215) );
  CLKBUFX3 U1148 ( .A(n85), .Y(n1198) );
  CLKBUFX3 U1149 ( .A(n85), .Y(n1199) );
  CLKBUFX3 U1150 ( .A(n78), .Y(n1207) );
  CLKBUFX3 U1151 ( .A(n78), .Y(n1208) );
  CLKBUFX3 U1152 ( .A(n74), .Y(n1211) );
  CLKBUFX3 U1153 ( .A(n74), .Y(n1212) );
  CLKBUFX3 U1154 ( .A(n504), .Y(n1196) );
  CLKBUFX3 U1155 ( .A(n80), .Y(n1206) );
  CLKBUFX3 U1156 ( .A(n72), .Y(n1216) );
  CLKBUFX3 U1157 ( .A(n70), .Y(n1219) );
  CLKBUFX3 U1158 ( .A(n83), .Y(n1203) );
  CLKBUFX3 U1159 ( .A(n85), .Y(n1200) );
  CLKBUFX3 U1160 ( .A(n1306), .Y(n1171) );
  CLKBUFX3 U1161 ( .A(n1306), .Y(n1170) );
  CLKBUFX3 U1162 ( .A(n504), .Y(n1197) );
  CLKBUFX3 U1163 ( .A(n78), .Y(n1209) );
  CLKBUFX3 U1164 ( .A(n74), .Y(n1213) );
  CLKBUFX3 U1165 ( .A(n1306), .Y(n1172) );
  CLKBUFX3 U1166 ( .A(n33), .Y(n1225) );
  CLKBUFX3 U1167 ( .A(n514), .Y(n1186) );
  CLKBUFX3 U1168 ( .A(n514), .Y(n1187) );
  CLKBUFX3 U1169 ( .A(n545), .Y(n1183) );
  CLKBUFX3 U1170 ( .A(n545), .Y(n1182) );
  CLKBUFX3 U1171 ( .A(n505), .Y(n1195) );
  CLKBUFX3 U1172 ( .A(n505), .Y(n1194) );
  CLKBUFX3 U1173 ( .A(n1158), .Y(n1159) );
  CLKBUFX3 U1174 ( .A(n1158), .Y(n1160) );
  CLKBUFX3 U1175 ( .A(n1247), .Y(n1246) );
  CLKBUFX3 U1176 ( .A(n1264), .Y(n1263) );
  CLKINVX1 U1177 ( .A(n20), .Y(n1463) );
  CLKINVX1 U1178 ( .A(n24), .Y(n1465) );
  CLKINVX1 U1179 ( .A(n28), .Y(n1468) );
  CLKINVX1 U1180 ( .A(n32), .Y(n1470) );
  OAI222X4 U1181 ( .A0(n1639), .A1(n1226), .B0(n1335), .B1(n1197), .C0(n505), 
        .C1(n1507), .Y(block_next[0]) );
  OAI222X4 U1182 ( .A0(n1638), .A1(n1228), .B0(n1336), .B1(n1196), .C0(n1195), 
        .C1(n1506), .Y(block_next[1]) );
  OAI222X4 U1183 ( .A0(n1637), .A1(n1228), .B0(n1337), .B1(n1197), .C0(n1194), 
        .C1(n1505), .Y(block_next[2]) );
  OAI222X4 U1184 ( .A0(n1636), .A1(n1229), .B0(n1338), .B1(n1197), .C0(n1194), 
        .C1(n1504), .Y(block_next[3]) );
  OAI222X4 U1185 ( .A0(n1635), .A1(n1229), .B0(n1339), .B1(n1197), .C0(n1194), 
        .C1(n1503), .Y(block_next[4]) );
  OAI222X4 U1186 ( .A0(n1634), .A1(n1230), .B0(n1340), .B1(n1197), .C0(n1194), 
        .C1(n1502), .Y(block_next[5]) );
  OAI222X4 U1187 ( .A0(n1633), .A1(n1231), .B0(n1341), .B1(n1196), .C0(n1194), 
        .C1(n1501), .Y(block_next[6]) );
  OAI222X4 U1188 ( .A0(n1632), .A1(n1231), .B0(n1342), .B1(n1197), .C0(n1194), 
        .C1(n1500), .Y(block_next[7]) );
  OAI222X4 U1189 ( .A0(n1631), .A1(n1232), .B0(n1343), .B1(n504), .C0(n1194), 
        .C1(n1499), .Y(block_next[8]) );
  OAI222X4 U1190 ( .A0(n1630), .A1(n1232), .B0(n1344), .B1(n504), .C0(n1194), 
        .C1(n1498), .Y(block_next[9]) );
  OAI222X4 U1191 ( .A0(n1629), .A1(n1226), .B0(n1345), .B1(n1197), .C0(n505), 
        .C1(n1497), .Y(block_next[10]) );
  OAI222X4 U1192 ( .A0(n1628), .A1(n1227), .B0(n1346), .B1(n1197), .C0(n1195), 
        .C1(n1496), .Y(block_next[11]) );
  OAI222X4 U1193 ( .A0(n1627), .A1(n1227), .B0(n1347), .B1(n1197), .C0(n1194), 
        .C1(n1495), .Y(block_next[12]) );
  OAI222X4 U1194 ( .A0(n1626), .A1(n1227), .B0(n1348), .B1(n1197), .C0(n1195), 
        .C1(n1494), .Y(block_next[13]) );
  OAI222X4 U1195 ( .A0(n1625), .A1(n1227), .B0(n1349), .B1(n1197), .C0(n1194), 
        .C1(n1493), .Y(block_next[14]) );
  OAI222X4 U1196 ( .A0(n1624), .A1(n1228), .B0(n1350), .B1(n1197), .C0(n505), 
        .C1(n1492), .Y(block_next[15]) );
  OAI222X4 U1197 ( .A0(n1623), .A1(n1228), .B0(n1351), .B1(n1197), .C0(n505), 
        .C1(n1491), .Y(block_next[16]) );
  OAI222X4 U1198 ( .A0(n1622), .A1(n1230), .B0(n1352), .B1(n1196), .C0(n1195), 
        .C1(n1490), .Y(block_next[17]) );
  OAI222X4 U1199 ( .A0(n1621), .A1(n1228), .B0(n1353), .B1(n1196), .C0(n1195), 
        .C1(n1489), .Y(block_next[18]) );
  OAI222X4 U1200 ( .A0(n1620), .A1(n1228), .B0(n1354), .B1(n1196), .C0(n1195), 
        .C1(n1488), .Y(block_next[19]) );
  OAI222X4 U1201 ( .A0(n1619), .A1(n1228), .B0(n1355), .B1(n1196), .C0(n1195), 
        .C1(n1487), .Y(block_next[20]) );
  OAI222X4 U1202 ( .A0(n1618), .A1(n1228), .B0(n1356), .B1(n1196), .C0(n1195), 
        .C1(n1486), .Y(block_next[21]) );
  OAI222X4 U1203 ( .A0(n1617), .A1(n1228), .B0(n1357), .B1(n1196), .C0(n1195), 
        .C1(n1485), .Y(block_next[22]) );
  OAI222X4 U1204 ( .A0(n1616), .A1(n1228), .B0(n1358), .B1(n1196), .C0(n1195), 
        .C1(n1484), .Y(block_next[23]) );
  OAI222X4 U1205 ( .A0(n1615), .A1(n1228), .B0(n1359), .B1(n1196), .C0(n1195), 
        .C1(n1483), .Y(block_next[24]) );
  OAI222X4 U1206 ( .A0(n1614), .A1(n1228), .B0(n1360), .B1(n1196), .C0(n1195), 
        .C1(n1482), .Y(block_next[25]) );
  OAI222X4 U1207 ( .A0(n1613), .A1(n1228), .B0(n1361), .B1(n1196), .C0(n1195), 
        .C1(n1481), .Y(block_next[26]) );
  OAI222X4 U1208 ( .A0(n1612), .A1(n1228), .B0(n1362), .B1(n1196), .C0(n1195), 
        .C1(n1480), .Y(block_next[27]) );
  OAI222X4 U1209 ( .A0(n1611), .A1(n1228), .B0(n1363), .B1(n1196), .C0(n1194), 
        .C1(n1479), .Y(block_next[28]) );
  OAI222X4 U1210 ( .A0(n1610), .A1(n1228), .B0(n1364), .B1(n1197), .C0(n1194), 
        .C1(n1478), .Y(block_next[29]) );
  OAI222X4 U1211 ( .A0(n1609), .A1(n1228), .B0(n1365), .B1(n504), .C0(n1194), 
        .C1(n1477), .Y(block_next[30]) );
  OAI222X4 U1212 ( .A0(n1608), .A1(n1228), .B0(n1366), .B1(n504), .C0(n1194), 
        .C1(n1476), .Y(block_next[31]) );
  OAI222X4 U1213 ( .A0(n1607), .A1(n1228), .B0(n1367), .B1(n1185), .C0(n1507), 
        .C1(n1183), .Y(block_next[32]) );
  OAI222X4 U1214 ( .A0(n1606), .A1(n1229), .B0(n1368), .B1(n1185), .C0(n1506), 
        .C1(n1182), .Y(block_next[33]) );
  OAI222X4 U1215 ( .A0(n1605), .A1(n1229), .B0(n1369), .B1(n1184), .C0(n1505), 
        .C1(n1183), .Y(block_next[34]) );
  OAI222X4 U1216 ( .A0(n1604), .A1(n1229), .B0(n1370), .B1(n1184), .C0(n1504), 
        .C1(n1182), .Y(block_next[35]) );
  OAI222X4 U1217 ( .A0(n1603), .A1(n1229), .B0(n1371), .B1(n1184), .C0(n1503), 
        .C1(n545), .Y(block_next[36]) );
  OAI222X4 U1218 ( .A0(n1602), .A1(n1229), .B0(n1372), .B1(n1184), .C0(n1502), 
        .C1(n545), .Y(block_next[37]) );
  OAI222X4 U1219 ( .A0(n1601), .A1(n1229), .B0(n1373), .B1(n1184), .C0(n1501), 
        .C1(n545), .Y(block_next[38]) );
  OAI222X4 U1220 ( .A0(n1600), .A1(n1229), .B0(n1374), .B1(n1184), .C0(n1500), 
        .C1(n545), .Y(block_next[39]) );
  OAI222X4 U1221 ( .A0(n1599), .A1(n1229), .B0(n1375), .B1(n1185), .C0(n1499), 
        .C1(n1183), .Y(block_next[40]) );
  OAI222X4 U1222 ( .A0(n1598), .A1(n1229), .B0(n1376), .B1(n1185), .C0(n1498), 
        .C1(n1183), .Y(block_next[41]) );
  OAI222X4 U1223 ( .A0(n1597), .A1(n1229), .B0(n1377), .B1(n1185), .C0(n1497), 
        .C1(n1183), .Y(block_next[42]) );
  OAI222X4 U1224 ( .A0(n1596), .A1(n1229), .B0(n1378), .B1(n1185), .C0(n1496), 
        .C1(n1183), .Y(block_next[43]) );
  OAI222X4 U1225 ( .A0(n1595), .A1(n1229), .B0(n1379), .B1(n1185), .C0(n1495), 
        .C1(n1183), .Y(block_next[44]) );
  OAI222X4 U1226 ( .A0(n1594), .A1(n1229), .B0(n1380), .B1(n1185), .C0(n1494), 
        .C1(n1183), .Y(block_next[45]) );
  OAI222X4 U1227 ( .A0(n1593), .A1(n1229), .B0(n1381), .B1(n1185), .C0(n1493), 
        .C1(n1183), .Y(block_next[46]) );
  OAI222X4 U1228 ( .A0(n1592), .A1(n1229), .B0(n1382), .B1(n1185), .C0(n1492), 
        .C1(n1183), .Y(block_next[47]) );
  OAI222X4 U1229 ( .A0(n1591), .A1(n1229), .B0(n1383), .B1(n1185), .C0(n1491), 
        .C1(n1183), .Y(block_next[48]) );
  OAI222X4 U1230 ( .A0(n1590), .A1(n1229), .B0(n1384), .B1(n1185), .C0(n1490), 
        .C1(n1183), .Y(block_next[49]) );
  OAI222X4 U1231 ( .A0(n1589), .A1(n1230), .B0(n1385), .B1(n1185), .C0(n1489), 
        .C1(n1183), .Y(block_next[50]) );
  OAI222X4 U1232 ( .A0(n1588), .A1(n1230), .B0(n1386), .B1(n1185), .C0(n1488), 
        .C1(n1183), .Y(block_next[51]) );
  OAI222X4 U1233 ( .A0(n1587), .A1(n1230), .B0(n1387), .B1(n1184), .C0(n1487), 
        .C1(n1182), .Y(block_next[52]) );
  OAI222X4 U1234 ( .A0(n1586), .A1(n1230), .B0(n1388), .B1(n1184), .C0(n1486), 
        .C1(n1182), .Y(block_next[53]) );
  OAI222X4 U1235 ( .A0(n1585), .A1(n1230), .B0(n1389), .B1(n1184), .C0(n1485), 
        .C1(n1182), .Y(block_next[54]) );
  OAI222X4 U1236 ( .A0(n1584), .A1(n1230), .B0(n1390), .B1(n1184), .C0(n1484), 
        .C1(n1182), .Y(block_next[55]) );
  OAI222X4 U1237 ( .A0(n1583), .A1(n1230), .B0(n1391), .B1(n1184), .C0(n1483), 
        .C1(n1182), .Y(block_next[56]) );
  OAI222X4 U1238 ( .A0(n1582), .A1(n1230), .B0(n1392), .B1(n1184), .C0(n1482), 
        .C1(n1182), .Y(block_next[57]) );
  OAI222X4 U1239 ( .A0(n1581), .A1(n1230), .B0(n1393), .B1(n1184), .C0(n1481), 
        .C1(n1182), .Y(block_next[58]) );
  OAI222X4 U1240 ( .A0(n1580), .A1(n1230), .B0(n1394), .B1(n1184), .C0(n1480), 
        .C1(n1182), .Y(block_next[59]) );
  OAI222X4 U1241 ( .A0(n1579), .A1(n1230), .B0(n1395), .B1(n1184), .C0(n1479), 
        .C1(n1182), .Y(block_next[60]) );
  OAI222X4 U1242 ( .A0(n1578), .A1(n1230), .B0(n1396), .B1(n1184), .C0(n1478), 
        .C1(n1182), .Y(block_next[61]) );
  OAI222X4 U1243 ( .A0(n1577), .A1(n1230), .B0(n1397), .B1(n1184), .C0(n1477), 
        .C1(n1182), .Y(block_next[62]) );
  OAI222X4 U1244 ( .A0(n1576), .A1(n1230), .B0(n1398), .B1(n544), .C0(n1476), 
        .C1(n1182), .Y(block_next[63]) );
  OAI222X4 U1245 ( .A0(n1575), .A1(n1230), .B0(n1399), .B1(n1188), .C0(n1507), 
        .C1(n1186), .Y(block_next[64]) );
  OAI222X4 U1246 ( .A0(n1574), .A1(n1230), .B0(n1400), .B1(n1189), .C0(n1506), 
        .C1(n1186), .Y(block_next[65]) );
  OAI222X4 U1247 ( .A0(n1573), .A1(n1230), .B0(n1401), .B1(n1188), .C0(n1505), 
        .C1(n1186), .Y(block_next[66]) );
  OAI222X4 U1248 ( .A0(n1572), .A1(n1231), .B0(n1402), .B1(n1188), .C0(n1504), 
        .C1(n1186), .Y(block_next[67]) );
  OAI222X4 U1249 ( .A0(n1571), .A1(n1231), .B0(n1403), .B1(n1188), .C0(n1186), 
        .C1(n1503), .Y(block_next[68]) );
  OAI222X4 U1250 ( .A0(n1570), .A1(n1231), .B0(n1404), .B1(n1188), .C0(n1186), 
        .C1(n1502), .Y(block_next[69]) );
  OAI222X4 U1251 ( .A0(n1569), .A1(n1231), .B0(n1405), .B1(n1188), .C0(n1186), 
        .C1(n1501), .Y(block_next[70]) );
  OAI222X4 U1252 ( .A0(n1568), .A1(n1231), .B0(n1406), .B1(n1188), .C0(n1186), 
        .C1(n1500), .Y(block_next[71]) );
  OAI222X4 U1253 ( .A0(n1567), .A1(n1231), .B0(n1407), .B1(n1188), .C0(n1187), 
        .C1(n1499), .Y(block_next[72]) );
  OAI222X4 U1254 ( .A0(n1566), .A1(n1231), .B0(n1408), .B1(n1188), .C0(n1498), 
        .C1(n1186), .Y(block_next[73]) );
  OAI222X4 U1255 ( .A0(n1565), .A1(n1231), .B0(n1409), .B1(n1188), .C0(n1186), 
        .C1(n1497), .Y(block_next[74]) );
  OAI222X4 U1256 ( .A0(n1564), .A1(n1231), .B0(n1410), .B1(n1188), .C0(n1186), 
        .C1(n1496), .Y(block_next[75]) );
  OAI222X4 U1257 ( .A0(n1563), .A1(n1231), .B0(n1411), .B1(n1188), .C0(n1186), 
        .C1(n1495), .Y(block_next[76]) );
  OAI222X4 U1258 ( .A0(n1562), .A1(n1231), .B0(n1412), .B1(n1188), .C0(n1187), 
        .C1(n1494), .Y(block_next[77]) );
  OAI222X4 U1259 ( .A0(n1561), .A1(n1231), .B0(n1413), .B1(n1188), .C0(n1187), 
        .C1(n1493), .Y(block_next[78]) );
  OAI222X4 U1260 ( .A0(n1560), .A1(n1231), .B0(n1414), .B1(n1188), .C0(n1187), 
        .C1(n1492), .Y(block_next[79]) );
  OAI222X4 U1261 ( .A0(n1559), .A1(n1231), .B0(n1415), .B1(n1188), .C0(n1187), 
        .C1(n1491), .Y(block_next[80]) );
  OAI222X4 U1262 ( .A0(n1558), .A1(n1231), .B0(n1416), .B1(n513), .C0(n1187), 
        .C1(n1490), .Y(block_next[81]) );
  OAI222X4 U1263 ( .A0(n1557), .A1(n1231), .B0(n1417), .B1(n1188), .C0(n1187), 
        .C1(n1489), .Y(block_next[82]) );
  OAI222X4 U1264 ( .A0(n1556), .A1(n1231), .B0(n1418), .B1(n1188), .C0(n1187), 
        .C1(n1488), .Y(block_next[83]) );
  OAI222X4 U1265 ( .A0(n1555), .A1(n1232), .B0(n1419), .B1(n1189), .C0(n1187), 
        .C1(n1487), .Y(block_next[84]) );
  OAI222X4 U1266 ( .A0(n1554), .A1(n1232), .B0(n1420), .B1(n1189), .C0(n1187), 
        .C1(n1486), .Y(block_next[85]) );
  OAI222X4 U1267 ( .A0(n1553), .A1(n1232), .B0(n1421), .B1(n1189), .C0(n1187), 
        .C1(n1485), .Y(block_next[86]) );
  OAI222X4 U1268 ( .A0(n1552), .A1(n1232), .B0(n1422), .B1(n1189), .C0(n1187), 
        .C1(n1484), .Y(block_next[87]) );
  OAI222X4 U1269 ( .A0(n1551), .A1(n1232), .B0(n1423), .B1(n1189), .C0(n1187), 
        .C1(n1483), .Y(block_next[88]) );
  OAI222X4 U1270 ( .A0(n1550), .A1(n1232), .B0(n1424), .B1(n1189), .C0(n1186), 
        .C1(n1482), .Y(block_next[89]) );
  OAI222X4 U1271 ( .A0(n1549), .A1(n1232), .B0(n1425), .B1(n1189), .C0(n1187), 
        .C1(n1481), .Y(block_next[90]) );
  OAI222X4 U1272 ( .A0(n1548), .A1(n1232), .B0(n1426), .B1(n1189), .C0(n1186), 
        .C1(n1480), .Y(block_next[91]) );
  OAI222X4 U1273 ( .A0(n1547), .A1(n1232), .B0(n1427), .B1(n1189), .C0(n1187), 
        .C1(n1479), .Y(block_next[92]) );
  OAI222X4 U1274 ( .A0(n1546), .A1(n1232), .B0(n1428), .B1(n1189), .C0(n514), 
        .C1(n1478), .Y(block_next[93]) );
  OAI222X4 U1275 ( .A0(n1545), .A1(n1232), .B0(n1429), .B1(n1189), .C0(n514), 
        .C1(n1477), .Y(block_next[94]) );
  OAI222X4 U1276 ( .A0(n1544), .A1(n1232), .B0(n1430), .B1(n1189), .C0(n1186), 
        .C1(n1476), .Y(block_next[95]) );
  OAI222X4 U1277 ( .A0(n1543), .A1(n1232), .B0(n1431), .B1(n1193), .C0(n1191), 
        .C1(n1507), .Y(block_next[96]) );
  OAI222X4 U1278 ( .A0(n1542), .A1(n1232), .B0(n1432), .B1(n1193), .C0(n508), 
        .C1(n1506), .Y(block_next[97]) );
  OAI222X4 U1279 ( .A0(n1541), .A1(n1232), .B0(n1433), .B1(n1193), .C0(n508), 
        .C1(n1505), .Y(block_next[98]) );
  OAI222X4 U1280 ( .A0(n1540), .A1(n1232), .B0(n1434), .B1(n1193), .C0(n1190), 
        .C1(n1504), .Y(block_next[99]) );
  OAI222X4 U1281 ( .A0(n1539), .A1(n1226), .B0(n1435), .B1(n1192), .C0(n1191), 
        .C1(n1503), .Y(block_next[100]) );
  OAI222X4 U1282 ( .A0(n1538), .A1(n1226), .B0(n1436), .B1(n1193), .C0(n1190), 
        .C1(n1502), .Y(block_next[101]) );
  OAI222X4 U1283 ( .A0(n1537), .A1(n1226), .B0(n1437), .B1(n1192), .C0(n1190), 
        .C1(n1501), .Y(block_next[102]) );
  OAI222X4 U1284 ( .A0(n1536), .A1(n1226), .B0(n1438), .B1(n1192), .C0(n1190), 
        .C1(n1500), .Y(block_next[103]) );
  OAI222X4 U1285 ( .A0(n1535), .A1(n1226), .B0(n1439), .B1(n1192), .C0(n1190), 
        .C1(n1499), .Y(block_next[104]) );
  OAI222X4 U1286 ( .A0(n1534), .A1(n1226), .B0(n1440), .B1(n1192), .C0(n1498), 
        .C1(n1190), .Y(block_next[105]) );
  OAI222X4 U1287 ( .A0(n1533), .A1(n1226), .B0(n1441), .B1(n1192), .C0(n1190), 
        .C1(n1497), .Y(block_next[106]) );
  OAI222X4 U1288 ( .A0(n1532), .A1(n1226), .B0(n1442), .B1(n1192), .C0(n1190), 
        .C1(n1496), .Y(block_next[107]) );
  OAI222X4 U1289 ( .A0(n1531), .A1(n1226), .B0(n1443), .B1(n1192), .C0(n1190), 
        .C1(n1495), .Y(block_next[108]) );
  OAI222X4 U1290 ( .A0(n1530), .A1(n1226), .B0(n1444), .B1(n1192), .C0(n1190), 
        .C1(n1494), .Y(block_next[109]) );
  OAI222X4 U1291 ( .A0(n1529), .A1(n1226), .B0(n1445), .B1(n1192), .C0(n1190), 
        .C1(n1493), .Y(block_next[110]) );
  OAI222X4 U1292 ( .A0(n1528), .A1(n1226), .B0(n1446), .B1(n507), .C0(n1190), 
        .C1(n1492), .Y(block_next[111]) );
  OAI222X4 U1293 ( .A0(n1527), .A1(n1227), .B0(n1447), .B1(n1192), .C0(n1190), 
        .C1(n1491), .Y(block_next[112]) );
  OAI222X4 U1294 ( .A0(n1526), .A1(n1226), .B0(n1448), .B1(n1192), .C0(n1191), 
        .C1(n1490), .Y(block_next[113]) );
  OAI222X4 U1295 ( .A0(n1525), .A1(n1227), .B0(n1449), .B1(n1192), .C0(n1191), 
        .C1(n1489), .Y(block_next[114]) );
  OAI222X4 U1296 ( .A0(n1524), .A1(n1227), .B0(n1450), .B1(n1192), .C0(n1191), 
        .C1(n1488), .Y(block_next[115]) );
  OAI222X4 U1297 ( .A0(n1523), .A1(n1227), .B0(n1451), .B1(n1192), .C0(n1191), 
        .C1(n1487), .Y(block_next[116]) );
  OAI222X4 U1298 ( .A0(n1522), .A1(n1227), .B0(n1452), .B1(n1192), .C0(n1191), 
        .C1(n1486), .Y(block_next[117]) );
  OAI222X4 U1299 ( .A0(n1521), .A1(n1227), .B0(n1453), .B1(n1192), .C0(n1191), 
        .C1(n1485), .Y(block_next[118]) );
  OAI222X4 U1300 ( .A0(n1520), .A1(n1227), .B0(n1454), .B1(n1192), .C0(n1191), 
        .C1(n1484), .Y(block_next[119]) );
  OAI222X4 U1301 ( .A0(n1519), .A1(n1227), .B0(n1455), .B1(n1193), .C0(n1191), 
        .C1(n1483), .Y(block_next[120]) );
  OAI222X4 U1302 ( .A0(n1518), .A1(n1227), .B0(n1456), .B1(n1193), .C0(n1191), 
        .C1(n1482), .Y(block_next[121]) );
  OAI222X4 U1303 ( .A0(n1517), .A1(n1227), .B0(n1457), .B1(n1193), .C0(n1191), 
        .C1(n1481), .Y(block_next[122]) );
  OAI222X4 U1304 ( .A0(n1516), .A1(n1227), .B0(n1458), .B1(n1193), .C0(n1191), 
        .C1(n1480), .Y(block_next[123]) );
  OAI222X4 U1305 ( .A0(n1515), .A1(n1227), .B0(n1459), .B1(n1193), .C0(n1191), 
        .C1(n1479), .Y(block_next[124]) );
  OAI222X4 U1306 ( .A0(n1514), .A1(n1227), .B0(n1460), .B1(n1193), .C0(n1190), 
        .C1(n1478), .Y(block_next[125]) );
  OAI222X4 U1307 ( .A0(n1513), .A1(n1227), .B0(n1461), .B1(n1193), .C0(n1191), 
        .C1(n1477), .Y(block_next[126]) );
  OAI222X4 U1308 ( .A0(n1512), .A1(n1227), .B0(n1462), .B1(n1193), .C0(n1190), 
        .C1(n1476), .Y(block_next[127]) );
  OAI222XL U1309 ( .A0(n1213), .A1(n1615), .B0(n1210), .B1(n1583), .C0(n1209), 
        .C1(n1519), .Y(n365) );
  OAI222XL U1310 ( .A0(n1213), .A1(n1614), .B0(n1210), .B1(n1582), .C0(n1209), 
        .C1(n1518), .Y(n377) );
  OAI222XL U1311 ( .A0(n1213), .A1(n1613), .B0(n1210), .B1(n1581), .C0(n1209), 
        .C1(n1517), .Y(n389) );
  OAI222XL U1312 ( .A0(n1213), .A1(n1612), .B0(n1210), .B1(n1580), .C0(n1209), 
        .C1(n1516), .Y(n401) );
  OAI222XL U1313 ( .A0(n1213), .A1(n1611), .B0(n1210), .B1(n1579), .C0(n1209), 
        .C1(n1515), .Y(n413) );
  OAI222XL U1314 ( .A0(n1213), .A1(n1610), .B0(n1210), .B1(n1578), .C0(n1209), 
        .C1(n1514), .Y(n425) );
  OAI222XL U1315 ( .A0(n1213), .A1(n1609), .B0(n1210), .B1(n1577), .C0(n1209), 
        .C1(n1513), .Y(n437) );
  OAI222XL U1316 ( .A0(n1213), .A1(n1608), .B0(n1210), .B1(n1576), .C0(n1209), 
        .C1(n1512), .Y(n449) );
  OR4X1 U1317 ( .A(n34), .B(n460), .C(n456), .D(n455), .Y(n546) );
  CLKINVX1 U1318 ( .A(n454), .Y(n1509) );
  NAND2X1 U1319 ( .A(n10), .B(n1333), .Y(n6) );
  NAND2X1 U1320 ( .A(n10), .B(n64), .Y(n65) );
  NOR2X1 U1321 ( .A(n1509), .B(n1508), .Y(n33) );
  NOR4X1 U1322 ( .A(n481), .B(n482), .C(n483), .D(n484), .Y(n472) );
  NOR4X1 U1323 ( .A(n474), .B(n475), .C(n476), .D(n477), .Y(n473) );
  CLKINVX1 U1324 ( .A(n34), .Y(n1307) );
  NAND2BX1 U1325 ( .AN(n461), .B(n1307), .Y(n543) );
  NAND4X1 U1326 ( .A(n466), .B(n11), .C(n65), .D(n9), .Y(proc_stall_next) );
  NAND2X1 U1327 ( .A(n454), .B(n1508), .Y(n466) );
  CLKINVX1 U1328 ( .A(dirty), .Y(n1334) );
  CLKBUFX3 U1329 ( .A(n650), .Y(n1174) );
  CLKBUFX3 U1330 ( .A(n650), .Y(n1173) );
  CLKBUFX3 U1331 ( .A(n1473), .Y(n1124) );
  NAND2X1 U1332 ( .A(n1509), .B(n9), .Y(n13) );
  CLKBUFX3 U1333 ( .A(n544), .Y(n1184) );
  OAI31XL U1334 ( .A0(n543), .A1(n455), .A2(n460), .B0(n1233), .Y(n544) );
  CLKBUFX3 U1335 ( .A(n513), .Y(n1188) );
  OAI31XL U1336 ( .A0(n543), .A1(n456), .A2(n460), .B0(n1232), .Y(n513) );
  CLKBUFX3 U1337 ( .A(n507), .Y(n1192) );
  OAI31XL U1338 ( .A0(n543), .A1(n455), .A2(n456), .B0(n1233), .Y(n507) );
  NOR2X2 U1339 ( .A(valid), .B(n1236), .Y(n35) );
  OA21X2 U1340 ( .A0(n1236), .A1(n1334), .B0(n34), .Y(n17) );
  NOR2X2 U1341 ( .A(n1474), .B(n1475), .Y(n460) );
  NAND2X1 U1342 ( .A(n550), .B(n1473), .Y(n20) );
  NAND2X1 U1343 ( .A(n554), .B(n1473), .Y(n24) );
  NAND2X1 U1344 ( .A(n555), .B(n1473), .Y(n28) );
  NAND2X1 U1345 ( .A(n556), .B(n1473), .Y(n32) );
  CLKINVX1 U1346 ( .A(blockdata[64]), .Y(n1399) );
  CLKINVX1 U1347 ( .A(blockdata[65]), .Y(n1400) );
  CLKINVX1 U1348 ( .A(blockdata[66]), .Y(n1401) );
  CLKINVX1 U1349 ( .A(blockdata[67]), .Y(n1402) );
  CLKINVX1 U1350 ( .A(blockdata[68]), .Y(n1403) );
  CLKINVX1 U1351 ( .A(blockdata[69]), .Y(n1404) );
  CLKINVX1 U1352 ( .A(blockdata[70]), .Y(n1405) );
  CLKINVX1 U1353 ( .A(blockdata[71]), .Y(n1406) );
  CLKINVX1 U1354 ( .A(blockdata[72]), .Y(n1407) );
  CLKINVX1 U1355 ( .A(blockdata[73]), .Y(n1408) );
  CLKINVX1 U1356 ( .A(blockdata[74]), .Y(n1409) );
  CLKINVX1 U1357 ( .A(blockdata[75]), .Y(n1410) );
  CLKINVX1 U1358 ( .A(blockdata[76]), .Y(n1411) );
  CLKINVX1 U1359 ( .A(blockdata[77]), .Y(n1412) );
  CLKINVX1 U1360 ( .A(blockdata[78]), .Y(n1413) );
  CLKINVX1 U1361 ( .A(blockdata[79]), .Y(n1414) );
  CLKINVX1 U1362 ( .A(blockdata[80]), .Y(n1415) );
  CLKINVX1 U1363 ( .A(blockdata[81]), .Y(n1416) );
  CLKINVX1 U1364 ( .A(blockdata[82]), .Y(n1417) );
  CLKINVX1 U1365 ( .A(blockdata[83]), .Y(n1418) );
  CLKINVX1 U1366 ( .A(blockdata[84]), .Y(n1419) );
  CLKINVX1 U1367 ( .A(blockdata[85]), .Y(n1420) );
  CLKINVX1 U1368 ( .A(blockdata[86]), .Y(n1421) );
  CLKINVX1 U1369 ( .A(blockdata[87]), .Y(n1422) );
  CLKINVX1 U1370 ( .A(blockdata[88]), .Y(n1423) );
  CLKINVX1 U1371 ( .A(blockdata[89]), .Y(n1424) );
  CLKINVX1 U1372 ( .A(blockdata[90]), .Y(n1425) );
  CLKINVX1 U1373 ( .A(blockdata[91]), .Y(n1426) );
  CLKINVX1 U1374 ( .A(blockdata[92]), .Y(n1427) );
  CLKINVX1 U1375 ( .A(blockdata[93]), .Y(n1428) );
  CLKINVX1 U1376 ( .A(blockdata[94]), .Y(n1429) );
  CLKINVX1 U1377 ( .A(blockdata[95]), .Y(n1430) );
  CLKINVX1 U1378 ( .A(blockdata[32]), .Y(n1367) );
  CLKINVX1 U1379 ( .A(blockdata[96]), .Y(n1431) );
  CLKINVX1 U1380 ( .A(blockdata[33]), .Y(n1368) );
  CLKINVX1 U1381 ( .A(blockdata[97]), .Y(n1432) );
  CLKINVX1 U1382 ( .A(blockdata[34]), .Y(n1369) );
  CLKINVX1 U1383 ( .A(blockdata[98]), .Y(n1433) );
  CLKINVX1 U1384 ( .A(blockdata[35]), .Y(n1370) );
  CLKINVX1 U1385 ( .A(blockdata[99]), .Y(n1434) );
  CLKINVX1 U1386 ( .A(blockdata[36]), .Y(n1371) );
  CLKINVX1 U1387 ( .A(blockdata[100]), .Y(n1435) );
  CLKINVX1 U1388 ( .A(blockdata[37]), .Y(n1372) );
  CLKINVX1 U1389 ( .A(blockdata[101]), .Y(n1436) );
  CLKINVX1 U1390 ( .A(blockdata[38]), .Y(n1373) );
  CLKINVX1 U1391 ( .A(blockdata[102]), .Y(n1437) );
  CLKINVX1 U1392 ( .A(blockdata[39]), .Y(n1374) );
  CLKINVX1 U1393 ( .A(blockdata[103]), .Y(n1438) );
  CLKINVX1 U1394 ( .A(blockdata[40]), .Y(n1375) );
  CLKINVX1 U1395 ( .A(blockdata[104]), .Y(n1439) );
  CLKINVX1 U1396 ( .A(blockdata[41]), .Y(n1376) );
  CLKINVX1 U1397 ( .A(blockdata[105]), .Y(n1440) );
  CLKINVX1 U1398 ( .A(blockdata[42]), .Y(n1377) );
  CLKINVX1 U1399 ( .A(blockdata[106]), .Y(n1441) );
  CLKINVX1 U1400 ( .A(blockdata[43]), .Y(n1378) );
  CLKINVX1 U1401 ( .A(blockdata[107]), .Y(n1442) );
  CLKINVX1 U1402 ( .A(blockdata[44]), .Y(n1379) );
  CLKINVX1 U1403 ( .A(blockdata[108]), .Y(n1443) );
  CLKINVX1 U1404 ( .A(blockdata[45]), .Y(n1380) );
  CLKINVX1 U1405 ( .A(blockdata[109]), .Y(n1444) );
  CLKINVX1 U1406 ( .A(blockdata[46]), .Y(n1381) );
  CLKINVX1 U1407 ( .A(blockdata[110]), .Y(n1445) );
  CLKINVX1 U1408 ( .A(blockdata[47]), .Y(n1382) );
  CLKINVX1 U1409 ( .A(blockdata[111]), .Y(n1446) );
  CLKINVX1 U1410 ( .A(blockdata[48]), .Y(n1383) );
  CLKINVX1 U1411 ( .A(blockdata[112]), .Y(n1447) );
  CLKINVX1 U1412 ( .A(blockdata[49]), .Y(n1384) );
  CLKINVX1 U1413 ( .A(blockdata[113]), .Y(n1448) );
  CLKINVX1 U1414 ( .A(blockdata[50]), .Y(n1385) );
  CLKINVX1 U1415 ( .A(blockdata[114]), .Y(n1449) );
  CLKINVX1 U1416 ( .A(blockdata[51]), .Y(n1386) );
  CLKINVX1 U1417 ( .A(blockdata[115]), .Y(n1450) );
  CLKINVX1 U1418 ( .A(blockdata[52]), .Y(n1387) );
  CLKINVX1 U1419 ( .A(blockdata[116]), .Y(n1451) );
  CLKINVX1 U1420 ( .A(blockdata[53]), .Y(n1388) );
  CLKINVX1 U1421 ( .A(blockdata[117]), .Y(n1452) );
  CLKINVX1 U1422 ( .A(blockdata[54]), .Y(n1389) );
  CLKINVX1 U1423 ( .A(blockdata[118]), .Y(n1453) );
  CLKINVX1 U1424 ( .A(blockdata[55]), .Y(n1390) );
  CLKINVX1 U1425 ( .A(blockdata[119]), .Y(n1454) );
  CLKINVX1 U1426 ( .A(blockdata[56]), .Y(n1391) );
  CLKINVX1 U1427 ( .A(blockdata[120]), .Y(n1455) );
  CLKINVX1 U1428 ( .A(blockdata[57]), .Y(n1392) );
  CLKINVX1 U1429 ( .A(blockdata[121]), .Y(n1456) );
  CLKINVX1 U1430 ( .A(blockdata[58]), .Y(n1393) );
  CLKINVX1 U1431 ( .A(blockdata[122]), .Y(n1457) );
  CLKINVX1 U1432 ( .A(blockdata[59]), .Y(n1394) );
  CLKINVX1 U1433 ( .A(blockdata[123]), .Y(n1458) );
  CLKINVX1 U1434 ( .A(blockdata[60]), .Y(n1395) );
  CLKINVX1 U1435 ( .A(blockdata[124]), .Y(n1459) );
  CLKINVX1 U1436 ( .A(blockdata[61]), .Y(n1396) );
  CLKINVX1 U1437 ( .A(blockdata[125]), .Y(n1460) );
  CLKINVX1 U1438 ( .A(blockdata[62]), .Y(n1397) );
  CLKINVX1 U1439 ( .A(blockdata[126]), .Y(n1461) );
  CLKINVX1 U1440 ( .A(blockdata[63]), .Y(n1398) );
  CLKINVX1 U1441 ( .A(blockdata[127]), .Y(n1462) );
  CLKINVX1 U1442 ( .A(blockdata[0]), .Y(n1335) );
  CLKINVX1 U1443 ( .A(blockdata[1]), .Y(n1336) );
  CLKINVX1 U1444 ( .A(blockdata[2]), .Y(n1337) );
  CLKINVX1 U1445 ( .A(blockdata[3]), .Y(n1338) );
  CLKINVX1 U1446 ( .A(blockdata[4]), .Y(n1339) );
  CLKINVX1 U1447 ( .A(blockdata[5]), .Y(n1340) );
  CLKINVX1 U1448 ( .A(blockdata[6]), .Y(n1341) );
  CLKINVX1 U1449 ( .A(blockdata[7]), .Y(n1342) );
  CLKINVX1 U1450 ( .A(blockdata[8]), .Y(n1343) );
  CLKINVX1 U1451 ( .A(blockdata[9]), .Y(n1344) );
  CLKINVX1 U1452 ( .A(blockdata[10]), .Y(n1345) );
  CLKINVX1 U1453 ( .A(blockdata[11]), .Y(n1346) );
  CLKINVX1 U1454 ( .A(blockdata[12]), .Y(n1347) );
  CLKINVX1 U1455 ( .A(blockdata[13]), .Y(n1348) );
  CLKINVX1 U1456 ( .A(blockdata[14]), .Y(n1349) );
  CLKINVX1 U1457 ( .A(blockdata[15]), .Y(n1350) );
  CLKINVX1 U1458 ( .A(blockdata[16]), .Y(n1351) );
  CLKINVX1 U1459 ( .A(blockdata[17]), .Y(n1352) );
  CLKINVX1 U1460 ( .A(blockdata[18]), .Y(n1353) );
  CLKINVX1 U1461 ( .A(blockdata[19]), .Y(n1354) );
  CLKINVX1 U1462 ( .A(blockdata[20]), .Y(n1355) );
  CLKINVX1 U1463 ( .A(blockdata[21]), .Y(n1356) );
  CLKINVX1 U1464 ( .A(blockdata[22]), .Y(n1357) );
  CLKINVX1 U1465 ( .A(blockdata[23]), .Y(n1358) );
  CLKINVX1 U1466 ( .A(blockdata[24]), .Y(n1359) );
  CLKINVX1 U1467 ( .A(blockdata[25]), .Y(n1360) );
  CLKINVX1 U1468 ( .A(blockdata[26]), .Y(n1361) );
  CLKINVX1 U1469 ( .A(blockdata[27]), .Y(n1362) );
  CLKINVX1 U1470 ( .A(blockdata[28]), .Y(n1363) );
  CLKINVX1 U1471 ( .A(blockdata[29]), .Y(n1364) );
  CLKINVX1 U1472 ( .A(blockdata[30]), .Y(n1365) );
  CLKINVX1 U1473 ( .A(blockdata[31]), .Y(n1366) );
  CLKINVX1 U1474 ( .A(n503), .Y(n1511) );
  CLKBUFX3 U1475 ( .A(N965), .Y(n1237) );
  CLKBUFX3 U1476 ( .A(N960), .Y(n1271) );
  CLKBUFX3 U1477 ( .A(N957), .Y(n1288) );
  CLKBUFX3 U1478 ( .A(N962), .Y(n1254) );
  CLKBUFX3 U1479 ( .A(n695), .Y(n1247) );
  CLKBUFX3 U1480 ( .A(n696), .Y(n1264) );
  CLKINVX1 U1481 ( .A(n22), .Y(n1466) );
  CLKINVX1 U1482 ( .A(n26), .Y(n1469) );
  CLKINVX1 U1483 ( .A(n30), .Y(n1471) );
  CLKINVX1 U1484 ( .A(n18), .Y(n1464) );
  MXI2X1 U1485 ( .A(n1055), .B(n1056), .S0(n1160), .Y(tag[19]) );
  MXI4X1 U1486 ( .A(\blocktag[0][19] ), .B(\blocktag[1][19] ), .C(
        \blocktag[2][19] ), .D(\blocktag[3][19] ), .S0(n1106), .S1(n1134), .Y(
        n1055) );
  MXI4X1 U1487 ( .A(\blocktag[4][19] ), .B(\blocktag[5][19] ), .C(
        \blocktag[6][19] ), .D(\blocktag[7][19] ), .S0(n1106), .S1(n1134), .Y(
        n1056) );
  MXI2X1 U1488 ( .A(n1093), .B(n1094), .S0(n1163), .Y(tag[0]) );
  MXI4X1 U1489 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(
        \blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n1103), .S1(n1131), .Y(
        n1093) );
  MXI4X1 U1490 ( .A(\blocktag[4][0] ), .B(\blocktag[5][0] ), .C(
        \blocktag[6][0] ), .D(\blocktag[7][0] ), .S0(n1103), .S1(n1131), .Y(
        n1094) );
  MXI2X1 U1491 ( .A(n1091), .B(n1092), .S0(n1163), .Y(tag[1]) );
  MXI4X1 U1492 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(
        \blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n1103), .S1(n1131), .Y(
        n1091) );
  MXI4X1 U1493 ( .A(\blocktag[4][1] ), .B(\blocktag[5][1] ), .C(
        \blocktag[6][1] ), .D(\blocktag[7][1] ), .S0(n1103), .S1(n1131), .Y(
        n1092) );
  MXI2X1 U1494 ( .A(n1087), .B(n1088), .S0(n1163), .Y(tag[3]) );
  MXI4X1 U1495 ( .A(\blocktag[0][3] ), .B(\blocktag[1][3] ), .C(
        \blocktag[2][3] ), .D(\blocktag[3][3] ), .S0(n1103), .S1(n1131), .Y(
        n1087) );
  MXI4X1 U1496 ( .A(\blocktag[4][3] ), .B(\blocktag[5][3] ), .C(
        \blocktag[6][3] ), .D(\blocktag[7][3] ), .S0(n1103), .S1(n1131), .Y(
        n1088) );
  MXI2X1 U1497 ( .A(n1077), .B(n1078), .S0(n1163), .Y(tag[8]) );
  MXI4X1 U1498 ( .A(\blocktag[0][8] ), .B(\blocktag[1][8] ), .C(
        \blocktag[2][8] ), .D(\blocktag[3][8] ), .S0(n687), .S1(n1132), .Y(
        n1077) );
  MXI4X1 U1499 ( .A(\blocktag[4][8] ), .B(\blocktag[5][8] ), .C(
        \blocktag[6][8] ), .D(\blocktag[7][8] ), .S0(n688), .S1(n1132), .Y(
        n1078) );
  MXI2X1 U1500 ( .A(n1069), .B(n1070), .S0(n1160), .Y(tag[12]) );
  MXI4X1 U1501 ( .A(\blocktag[0][12] ), .B(\blocktag[1][12] ), .C(
        \blocktag[2][12] ), .D(\blocktag[3][12] ), .S0(n1105), .S1(n1133), .Y(
        n1069) );
  MXI4X1 U1502 ( .A(\blocktag[4][12] ), .B(\blocktag[5][12] ), .C(
        \blocktag[6][12] ), .D(\blocktag[7][12] ), .S0(n1105), .S1(n1133), .Y(
        n1070) );
  MXI2X1 U1503 ( .A(n1083), .B(n1084), .S0(n1163), .Y(tag[5]) );
  MXI2X1 U1504 ( .A(n1079), .B(n1080), .S0(n1163), .Y(tag[7]) );
  MXI2X1 U1505 ( .A(n1061), .B(n1062), .S0(n1160), .Y(tag[16]) );
  MXI2X1 U1506 ( .A(n1085), .B(n1086), .S0(n1163), .Y(tag[4]) );
  MXI2X1 U1507 ( .A(n1043), .B(n1044), .S0(n1164), .Y(dirty) );
  MXI2X1 U1508 ( .A(n1041), .B(n1042), .S0(n1164), .Y(valid) );
  NAND3X1 U1509 ( .A(n485), .B(n486), .C(n487), .Y(n481) );
  XNOR2X1 U1510 ( .A(dataTag[12]), .B(n693), .Y(n485) );
  XNOR2X1 U1511 ( .A(dataTag[8]), .B(n690), .Y(n487) );
  XNOR2X1 U1512 ( .A(dataTag[20]), .B(tag[20]), .Y(n486) );
  XOR2X1 U1513 ( .A(n689), .B(dataTag[21]), .Y(n477) );
  XOR2X1 U1514 ( .A(tag[17]), .B(dataTag[17]), .Y(n484) );
  XOR2X1 U1515 ( .A(tag[6]), .B(dataTag[6]), .Y(n499) );
  NOR3BXL U1516 ( .AN(state[0]), .B(state[2]), .C(n1510), .Y(state_next[2]) );
  XOR2X1 U1517 ( .A(tag[22]), .B(dataTag[22]), .Y(n476) );
  XOR2X1 U1518 ( .A(tag[7]), .B(dataTag[7]), .Y(n483) );
  XOR2X1 U1519 ( .A(tag[2]), .B(dataTag[2]), .Y(n498) );
  XOR2X1 U1520 ( .A(tag[23]), .B(dataTag[23]), .Y(n475) );
  XOR2X1 U1521 ( .A(n692), .B(dataTag[4]), .Y(n497) );
  XNOR2X1 U1522 ( .A(dataTag[19]), .B(n694), .Y(n495) );
  NOR4X1 U1523 ( .A(n488), .B(n489), .C(n490), .D(n491), .Y(n471) );
  XOR2X1 U1524 ( .A(tag[18]), .B(dataTag[18]), .Y(n489) );
  XOR2X1 U1525 ( .A(tag[24]), .B(dataTag[24]), .Y(n490) );
  XOR2X1 U1526 ( .A(n691), .B(dataTag[5]), .Y(n491) );
  NAND4X1 U1527 ( .A(n492), .B(n493), .C(n494), .D(n495), .Y(n488) );
  XNOR2X1 U1528 ( .A(dataTag[9]), .B(tag[9]), .Y(n494) );
  NAND4X1 U1529 ( .A(n478), .B(n479), .C(n480), .D(valid), .Y(n474) );
  XNOR2X1 U1530 ( .A(dataTag[3]), .B(n685), .Y(n478) );
  XNOR2X1 U1531 ( .A(dataTag[1]), .B(n684), .Y(n479) );
  XNOR2X1 U1532 ( .A(dataTag[0]), .B(n683), .Y(n480) );
  NAND3X1 U1533 ( .A(state_next[2]), .B(n1308), .C(proc_write_r), .Y(n34) );
  OAI21XL U1534 ( .A0(mem_ready_r), .A1(n1509), .B0(n63), .Y(mem_read_next) );
  OAI2BB2XL U1535 ( .B0(mem_ready_r), .B1(n9), .A0N(n10), .A1N(dirty), .Y(n7)
         );
  NAND3X1 U1536 ( .A(n500), .B(n501), .C(n502), .Y(n496) );
  XNOR2X1 U1537 ( .A(dataTag[11]), .B(tag[11]), .Y(n500) );
  XNOR2X1 U1538 ( .A(dataTag[13]), .B(tag[13]), .Y(n502) );
  XNOR2X1 U1539 ( .A(dataTag[10]), .B(tag[10]), .Y(n501) );
  OAI21XL U1540 ( .A0(proc_write_r), .A1(n1308), .B0(n10), .Y(n465) );
  AOI222XL U1541 ( .A0(mem_addr[3]), .A1(n1221), .B0(n38), .B1(dataTag[0]), 
        .C0(n683), .C1(n1173), .Y(n39) );
  AOI222XL U1542 ( .A0(mem_addr[4]), .A1(n1221), .B0(n38), .B1(dataTag[1]), 
        .C0(n684), .C1(n1173), .Y(n40) );
  AOI222XL U1543 ( .A0(mem_addr[5]), .A1(n1220), .B0(n38), .B1(dataTag[2]), 
        .C0(tag[2]), .C1(n1173), .Y(n41) );
  AOI222XL U1544 ( .A0(mem_addr[6]), .A1(n1221), .B0(n38), .B1(dataTag[3]), 
        .C0(n685), .C1(n1173), .Y(n42) );
  AOI222XL U1545 ( .A0(mem_addr[7]), .A1(n1220), .B0(n38), .B1(dataTag[4]), 
        .C0(n692), .C1(n1173), .Y(n43) );
  AOI222XL U1546 ( .A0(mem_addr[8]), .A1(n1220), .B0(n38), .B1(dataTag[5]), 
        .C0(n691), .C1(n1173), .Y(n44) );
  AOI222XL U1547 ( .A0(mem_addr[9]), .A1(n1220), .B0(n38), .B1(dataTag[6]), 
        .C0(tag[6]), .C1(n1173), .Y(n45) );
  AOI222XL U1548 ( .A0(mem_addr[10]), .A1(n1220), .B0(n38), .B1(dataTag[7]), 
        .C0(tag[7]), .C1(n1173), .Y(n46) );
  AOI222XL U1549 ( .A0(mem_addr[11]), .A1(n1221), .B0(n38), .B1(dataTag[8]), 
        .C0(n690), .C1(n1173), .Y(n47) );
  AOI222XL U1550 ( .A0(mem_addr[12]), .A1(n1220), .B0(n38), .B1(dataTag[9]), 
        .C0(tag[9]), .C1(n1173), .Y(n48) );
  AOI222XL U1551 ( .A0(mem_addr[13]), .A1(n1220), .B0(n38), .B1(dataTag[10]), 
        .C0(tag[10]), .C1(n1173), .Y(n49) );
  AOI222XL U1552 ( .A0(mem_addr[14]), .A1(n1220), .B0(n38), .B1(dataTag[11]), 
        .C0(tag[11]), .C1(n1174), .Y(n50) );
  AOI222XL U1553 ( .A0(mem_addr[15]), .A1(n1220), .B0(n38), .B1(dataTag[12]), 
        .C0(n693), .C1(n1174), .Y(n51) );
  AOI222XL U1554 ( .A0(mem_addr[16]), .A1(n1220), .B0(n38), .B1(dataTag[13]), 
        .C0(tag[13]), .C1(n1174), .Y(n52) );
  AOI222XL U1555 ( .A0(mem_addr[19]), .A1(n1220), .B0(n38), .B1(dataTag[16]), 
        .C0(tag[16]), .C1(n1174), .Y(n55) );
  AOI222XL U1556 ( .A0(mem_addr[20]), .A1(n1220), .B0(n38), .B1(dataTag[17]), 
        .C0(tag[17]), .C1(n1174), .Y(n56) );
  AOI222XL U1557 ( .A0(mem_addr[21]), .A1(n1220), .B0(n38), .B1(dataTag[18]), 
        .C0(tag[18]), .C1(n1174), .Y(n57) );
  AOI222XL U1558 ( .A0(mem_addr[22]), .A1(n1220), .B0(n38), .B1(dataTag[19]), 
        .C0(n694), .C1(n1174), .Y(n58) );
  AOI222XL U1559 ( .A0(mem_addr[23]), .A1(n1220), .B0(n38), .B1(dataTag[20]), 
        .C0(tag[20]), .C1(n1174), .Y(n59) );
  AOI222XL U1560 ( .A0(mem_addr[24]), .A1(n1220), .B0(n38), .B1(dataTag[21]), 
        .C0(n689), .C1(n1174), .Y(n60) );
  AOI222XL U1561 ( .A0(mem_addr[25]), .A1(n1220), .B0(n38), .B1(dataTag[22]), 
        .C0(tag[22]), .C1(n1174), .Y(n61) );
  AOI222XL U1562 ( .A0(mem_addr[26]), .A1(n1221), .B0(n38), .B1(dataTag[23]), 
        .C0(tag[23]), .C1(n1173), .Y(n62) );
  CLKINVX1 U1563 ( .A(n1222), .Y(n1221) );
  OR4X1 U1564 ( .A(n66), .B(n67), .C(n68), .D(n69), .Y(n651) );
  OAI22XL U1565 ( .A0(n1201), .A1(n1431), .B0(n1198), .B1(n1335), .Y(n66) );
  OAI22XL U1566 ( .A0(n1217), .A1(n1367), .B0(n1214), .B1(n1575), .Y(n69) );
  OAI2BB2XL U1567 ( .B0(n1204), .B1(n1399), .A0N(proc_rdata[0]), .A1N(n1172), 
        .Y(n67) );
  OR4X1 U1568 ( .A(n87), .B(n88), .C(n89), .D(n90), .Y(n652) );
  OAI22XL U1569 ( .A0(n1201), .A1(n1432), .B0(n1198), .B1(n1336), .Y(n87) );
  OAI22XL U1570 ( .A0(n1217), .A1(n1368), .B0(n1214), .B1(n1574), .Y(n90) );
  OAI2BB2XL U1571 ( .B0(n1204), .B1(n1400), .A0N(proc_rdata[1]), .A1N(n1172), 
        .Y(n88) );
  OR4X1 U1572 ( .A(n99), .B(n100), .C(n101), .D(n102), .Y(n653) );
  OAI22XL U1573 ( .A0(n1201), .A1(n1433), .B0(n1198), .B1(n1337), .Y(n99) );
  OAI22XL U1574 ( .A0(n1217), .A1(n1369), .B0(n1214), .B1(n1573), .Y(n102) );
  OAI2BB2XL U1575 ( .B0(n1204), .B1(n1401), .A0N(proc_rdata[2]), .A1N(n1172), 
        .Y(n100) );
  OR4X1 U1576 ( .A(n111), .B(n112), .C(n113), .D(n114), .Y(n654) );
  OAI22XL U1577 ( .A0(n1201), .A1(n1434), .B0(n1198), .B1(n1338), .Y(n111) );
  OAI22XL U1578 ( .A0(n1217), .A1(n1370), .B0(n1214), .B1(n1572), .Y(n114) );
  OAI2BB2XL U1579 ( .B0(n1204), .B1(n1402), .A0N(proc_rdata[3]), .A1N(n1172), 
        .Y(n112) );
  OR4X1 U1580 ( .A(n123), .B(n124), .C(n125), .D(n126), .Y(n655) );
  OAI22XL U1581 ( .A0(n1201), .A1(n1435), .B0(n1198), .B1(n1339), .Y(n123) );
  OAI22XL U1582 ( .A0(n1217), .A1(n1371), .B0(n1214), .B1(n1571), .Y(n126) );
  OAI2BB2XL U1583 ( .B0(n1204), .B1(n1403), .A0N(proc_rdata[4]), .A1N(n1172), 
        .Y(n124) );
  OR4X1 U1584 ( .A(n135), .B(n136), .C(n137), .D(n138), .Y(n656) );
  OAI22XL U1585 ( .A0(n1201), .A1(n1436), .B0(n1198), .B1(n1340), .Y(n135) );
  OAI22XL U1586 ( .A0(n1217), .A1(n1372), .B0(n1214), .B1(n1570), .Y(n138) );
  OAI2BB2XL U1587 ( .B0(n1204), .B1(n1404), .A0N(proc_rdata[5]), .A1N(n1172), 
        .Y(n136) );
  OR4X1 U1588 ( .A(n147), .B(n148), .C(n149), .D(n150), .Y(n657) );
  OAI22XL U1589 ( .A0(n1201), .A1(n1437), .B0(n1198), .B1(n1341), .Y(n147) );
  OAI22XL U1590 ( .A0(n1217), .A1(n1373), .B0(n1214), .B1(n1569), .Y(n150) );
  OAI2BB2XL U1591 ( .B0(n1204), .B1(n1405), .A0N(proc_rdata[6]), .A1N(n1172), 
        .Y(n148) );
  OR4X1 U1592 ( .A(n159), .B(n160), .C(n161), .D(n162), .Y(n658) );
  OAI22XL U1593 ( .A0(n1201), .A1(n1438), .B0(n1198), .B1(n1342), .Y(n159) );
  OAI22XL U1594 ( .A0(n1217), .A1(n1374), .B0(n1214), .B1(n1568), .Y(n162) );
  OAI2BB2XL U1595 ( .B0(n1204), .B1(n1406), .A0N(proc_rdata[7]), .A1N(n1172), 
        .Y(n160) );
  OR4X1 U1596 ( .A(n171), .B(n172), .C(n173), .D(n174), .Y(n659) );
  OAI22XL U1597 ( .A0(n1201), .A1(n1439), .B0(n1198), .B1(n1343), .Y(n171) );
  OAI22XL U1598 ( .A0(n1217), .A1(n1375), .B0(n1214), .B1(n1567), .Y(n174) );
  OAI2BB2XL U1599 ( .B0(n1204), .B1(n1407), .A0N(proc_rdata[8]), .A1N(n1171), 
        .Y(n172) );
  OR4X1 U1600 ( .A(n183), .B(n184), .C(n185), .D(n186), .Y(n660) );
  OAI22XL U1601 ( .A0(n1201), .A1(n1440), .B0(n1198), .B1(n1344), .Y(n183) );
  OAI22XL U1602 ( .A0(n1217), .A1(n1376), .B0(n1214), .B1(n1566), .Y(n186) );
  OAI2BB2XL U1603 ( .B0(n1204), .B1(n1408), .A0N(proc_rdata[9]), .A1N(n1171), 
        .Y(n184) );
  OR4X1 U1604 ( .A(n195), .B(n196), .C(n197), .D(n198), .Y(n661) );
  OAI22XL U1605 ( .A0(n1201), .A1(n1441), .B0(n1198), .B1(n1345), .Y(n195) );
  OAI22XL U1606 ( .A0(n1217), .A1(n1377), .B0(n1214), .B1(n1565), .Y(n198) );
  OAI2BB2XL U1607 ( .B0(n1204), .B1(n1409), .A0N(proc_rdata[10]), .A1N(n1171), 
        .Y(n196) );
  OR4X1 U1608 ( .A(n207), .B(n208), .C(n209), .D(n210), .Y(n662) );
  OAI22XL U1609 ( .A0(n1201), .A1(n1442), .B0(n1198), .B1(n1346), .Y(n207) );
  OAI22XL U1610 ( .A0(n1217), .A1(n1378), .B0(n1214), .B1(n1564), .Y(n210) );
  OAI2BB2XL U1611 ( .B0(n1204), .B1(n1410), .A0N(proc_rdata[11]), .A1N(n1171), 
        .Y(n208) );
  OR4X1 U1612 ( .A(n219), .B(n220), .C(n221), .D(n222), .Y(n663) );
  OAI22XL U1613 ( .A0(n1202), .A1(n1443), .B0(n1199), .B1(n1347), .Y(n219) );
  OAI22XL U1614 ( .A0(n1218), .A1(n1379), .B0(n1215), .B1(n1563), .Y(n222) );
  OAI2BB2XL U1615 ( .B0(n1205), .B1(n1411), .A0N(proc_rdata[12]), .A1N(n1171), 
        .Y(n220) );
  OR4X1 U1616 ( .A(n231), .B(n232), .C(n233), .D(n234), .Y(n664) );
  OAI22XL U1617 ( .A0(n1202), .A1(n1444), .B0(n1199), .B1(n1348), .Y(n231) );
  OAI22XL U1618 ( .A0(n1218), .A1(n1380), .B0(n1215), .B1(n1562), .Y(n234) );
  OAI2BB2XL U1619 ( .B0(n1205), .B1(n1412), .A0N(proc_rdata[13]), .A1N(n1171), 
        .Y(n232) );
  OR4X1 U1620 ( .A(n243), .B(n244), .C(n245), .D(n246), .Y(n665) );
  OAI22XL U1621 ( .A0(n1202), .A1(n1445), .B0(n1199), .B1(n1349), .Y(n243) );
  OAI22XL U1622 ( .A0(n1218), .A1(n1381), .B0(n1215), .B1(n1561), .Y(n246) );
  OAI2BB2XL U1623 ( .B0(n1205), .B1(n1413), .A0N(proc_rdata[14]), .A1N(n1171), 
        .Y(n244) );
  OR4X1 U1624 ( .A(n255), .B(n256), .C(n257), .D(n258), .Y(n666) );
  OAI22XL U1625 ( .A0(n1202), .A1(n1446), .B0(n1199), .B1(n1350), .Y(n255) );
  OAI22XL U1626 ( .A0(n1218), .A1(n1382), .B0(n1215), .B1(n1560), .Y(n258) );
  OAI2BB2XL U1627 ( .B0(n1205), .B1(n1414), .A0N(proc_rdata[15]), .A1N(n1171), 
        .Y(n256) );
  OR4X1 U1628 ( .A(n267), .B(n268), .C(n269), .D(n270), .Y(n667) );
  OAI22XL U1629 ( .A0(n1202), .A1(n1447), .B0(n1199), .B1(n1351), .Y(n267) );
  OAI22XL U1630 ( .A0(n1218), .A1(n1383), .B0(n1215), .B1(n1559), .Y(n270) );
  OAI2BB2XL U1631 ( .B0(n1205), .B1(n1415), .A0N(proc_rdata[16]), .A1N(n1171), 
        .Y(n268) );
  OR4X1 U1632 ( .A(n279), .B(n280), .C(n281), .D(n282), .Y(n668) );
  OAI22XL U1633 ( .A0(n1202), .A1(n1448), .B0(n1199), .B1(n1352), .Y(n279) );
  OAI22XL U1634 ( .A0(n1218), .A1(n1384), .B0(n1215), .B1(n1558), .Y(n282) );
  OAI2BB2XL U1635 ( .B0(n1205), .B1(n1416), .A0N(proc_rdata[17]), .A1N(n1171), 
        .Y(n280) );
  OR4X1 U1636 ( .A(n291), .B(n292), .C(n293), .D(n294), .Y(n669) );
  OAI22XL U1637 ( .A0(n1202), .A1(n1449), .B0(n1199), .B1(n1353), .Y(n291) );
  OAI22XL U1638 ( .A0(n1218), .A1(n1385), .B0(n1215), .B1(n1557), .Y(n294) );
  OAI2BB2XL U1639 ( .B0(n1205), .B1(n1417), .A0N(proc_rdata[18]), .A1N(n1171), 
        .Y(n292) );
  OR4X1 U1640 ( .A(n303), .B(n304), .C(n305), .D(n306), .Y(n670) );
  OAI22XL U1641 ( .A0(n1202), .A1(n1450), .B0(n1199), .B1(n1354), .Y(n303) );
  OAI22XL U1642 ( .A0(n1218), .A1(n1386), .B0(n1215), .B1(n1556), .Y(n306) );
  OAI2BB2XL U1643 ( .B0(n1205), .B1(n1418), .A0N(proc_rdata[19]), .A1N(n1171), 
        .Y(n304) );
  OR4X1 U1644 ( .A(n315), .B(n316), .C(n317), .D(n318), .Y(n671) );
  OAI22XL U1645 ( .A0(n1202), .A1(n1451), .B0(n1199), .B1(n1355), .Y(n315) );
  OAI22XL U1646 ( .A0(n1218), .A1(n1387), .B0(n1215), .B1(n1555), .Y(n318) );
  OAI2BB2XL U1647 ( .B0(n1205), .B1(n1419), .A0N(proc_rdata[20]), .A1N(n1170), 
        .Y(n316) );
  OR4X1 U1648 ( .A(n327), .B(n328), .C(n329), .D(n330), .Y(n672) );
  OAI22XL U1649 ( .A0(n1202), .A1(n1452), .B0(n1199), .B1(n1356), .Y(n327) );
  OAI22XL U1650 ( .A0(n1218), .A1(n1388), .B0(n1215), .B1(n1554), .Y(n330) );
  OAI2BB2XL U1651 ( .B0(n1205), .B1(n1420), .A0N(proc_rdata[21]), .A1N(n1170), 
        .Y(n328) );
  OR4X1 U1652 ( .A(n339), .B(n340), .C(n341), .D(n342), .Y(n673) );
  OAI22XL U1653 ( .A0(n1202), .A1(n1453), .B0(n1199), .B1(n1357), .Y(n339) );
  OAI22XL U1654 ( .A0(n1218), .A1(n1389), .B0(n1215), .B1(n1553), .Y(n342) );
  OAI2BB2XL U1655 ( .B0(n1205), .B1(n1421), .A0N(proc_rdata[22]), .A1N(n1170), 
        .Y(n340) );
  OR4X1 U1656 ( .A(n351), .B(n352), .C(n353), .D(n354), .Y(n674) );
  OAI22XL U1657 ( .A0(n1202), .A1(n1454), .B0(n1199), .B1(n1358), .Y(n351) );
  OAI22XL U1658 ( .A0(n1218), .A1(n1390), .B0(n1215), .B1(n1552), .Y(n354) );
  OAI2BB2XL U1659 ( .B0(n1205), .B1(n1422), .A0N(proc_rdata[23]), .A1N(n1170), 
        .Y(n352) );
  OR4X1 U1660 ( .A(n363), .B(n364), .C(n365), .D(n366), .Y(n675) );
  OAI22XL U1661 ( .A0(n1203), .A1(n1455), .B0(n1200), .B1(n1359), .Y(n363) );
  OAI22XL U1662 ( .A0(n1219), .A1(n1391), .B0(n1216), .B1(n1551), .Y(n366) );
  OAI2BB2XL U1663 ( .B0(n1206), .B1(n1423), .A0N(proc_rdata[24]), .A1N(n1170), 
        .Y(n364) );
  OR4X1 U1664 ( .A(n375), .B(n376), .C(n377), .D(n378), .Y(n676) );
  OAI22XL U1665 ( .A0(n1203), .A1(n1456), .B0(n1200), .B1(n1360), .Y(n375) );
  OAI22XL U1666 ( .A0(n1219), .A1(n1392), .B0(n1216), .B1(n1550), .Y(n378) );
  OAI2BB2XL U1667 ( .B0(n1206), .B1(n1424), .A0N(proc_rdata[25]), .A1N(n1170), 
        .Y(n376) );
  OR4X1 U1668 ( .A(n387), .B(n388), .C(n389), .D(n390), .Y(n677) );
  OAI22XL U1669 ( .A0(n1203), .A1(n1457), .B0(n1200), .B1(n1361), .Y(n387) );
  OAI22XL U1670 ( .A0(n1219), .A1(n1393), .B0(n1216), .B1(n1549), .Y(n390) );
  OAI2BB2XL U1671 ( .B0(n1206), .B1(n1425), .A0N(proc_rdata[26]), .A1N(n1170), 
        .Y(n388) );
  OR4X1 U1672 ( .A(n399), .B(n400), .C(n401), .D(n402), .Y(n678) );
  OAI22XL U1673 ( .A0(n1203), .A1(n1458), .B0(n1200), .B1(n1362), .Y(n399) );
  OAI22XL U1674 ( .A0(n1219), .A1(n1394), .B0(n1216), .B1(n1548), .Y(n402) );
  OAI2BB2XL U1675 ( .B0(n1206), .B1(n1426), .A0N(proc_rdata[27]), .A1N(n1170), 
        .Y(n400) );
  OR4X1 U1676 ( .A(n411), .B(n412), .C(n413), .D(n414), .Y(n679) );
  OAI22XL U1677 ( .A0(n1203), .A1(n1459), .B0(n1200), .B1(n1363), .Y(n411) );
  OAI22XL U1678 ( .A0(n1219), .A1(n1395), .B0(n1216), .B1(n1547), .Y(n414) );
  OAI2BB2XL U1679 ( .B0(n1206), .B1(n1427), .A0N(proc_rdata[28]), .A1N(n1170), 
        .Y(n412) );
  OR4X1 U1680 ( .A(n423), .B(n424), .C(n425), .D(n426), .Y(n680) );
  OAI22XL U1681 ( .A0(n1203), .A1(n1460), .B0(n1200), .B1(n1364), .Y(n423) );
  OAI22XL U1682 ( .A0(n1219), .A1(n1396), .B0(n1216), .B1(n1546), .Y(n426) );
  OAI2BB2XL U1683 ( .B0(n1206), .B1(n1428), .A0N(proc_rdata[29]), .A1N(n1170), 
        .Y(n424) );
  OR4X1 U1684 ( .A(n435), .B(n436), .C(n437), .D(n438), .Y(n681) );
  OAI22XL U1685 ( .A0(n1203), .A1(n1461), .B0(n1200), .B1(n1365), .Y(n435) );
  OAI22XL U1686 ( .A0(n1219), .A1(n1397), .B0(n1216), .B1(n1545), .Y(n438) );
  OAI2BB2XL U1687 ( .B0(n1206), .B1(n1429), .A0N(proc_rdata[30]), .A1N(n1170), 
        .Y(n436) );
  OR4X1 U1688 ( .A(n447), .B(n448), .C(n449), .D(n450), .Y(n682) );
  OAI22XL U1689 ( .A0(n1203), .A1(n1462), .B0(n1200), .B1(n1366), .Y(n447) );
  OAI22XL U1690 ( .A0(n1219), .A1(n1398), .B0(n1216), .B1(n1544), .Y(n450) );
  OAI2BB2XL U1691 ( .B0(n1206), .B1(n1430), .A0N(proc_rdata[31]), .A1N(n1170), 
        .Y(n448) );
  CLKINVX1 U1692 ( .A(N87), .Y(n1467) );
  NOR2X2 U1693 ( .A(n1475), .B(wordIndex[1]), .Y(n456) );
  NOR2X2 U1694 ( .A(n1474), .B(wordIndex[0]), .Y(n455) );
  OAI21X1 U1695 ( .A0(state[2]), .A1(state[0]), .B0(n1511), .Y(n11) );
  AO22X2 U1696 ( .A0(dataTag[0]), .A1(n1236), .B0(n1233), .B1(n683), .Y(
        blocktag_next[0]) );
  AO22X2 U1697 ( .A0(dataTag[10]), .A1(n1234), .B0(n1230), .B1(tag[10]), .Y(
        blocktag_next[10]) );
  AO22X2 U1698 ( .A0(dataTag[11]), .A1(n1234), .B0(n1233), .B1(tag[11]), .Y(
        blocktag_next[11]) );
  AO22X2 U1699 ( .A0(dataTag[12]), .A1(n1235), .B0(n1233), .B1(n693), .Y(
        blocktag_next[12]) );
  AO22X2 U1700 ( .A0(dataTag[13]), .A1(n1236), .B0(n1233), .B1(tag[13]), .Y(
        blocktag_next[13]) );
  AO22X2 U1701 ( .A0(dataTag[14]), .A1(n1236), .B0(n1231), .B1(n699), .Y(
        blocktag_next[14]) );
  AO22X2 U1702 ( .A0(dataTag[15]), .A1(n1236), .B0(n1233), .B1(n700), .Y(
        blocktag_next[15]) );
  AO22X2 U1703 ( .A0(dataTag[19]), .A1(n1236), .B0(n1233), .B1(n694), .Y(
        blocktag_next[19]) );
  AO22X2 U1704 ( .A0(dataTag[1]), .A1(n1236), .B0(n1229), .B1(n684), .Y(
        blocktag_next[1]) );
  AO22X2 U1705 ( .A0(dataTag[20]), .A1(n1236), .B0(n1233), .B1(tag[20]), .Y(
        blocktag_next[20]) );
  AO22X2 U1706 ( .A0(dataTag[3]), .A1(n1236), .B0(n1233), .B1(n685), .Y(
        blocktag_next[3]) );
  AO22X2 U1707 ( .A0(dataTag[8]), .A1(n1236), .B0(n1228), .B1(n690), .Y(
        blocktag_next[8]) );
  AO22X2 U1708 ( .A0(dataTag[9]), .A1(n1236), .B0(n1227), .B1(tag[9]), .Y(
        blocktag_next[9]) );
  AO22X2 U1709 ( .A0(n1233), .A1(tag[16]), .B0(dataTag[16]), .B1(n1236), .Y(
        blocktag_next[16]) );
  AO22X2 U1710 ( .A0(n1233), .A1(tag[17]), .B0(dataTag[17]), .B1(n1224), .Y(
        blocktag_next[17]) );
  AO22X2 U1711 ( .A0(n1233), .A1(tag[18]), .B0(dataTag[18]), .B1(n1234), .Y(
        blocktag_next[18]) );
  AO22X2 U1712 ( .A0(n1233), .A1(n689), .B0(dataTag[21]), .B1(n1236), .Y(
        blocktag_next[21]) );
  AO22X2 U1713 ( .A0(n1233), .A1(tag[22]), .B0(dataTag[22]), .B1(n1225), .Y(
        blocktag_next[22]) );
  AO22X2 U1714 ( .A0(n1233), .A1(tag[23]), .B0(dataTag[23]), .B1(n1236), .Y(
        blocktag_next[23]) );
  AO22X2 U1715 ( .A0(n1233), .A1(tag[24]), .B0(dataTag[24]), .B1(n1236), .Y(
        blocktag_next[24]) );
  AO22X2 U1716 ( .A0(n1233), .A1(tag[2]), .B0(dataTag[2]), .B1(n1236), .Y(
        blocktag_next[2]) );
  AO22X2 U1717 ( .A0(n1233), .A1(n692), .B0(dataTag[4]), .B1(n1225), .Y(
        blocktag_next[4]) );
  AO22X2 U1718 ( .A0(n1233), .A1(n691), .B0(dataTag[5]), .B1(n33), .Y(
        blocktag_next[5]) );
  AO22X2 U1719 ( .A0(n1233), .A1(tag[6]), .B0(dataTag[6]), .B1(n33), .Y(
        blocktag_next[6]) );
  AO22X2 U1720 ( .A0(n1233), .A1(tag[7]), .B0(dataTag[7]), .B1(n33), .Y(
        blocktag_next[7]) );
  NAND2X1 U1721 ( .A(n554), .B(N85), .Y(n22) );
  NAND2X1 U1722 ( .A(n555), .B(N85), .Y(n26) );
  NAND2X1 U1723 ( .A(n556), .B(N85), .Y(n30) );
  NAND2X1 U1724 ( .A(N85), .B(n550), .Y(n18) );
  NOR2X1 U1725 ( .A(n703), .B(n18), .Y(N965) );
  NOR2X1 U1726 ( .A(n703), .B(n22), .Y(N962) );
  NOR2X1 U1727 ( .A(n703), .B(n26), .Y(N960) );
  NOR2X1 U1728 ( .A(n703), .B(n30), .Y(N957) );
  MXI2X1 U1729 ( .A(n1039), .B(n1040), .S0(n1164), .Y(blockdata[0]) );
  MXI2X1 U1730 ( .A(n1037), .B(n1038), .S0(n1164), .Y(blockdata[1]) );
  MXI2X1 U1731 ( .A(n1035), .B(n1036), .S0(n1164), .Y(blockdata[2]) );
  MXI2X1 U1732 ( .A(n1033), .B(n1034), .S0(n1164), .Y(blockdata[3]) );
  MXI2X1 U1733 ( .A(n1031), .B(n1032), .S0(n1164), .Y(blockdata[4]) );
  MXI4X1 U1734 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n1122), .S1(n1136), .Y(n1032) );
  MXI2X1 U1735 ( .A(n1029), .B(n1030), .S0(n1164), .Y(blockdata[5]) );
  MXI4X1 U1736 ( .A(\block[0][5] ), .B(\block[1][5] ), .C(\block[2][5] ), .D(
        \block[3][5] ), .S0(n1123), .S1(n1136), .Y(n1029) );
  MXI4X1 U1737 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n1115), .S1(n1136), .Y(n1030) );
  MXI2X1 U1738 ( .A(n1027), .B(n1028), .S0(n1164), .Y(blockdata[6]) );
  MXI4X1 U1739 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n1098), .S1(n1136), .Y(n1027) );
  MXI4X1 U1740 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n1119), .S1(n1136), .Y(n1028) );
  MXI2X1 U1741 ( .A(n1025), .B(n1026), .S0(n1164), .Y(blockdata[7]) );
  MXI4X1 U1742 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n1110), .S1(n1136), .Y(n1025) );
  MXI4X1 U1743 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n1121), .S1(n1136), .Y(n1026) );
  MXI2X1 U1744 ( .A(n1023), .B(n1024), .S0(n1165), .Y(blockdata[8]) );
  MXI4X1 U1745 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n1098), .S1(n1137), .Y(n1023) );
  MXI4X1 U1746 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n1099), .S1(n1137), .Y(n1024) );
  MXI2X1 U1747 ( .A(n1021), .B(n1022), .S0(n1165), .Y(blockdata[9]) );
  MXI4X1 U1748 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n1109), .S1(n1137), .Y(n1021) );
  MXI4X1 U1749 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n1115), .S1(n1137), .Y(n1022) );
  MXI2X1 U1750 ( .A(n1019), .B(n1020), .S0(n1165), .Y(blockdata[10]) );
  MXI4X1 U1751 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n1099), .S1(n1137), .Y(n1019) );
  MXI4X1 U1752 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n1120), .S1(n1137), .Y(n1020) );
  MXI2X1 U1753 ( .A(n1017), .B(n1018), .S0(n1165), .Y(blockdata[11]) );
  MXI4X1 U1754 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n1108), .S1(n1137), .Y(n1017) );
  MXI4X1 U1755 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n1108), .S1(n1137), .Y(n1018) );
  MXI2X1 U1756 ( .A(n1015), .B(n1016), .S0(n1165), .Y(blockdata[12]) );
  MXI4X1 U1757 ( .A(\block[0][12] ), .B(\block[1][12] ), .C(\block[2][12] ), 
        .D(\block[3][12] ), .S0(n1108), .S1(n1137), .Y(n1015) );
  MXI4X1 U1758 ( .A(\block[4][12] ), .B(\block[5][12] ), .C(\block[6][12] ), 
        .D(\block[7][12] ), .S0(n1108), .S1(n1137), .Y(n1016) );
  MXI2X1 U1759 ( .A(n1013), .B(n1014), .S0(n1165), .Y(blockdata[13]) );
  MXI4X1 U1760 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n1108), .S1(n1137), .Y(n1013) );
  MXI4X1 U1761 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n1108), .S1(n1137), .Y(n1014) );
  MXI2X1 U1762 ( .A(n1011), .B(n1012), .S0(n1165), .Y(blockdata[14]) );
  MXI4X1 U1763 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n1108), .S1(n1138), .Y(n1011) );
  MXI4X1 U1764 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n1108), .S1(n1138), .Y(n1012) );
  MXI2X1 U1765 ( .A(n1009), .B(n1010), .S0(n1165), .Y(blockdata[15]) );
  MXI4X1 U1766 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n1108), .S1(n1138), .Y(n1009) );
  MXI4X1 U1767 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n1108), .S1(n1138), .Y(n1010) );
  MXI2X1 U1768 ( .A(n1007), .B(n1008), .S0(n1165), .Y(blockdata[16]) );
  MXI4X1 U1769 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n1108), .S1(n1138), .Y(n1007) );
  MXI4X1 U1770 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n1108), .S1(n1138), .Y(n1008) );
  MXI2X1 U1771 ( .A(n1005), .B(n1006), .S0(n1165), .Y(blockdata[17]) );
  MXI4X1 U1772 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n1108), .S1(n1138), .Y(n1005) );
  MXI4X1 U1773 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n1099), .S1(n1138), .Y(n1006) );
  MXI2X1 U1774 ( .A(n1003), .B(n1004), .S0(n1165), .Y(blockdata[18]) );
  MXI4X1 U1775 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n1110), .S1(n1138), .Y(n1003) );
  MXI4X1 U1776 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n1114), .S1(n1138), .Y(n1004) );
  MXI2X1 U1777 ( .A(n1001), .B(n1002), .S0(n1165), .Y(blockdata[19]) );
  MXI4X1 U1778 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n1111), .S1(n1138), .Y(n1001) );
  MXI4X1 U1779 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n1108), .S1(n1138), .Y(n1002) );
  MXI2X1 U1780 ( .A(n999), .B(n1000), .S0(n1166), .Y(blockdata[20]) );
  MXI4X1 U1781 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n1112), .S1(n1139), .Y(n999) );
  MXI4X1 U1782 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n1118), .S1(n1139), .Y(n1000) );
  MXI2X1 U1783 ( .A(n997), .B(n998), .S0(n1166), .Y(blockdata[21]) );
  MXI4X1 U1784 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n1099), .S1(n1139), .Y(n997) );
  MXI4X1 U1785 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n1108), .S1(n1139), .Y(n998) );
  MXI2X1 U1786 ( .A(n995), .B(n996), .S0(n1166), .Y(blockdata[22]) );
  MXI4X1 U1787 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n1113), .S1(n1139), .Y(n995) );
  MXI4X1 U1788 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n1108), .S1(n1139), .Y(n996) );
  MXI2X1 U1789 ( .A(n993), .B(n994), .S0(n1166), .Y(blockdata[23]) );
  MXI4X1 U1790 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n1099), .S1(n1139), .Y(n993) );
  MXI4X1 U1791 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n1109), .S1(n1139), .Y(n994) );
  MXI2X1 U1792 ( .A(n991), .B(n992), .S0(n1166), .Y(blockdata[24]) );
  MXI4X1 U1793 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n1109), .S1(n1139), .Y(n991) );
  MXI4X1 U1794 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n1109), .S1(n1139), .Y(n992) );
  MXI2X1 U1795 ( .A(n989), .B(n990), .S0(n1166), .Y(blockdata[25]) );
  MXI4X1 U1796 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n1109), .S1(n1139), .Y(n989) );
  MXI4X1 U1797 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n1109), .S1(n1139), .Y(n990) );
  MXI2X1 U1798 ( .A(n987), .B(n988), .S0(n1166), .Y(blockdata[26]) );
  MXI4X1 U1799 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n1109), .S1(n1140), .Y(n987) );
  MXI4X1 U1800 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n1109), .S1(n1140), .Y(n988) );
  MXI2X1 U1801 ( .A(n985), .B(n986), .S0(n1166), .Y(blockdata[27]) );
  MXI4X1 U1802 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n1109), .S1(n1140), .Y(n985) );
  MXI4X1 U1803 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n1109), .S1(n1140), .Y(n986) );
  MXI2X1 U1804 ( .A(n983), .B(n984), .S0(n1166), .Y(blockdata[28]) );
  MXI4X1 U1805 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n1109), .S1(n1140), .Y(n983) );
  MXI4X1 U1806 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n1109), .S1(n1140), .Y(n984) );
  MXI2X1 U1807 ( .A(n981), .B(n982), .S0(n1166), .Y(blockdata[29]) );
  MXI4X1 U1808 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n1109), .S1(n1140), .Y(n981) );
  MXI4X1 U1809 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n1109), .S1(n1140), .Y(n982) );
  MXI2X1 U1810 ( .A(n979), .B(n980), .S0(n1166), .Y(blockdata[30]) );
  MXI4X1 U1811 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n1109), .S1(n1140), .Y(n979) );
  MXI4X1 U1812 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n1110), .S1(n1140), .Y(n980) );
  MXI2X1 U1813 ( .A(n977), .B(n978), .S0(n1166), .Y(blockdata[31]) );
  MXI4X1 U1814 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n1110), .S1(n1140), .Y(n977) );
  MXI4X1 U1815 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n1110), .S1(n1140), .Y(n978) );
  MXI2X1 U1816 ( .A(n975), .B(n976), .S0(n1162), .Y(blockdata[32]) );
  MXI4X1 U1817 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n1110), .S1(n1141), .Y(n975) );
  MXI4X1 U1818 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n1110), .S1(n1141), .Y(n976) );
  MXI2X1 U1819 ( .A(n973), .B(n974), .S0(n1160), .Y(blockdata[33]) );
  MXI4X1 U1820 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n1110), .S1(n1141), .Y(n973) );
  MXI4X1 U1821 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n1110), .S1(n1141), .Y(n974) );
  MXI2X1 U1822 ( .A(n971), .B(n972), .S0(n1159), .Y(blockdata[34]) );
  MXI4X1 U1823 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n1110), .S1(n1141), .Y(n971) );
  MXI4X1 U1824 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n1110), .S1(n1141), .Y(n972) );
  MXI2X1 U1825 ( .A(n969), .B(n970), .S0(n1162), .Y(blockdata[35]) );
  MXI4X1 U1826 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n1110), .S1(n1141), .Y(n969) );
  MXI4X1 U1827 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n1110), .S1(n1141), .Y(n970) );
  MXI2X1 U1828 ( .A(n967), .B(n968), .S0(n1160), .Y(blockdata[36]) );
  MXI4X1 U1829 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n1110), .S1(n1141), .Y(n967) );
  MXI4X1 U1830 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n1110), .S1(n1141), .Y(n968) );
  MXI2X1 U1831 ( .A(n965), .B(n966), .S0(n1159), .Y(blockdata[37]) );
  MXI4X1 U1832 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n1111), .S1(n1141), .Y(n965) );
  MXI4X1 U1833 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n1111), .S1(n1141), .Y(n966) );
  MXI2X1 U1834 ( .A(n963), .B(n964), .S0(n1162), .Y(blockdata[38]) );
  MXI4X1 U1835 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n1111), .S1(n1142), .Y(n963) );
  MXI4X1 U1836 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n1111), .S1(n1142), .Y(n964) );
  MXI2X1 U1837 ( .A(n961), .B(n962), .S0(n1164), .Y(blockdata[39]) );
  MXI4X1 U1838 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n1111), .S1(n1142), .Y(n961) );
  MXI4X1 U1839 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n1111), .S1(n1142), .Y(n962) );
  MXI2X1 U1840 ( .A(n959), .B(n960), .S0(n1162), .Y(blockdata[40]) );
  MXI4X1 U1841 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n1111), .S1(n1142), .Y(n959) );
  MXI4X1 U1842 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n1111), .S1(n1142), .Y(n960) );
  MXI2X1 U1843 ( .A(n957), .B(n958), .S0(n1164), .Y(blockdata[41]) );
  MXI4X1 U1844 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n1111), .S1(n1142), .Y(n957) );
  MXI4X1 U1845 ( .A(\block[4][41] ), .B(\block[5][41] ), .C(\block[6][41] ), 
        .D(\block[7][41] ), .S0(n1111), .S1(n1142), .Y(n958) );
  MXI2X1 U1846 ( .A(n955), .B(n956), .S0(n1159), .Y(blockdata[42]) );
  MXI4X1 U1847 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n1111), .S1(n1142), .Y(n955) );
  MXI4X1 U1848 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n1111), .S1(n1142), .Y(n956) );
  MXI2X1 U1849 ( .A(n953), .B(n954), .S0(n1164), .Y(blockdata[43]) );
  MXI4X1 U1850 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n1111), .S1(n1142), .Y(n953) );
  MXI4X1 U1851 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n1112), .S1(n1142), .Y(n954) );
  MXI2X1 U1852 ( .A(n951), .B(n952), .S0(n1161), .Y(blockdata[44]) );
  MXI4X1 U1853 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n1112), .S1(n1143), .Y(n951) );
  MXI4X1 U1854 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n1112), .S1(n1143), .Y(n952) );
  MXI2X1 U1855 ( .A(n949), .B(n950), .S0(n1160), .Y(blockdata[45]) );
  MXI4X1 U1856 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n1112), .S1(n1143), .Y(n949) );
  MXI4X1 U1857 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n1112), .S1(n1143), .Y(n950) );
  MXI2X1 U1858 ( .A(n947), .B(n948), .S0(n1162), .Y(blockdata[46]) );
  MXI4X1 U1859 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n1112), .S1(n1143), .Y(n947) );
  MXI4X1 U1860 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n1112), .S1(n1143), .Y(n948) );
  MXI2X1 U1861 ( .A(n945), .B(n946), .S0(n1161), .Y(blockdata[47]) );
  MXI4X1 U1862 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n1112), .S1(n1143), .Y(n945) );
  MXI4X1 U1863 ( .A(\block[4][47] ), .B(\block[5][47] ), .C(\block[6][47] ), 
        .D(\block[7][47] ), .S0(n1112), .S1(n1143), .Y(n946) );
  MXI2X1 U1864 ( .A(n943), .B(n944), .S0(n1164), .Y(blockdata[48]) );
  MXI4X1 U1865 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n1112), .S1(n1143), .Y(n943) );
  MXI4X1 U1866 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n1112), .S1(n1143), .Y(n944) );
  MXI2X1 U1867 ( .A(n941), .B(n942), .S0(n1159), .Y(blockdata[49]) );
  MXI4X1 U1868 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n1112), .S1(n1143), .Y(n941) );
  MXI4X1 U1869 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n1112), .S1(n1143), .Y(n942) );
  MXI2X1 U1870 ( .A(n939), .B(n940), .S0(n1160), .Y(blockdata[50]) );
  MXI4X1 U1871 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n1113), .S1(n1144), .Y(n939) );
  MXI4X1 U1872 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n1113), .S1(n1144), .Y(n940) );
  MXI2X1 U1873 ( .A(n937), .B(n938), .S0(n1162), .Y(blockdata[51]) );
  MXI4X1 U1874 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n1113), .S1(n1144), .Y(n937) );
  MXI4X1 U1875 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n1113), .S1(n1144), .Y(n938) );
  MXI2X1 U1876 ( .A(n935), .B(n936), .S0(n1159), .Y(blockdata[52]) );
  MXI4X1 U1877 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n1113), .S1(n1144), .Y(n935) );
  MXI4X1 U1878 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n1113), .S1(n1144), .Y(n936) );
  MXI2X1 U1879 ( .A(n933), .B(n934), .S0(n1160), .Y(blockdata[53]) );
  MXI4X1 U1880 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n1113), .S1(n1144), .Y(n933) );
  MXI4X1 U1881 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n1113), .S1(n1144), .Y(n934) );
  MXI2X1 U1882 ( .A(n931), .B(n932), .S0(n1162), .Y(blockdata[54]) );
  MXI4X1 U1883 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n1113), .S1(n1144), .Y(n931) );
  MXI4X1 U1884 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n1113), .S1(n1144), .Y(n932) );
  MXI2X1 U1885 ( .A(n929), .B(n930), .S0(n1159), .Y(blockdata[55]) );
  MXI4X1 U1886 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n1113), .S1(n1144), .Y(n929) );
  MXI4X1 U1887 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n1113), .S1(n1144), .Y(n930) );
  MXI2X1 U1888 ( .A(n927), .B(n928), .S0(n1161), .Y(blockdata[56]) );
  MXI4X1 U1889 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n1113), .S1(n1145), .Y(n927) );
  MXI4X1 U1890 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n1114), .S1(n1145), .Y(n928) );
  MXI2X1 U1891 ( .A(n925), .B(n926), .S0(n1160), .Y(blockdata[57]) );
  MXI4X1 U1892 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n1114), .S1(n1145), .Y(n925) );
  MXI4X1 U1893 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n1114), .S1(n1145), .Y(n926) );
  MXI2X1 U1894 ( .A(n923), .B(n924), .S0(n1166), .Y(blockdata[58]) );
  MXI4X1 U1895 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n1114), .S1(n1145), .Y(n923) );
  MXI4X1 U1896 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n1114), .S1(n1145), .Y(n924) );
  MXI2X1 U1897 ( .A(n921), .B(n922), .S0(n1162), .Y(blockdata[59]) );
  MXI4X1 U1898 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n1114), .S1(n1145), .Y(n921) );
  MXI4X1 U1899 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n1114), .S1(n1145), .Y(n922) );
  MXI2X1 U1900 ( .A(n919), .B(n920), .S0(n1163), .Y(blockdata[60]) );
  MXI4X1 U1901 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n1114), .S1(n1145), .Y(n919) );
  MXI4X1 U1902 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n1114), .S1(n1145), .Y(n920) );
  MXI2X1 U1903 ( .A(n917), .B(n918), .S0(n1162), .Y(blockdata[61]) );
  MXI4X1 U1904 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n1114), .S1(n1145), .Y(n917) );
  MXI4X1 U1905 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n1114), .S1(n1145), .Y(n918) );
  MXI2X1 U1906 ( .A(n915), .B(n916), .S0(n1166), .Y(blockdata[62]) );
  MXI4X1 U1907 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n1114), .S1(n1146), .Y(n915) );
  MXI4X1 U1908 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n1114), .S1(n1146), .Y(n916) );
  MXI2X1 U1909 ( .A(n913), .B(n914), .S0(n1161), .Y(blockdata[63]) );
  MXI4X1 U1910 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n1113), .S1(n1146), .Y(n913) );
  MXI4X1 U1911 ( .A(\block[4][63] ), .B(\block[5][63] ), .C(\block[6][63] ), 
        .D(\block[7][63] ), .S0(n1112), .S1(n1146), .Y(n914) );
  MXI2X1 U1912 ( .A(n911), .B(n912), .S0(n1165), .Y(blockdata[64]) );
  MXI4X1 U1913 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n1111), .S1(n1146), .Y(n911) );
  MXI4X1 U1914 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n1115), .S1(n1146), .Y(n912) );
  MXI2X1 U1915 ( .A(n909), .B(n910), .S0(n1165), .Y(blockdata[65]) );
  MXI4X1 U1916 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n1114), .S1(n1146), .Y(n909) );
  MXI4X1 U1917 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n1111), .S1(n1146), .Y(n910) );
  MXI2X1 U1918 ( .A(n907), .B(n908), .S0(n1165), .Y(blockdata[66]) );
  MXI4X1 U1919 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n1123), .S1(n1146), .Y(n907) );
  MXI4X1 U1920 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n1114), .S1(n1146), .Y(n908) );
  MXI2X1 U1921 ( .A(n905), .B(n906), .S0(n1167), .Y(blockdata[67]) );
  MXI4X1 U1922 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n1118), .S1(n1146), .Y(n905) );
  MXI4X1 U1923 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n1123), .S1(n1146), .Y(n906) );
  MXI2X1 U1924 ( .A(n903), .B(n904), .S0(n1160), .Y(blockdata[68]) );
  MXI4X1 U1925 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n1119), .S1(n1147), .Y(n903) );
  MXI4X1 U1926 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n1122), .S1(n1147), .Y(n904) );
  MXI2X1 U1927 ( .A(n901), .B(n902), .S0(n1162), .Y(blockdata[69]) );
  MXI4X1 U1928 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n1122), .S1(n1147), .Y(n901) );
  MXI4X1 U1929 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n1115), .S1(n1147), .Y(n902) );
  MXI2X1 U1930 ( .A(n899), .B(n900), .S0(n1159), .Y(blockdata[70]) );
  MXI4X1 U1931 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n1115), .S1(n1147), .Y(n899) );
  MXI4X1 U1932 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n1115), .S1(n1147), .Y(n900) );
  MXI2X1 U1933 ( .A(n897), .B(n898), .S0(n1160), .Y(blockdata[71]) );
  MXI4X1 U1934 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n1115), .S1(n1147), .Y(n897) );
  MXI4X1 U1935 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n1115), .S1(n1147), .Y(n898) );
  MXI2X1 U1936 ( .A(n895), .B(n896), .S0(n1162), .Y(blockdata[72]) );
  MXI4X1 U1937 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n1115), .S1(n1147), .Y(n895) );
  MXI4X1 U1938 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n1115), .S1(n1147), .Y(n896) );
  MXI2X1 U1939 ( .A(n893), .B(n894), .S0(n1159), .Y(blockdata[73]) );
  MXI4X1 U1940 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n1115), .S1(n1147), .Y(n893) );
  MXI4X1 U1941 ( .A(\block[4][73] ), .B(\block[5][73] ), .C(\block[6][73] ), 
        .D(\block[7][73] ), .S0(n1115), .S1(n1147), .Y(n894) );
  MXI2X1 U1942 ( .A(n891), .B(n892), .S0(n1160), .Y(blockdata[74]) );
  MXI4X1 U1943 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n1115), .S1(n1148), .Y(n891) );
  MXI4X1 U1944 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n1115), .S1(n1148), .Y(n892) );
  MXI2X1 U1945 ( .A(n889), .B(n890), .S0(n1162), .Y(blockdata[75]) );
  MXI4X1 U1946 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n1115), .S1(n1148), .Y(n889) );
  MXI4X1 U1947 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n1115), .S1(n1148), .Y(n890) );
  MXI2X1 U1948 ( .A(n887), .B(n888), .S0(n1159), .Y(blockdata[76]) );
  MXI4X1 U1949 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n1116), .S1(n1148), .Y(n887) );
  MXI4X1 U1950 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n1116), .S1(n1148), .Y(n888) );
  MXI2X1 U1951 ( .A(n885), .B(n886), .S0(n1160), .Y(blockdata[77]) );
  MXI4X1 U1952 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n1116), .S1(n1148), .Y(n885) );
  MXI4X1 U1953 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n1116), .S1(n1148), .Y(n886) );
  MXI2X1 U1954 ( .A(n883), .B(n884), .S0(n1162), .Y(blockdata[78]) );
  MXI4X1 U1955 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n1116), .S1(n1148), .Y(n883) );
  MXI4X1 U1956 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n1116), .S1(n1148), .Y(n884) );
  MXI2X1 U1957 ( .A(n881), .B(n882), .S0(n1159), .Y(blockdata[79]) );
  MXI4X1 U1958 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n1116), .S1(n1148), .Y(n881) );
  MXI4X1 U1959 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n1116), .S1(n1148), .Y(n882) );
  MXI2X1 U1960 ( .A(n879), .B(n880), .S0(n1166), .Y(blockdata[80]) );
  MXI4X1 U1961 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n1116), .S1(n1149), .Y(n879) );
  MXI4X1 U1962 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n1116), .S1(n1149), .Y(n880) );
  MXI2X1 U1963 ( .A(n877), .B(n878), .S0(n1163), .Y(blockdata[81]) );
  MXI4X1 U1964 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n1116), .S1(n1149), .Y(n877) );
  MXI4X1 U1965 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n1116), .S1(n1149), .Y(n878) );
  MXI2X1 U1966 ( .A(n875), .B(n876), .S0(n1159), .Y(blockdata[82]) );
  MXI4X1 U1967 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n1116), .S1(n1149), .Y(n875) );
  MXI4X1 U1968 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n1117), .S1(n1149), .Y(n876) );
  MXI2X1 U1969 ( .A(n873), .B(n874), .S0(n1166), .Y(blockdata[83]) );
  MXI4X1 U1970 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n1117), .S1(n1149), .Y(n873) );
  MXI4X1 U1971 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n1117), .S1(n1149), .Y(n874) );
  MXI2X1 U1972 ( .A(n871), .B(n872), .S0(n1161), .Y(blockdata[84]) );
  MXI4X1 U1973 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n1117), .S1(n1149), .Y(n871) );
  MXI4X1 U1974 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n1117), .S1(n1149), .Y(n872) );
  MXI2X1 U1975 ( .A(n869), .B(n870), .S0(n1159), .Y(blockdata[85]) );
  MXI4X1 U1976 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n1117), .S1(n1149), .Y(n869) );
  MXI4X1 U1977 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n1117), .S1(n1149), .Y(n870) );
  MXI2X1 U1978 ( .A(n867), .B(n868), .S0(n1160), .Y(blockdata[86]) );
  MXI4X1 U1979 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n1117), .S1(n1150), .Y(n867) );
  MXI4X1 U1980 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n1117), .S1(n1150), .Y(n868) );
  MXI2X1 U1981 ( .A(n865), .B(n866), .S0(n1163), .Y(blockdata[87]) );
  MXI4X1 U1982 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n1117), .S1(n1150), .Y(n865) );
  MXI4X1 U1983 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n1117), .S1(n1150), .Y(n866) );
  MXI2X1 U1984 ( .A(n863), .B(n864), .S0(n1166), .Y(blockdata[88]) );
  MXI4X1 U1985 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n1117), .S1(n1150), .Y(n863) );
  MXI4X1 U1986 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n1117), .S1(n1150), .Y(n864) );
  MXI2X1 U1987 ( .A(n861), .B(n862), .S0(n1158), .Y(blockdata[89]) );
  MXI4X1 U1988 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n1118), .S1(n1150), .Y(n861) );
  MXI4X1 U1989 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n1118), .S1(n1150), .Y(n862) );
  MXI2X1 U1990 ( .A(n859), .B(n860), .S0(n1159), .Y(blockdata[90]) );
  MXI4X1 U1991 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n1118), .S1(n1150), .Y(n859) );
  MXI4X1 U1992 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n1118), .S1(n1150), .Y(n860) );
  MXI2X1 U1993 ( .A(n857), .B(n858), .S0(n1162), .Y(blockdata[91]) );
  MXI4X1 U1994 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n1118), .S1(n1150), .Y(n857) );
  MXI4X1 U1995 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n1118), .S1(n1150), .Y(n858) );
  MXI2X1 U1996 ( .A(n855), .B(n856), .S0(n1167), .Y(blockdata[92]) );
  MXI4X1 U1997 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n1118), .S1(n1151), .Y(n855) );
  MXI4X1 U1998 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n1118), .S1(n1151), .Y(n856) );
  MXI2X1 U1999 ( .A(n853), .B(n854), .S0(n1167), .Y(blockdata[93]) );
  MXI4X1 U2000 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n1118), .S1(n1151), .Y(n853) );
  MXI4X1 U2001 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n1118), .S1(n1151), .Y(n854) );
  MXI2X1 U2002 ( .A(n851), .B(n852), .S0(n1167), .Y(blockdata[94]) );
  MXI4X1 U2003 ( .A(\block[0][94] ), .B(\block[1][94] ), .C(\block[2][94] ), 
        .D(\block[3][94] ), .S0(n1118), .S1(n1151), .Y(n851) );
  MXI4X1 U2004 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), 
        .D(\block[7][94] ), .S0(n1118), .S1(n1151), .Y(n852) );
  MXI2X1 U2005 ( .A(n849), .B(n850), .S0(n1167), .Y(blockdata[95]) );
  MXI4X1 U2006 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n1118), .S1(n1151), .Y(n849) );
  MXI4X1 U2007 ( .A(\block[4][95] ), .B(\block[5][95] ), .C(\block[6][95] ), 
        .D(\block[7][95] ), .S0(n1119), .S1(n1151), .Y(n850) );
  MXI2X1 U2008 ( .A(n847), .B(n848), .S0(n1167), .Y(blockdata[96]) );
  MXI4X1 U2009 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n1119), .S1(n1151), .Y(n847) );
  MXI4X1 U2010 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n1119), .S1(n1151), .Y(n848) );
  MXI2X1 U2011 ( .A(n845), .B(n846), .S0(n1167), .Y(blockdata[97]) );
  MXI4X1 U2012 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n1119), .S1(n1151), .Y(n845) );
  MXI4X1 U2013 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n1119), .S1(n1151), .Y(n846) );
  MXI2X1 U2014 ( .A(n843), .B(n844), .S0(n1167), .Y(blockdata[98]) );
  MXI4X1 U2015 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n1119), .S1(n1152), .Y(n843) );
  MXI4X1 U2016 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n1119), .S1(n1152), .Y(n844) );
  MXI2X1 U2017 ( .A(n841), .B(n842), .S0(n1167), .Y(blockdata[99]) );
  MXI4X1 U2018 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n1119), .S1(n1152), .Y(n841) );
  MXI4X1 U2019 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n1119), .S1(n1152), .Y(n842) );
  MXI2X1 U2020 ( .A(n839), .B(n840), .S0(n1167), .Y(blockdata[100]) );
  MXI4X1 U2021 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n1119), .S1(n1152), .Y(n839) );
  MXI4X1 U2022 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n1119), .S1(n1152), .Y(n840) );
  MXI2X1 U2023 ( .A(n837), .B(n838), .S0(n1167), .Y(blockdata[101]) );
  MXI4X1 U2024 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n1119), .S1(n1152), .Y(n837) );
  MXI4X1 U2025 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n1119), .S1(n1152), .Y(n838) );
  MXI2X1 U2026 ( .A(n835), .B(n836), .S0(n1167), .Y(blockdata[102]) );
  MXI4X1 U2027 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n1120), .S1(n1152), .Y(n835) );
  MXI4X1 U2028 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n1120), .S1(n1152), .Y(n836) );
  MXI2X1 U2029 ( .A(n833), .B(n834), .S0(n1167), .Y(blockdata[103]) );
  MXI4X1 U2030 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n1120), .S1(n1152), .Y(n833) );
  MXI4X1 U2031 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n1120), .S1(n1152), .Y(n834) );
  MXI2X1 U2032 ( .A(n831), .B(n832), .S0(n1168), .Y(blockdata[104]) );
  MXI4X1 U2033 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n1120), .S1(n1153), .Y(n831) );
  MXI4X1 U2034 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n1120), .S1(n1153), .Y(n832) );
  MXI2X1 U2035 ( .A(n829), .B(n830), .S0(n1168), .Y(blockdata[105]) );
  MXI4X1 U2036 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n1120), .S1(n1153), .Y(n829) );
  MXI4X1 U2037 ( .A(\block[4][105] ), .B(\block[5][105] ), .C(\block[6][105] ), 
        .D(\block[7][105] ), .S0(n1120), .S1(n1153), .Y(n830) );
  MXI2X1 U2038 ( .A(n827), .B(n828), .S0(n1168), .Y(blockdata[106]) );
  MXI4X1 U2039 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n1120), .S1(n1153), .Y(n827) );
  MXI4X1 U2040 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n1120), .S1(n1153), .Y(n828) );
  MXI2X1 U2041 ( .A(n825), .B(n826), .S0(n1168), .Y(blockdata[107]) );
  MXI4X1 U2042 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n1120), .S1(n1153), .Y(n825) );
  MXI4X1 U2043 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n1120), .S1(n1153), .Y(n826) );
  MXI2X1 U2044 ( .A(n823), .B(n824), .S0(n1168), .Y(blockdata[108]) );
  MXI4X1 U2045 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n1120), .S1(n1153), .Y(n823) );
  MXI4X1 U2046 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n1121), .S1(n1153), .Y(n824) );
  MXI2X1 U2047 ( .A(n821), .B(n822), .S0(n1168), .Y(blockdata[109]) );
  MXI4X1 U2048 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n1121), .S1(n1153), .Y(n821) );
  MXI4X1 U2049 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n1121), .S1(n1153), .Y(n822) );
  MXI2X1 U2050 ( .A(n819), .B(n820), .S0(n1168), .Y(blockdata[110]) );
  MXI4X1 U2051 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n1121), .S1(n1154), .Y(n819) );
  MXI4X1 U2052 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n1121), .S1(n1154), .Y(n820) );
  MXI2X1 U2053 ( .A(n817), .B(n818), .S0(n1168), .Y(blockdata[111]) );
  MXI4X1 U2054 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n1121), .S1(n1154), .Y(n817) );
  MXI4X1 U2055 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n1121), .S1(n1154), .Y(n818) );
  MXI2X1 U2056 ( .A(n815), .B(n816), .S0(n1168), .Y(blockdata[112]) );
  MXI4X1 U2057 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n1121), .S1(n1154), .Y(n815) );
  MXI4X1 U2058 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n1121), .S1(n1154), .Y(n816) );
  MXI2X1 U2059 ( .A(n813), .B(n814), .S0(n1168), .Y(blockdata[113]) );
  MXI4X1 U2060 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n1121), .S1(n1154), .Y(n813) );
  MXI4X1 U2061 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n1121), .S1(n1154), .Y(n814) );
  MXI2X1 U2062 ( .A(n811), .B(n812), .S0(n1168), .Y(blockdata[114]) );
  MXI4X1 U2063 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n1121), .S1(n1154), .Y(n811) );
  MXI4X1 U2064 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n1121), .S1(n1154), .Y(n812) );
  MXI2X1 U2065 ( .A(n809), .B(n810), .S0(n1168), .Y(blockdata[115]) );
  MXI4X1 U2066 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n1122), .S1(n1154), .Y(n809) );
  MXI4X1 U2067 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n1122), .S1(n1154), .Y(n810) );
  MXI2X1 U2068 ( .A(n807), .B(n808), .S0(n1168), .Y(blockdata[116]) );
  MXI4X1 U2069 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n1122), .S1(n1155), .Y(n807) );
  MXI4X1 U2070 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n1122), .S1(n1155), .Y(n808) );
  MXI2X1 U2071 ( .A(n805), .B(n806), .S0(n1168), .Y(blockdata[117]) );
  MXI4X1 U2072 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n1122), .S1(n1155), .Y(n805) );
  MXI4X1 U2073 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n1122), .S1(n1155), .Y(n806) );
  MXI2X1 U2074 ( .A(n803), .B(n804), .S0(n1167), .Y(blockdata[118]) );
  MXI4X1 U2075 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n1122), .S1(n1155), .Y(n803) );
  MXI4X1 U2076 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n1122), .S1(n1155), .Y(n804) );
  MXI2X1 U2077 ( .A(n801), .B(n802), .S0(n1165), .Y(blockdata[119]) );
  MXI4X1 U2078 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n1122), .S1(n1155), .Y(n801) );
  MXI4X1 U2079 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n1122), .S1(n1155), .Y(n802) );
  MXI2X1 U2080 ( .A(n799), .B(n800), .S0(n1168), .Y(blockdata[120]) );
  MXI4X1 U2081 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n1122), .S1(n1155), .Y(n799) );
  MXI4X1 U2082 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n1122), .S1(n1155), .Y(n800) );
  MXI2X1 U2083 ( .A(n797), .B(n798), .S0(n1167), .Y(blockdata[121]) );
  MXI4X1 U2084 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n1122), .S1(n1155), .Y(n797) );
  MXI4X1 U2085 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n1123), .S1(n1155), .Y(n798) );
  MXI2X1 U2086 ( .A(n795), .B(n796), .S0(n1168), .Y(blockdata[122]) );
  MXI4X1 U2087 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n1123), .S1(n1156), .Y(n795) );
  MXI4X1 U2088 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n1123), .S1(n1156), .Y(n796) );
  MXI2X1 U2089 ( .A(n793), .B(n794), .S0(n1167), .Y(blockdata[123]) );
  MXI4X1 U2090 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n1123), .S1(n1156), .Y(n793) );
  MXI4X1 U2091 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n1123), .S1(n1156), .Y(n794) );
  MXI2X1 U2092 ( .A(n791), .B(n792), .S0(n1168), .Y(blockdata[124]) );
  MXI4X1 U2093 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n1123), .S1(n1156), .Y(n791) );
  MXI4X1 U2094 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n1123), .S1(n1156), .Y(n792) );
  MXI2X1 U2095 ( .A(n789), .B(n790), .S0(n1167), .Y(blockdata[125]) );
  MXI4X1 U2096 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n1123), .S1(n1156), .Y(n789) );
  MXI4X1 U2097 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n1123), .S1(n1156), .Y(n790) );
  MXI2X1 U2098 ( .A(n787), .B(n788), .S0(n1163), .Y(blockdata[126]) );
  MXI4X1 U2099 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n1123), .S1(n1156), .Y(n787) );
  MXI4X1 U2100 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n1123), .S1(n1156), .Y(n788) );
  MXI2X1 U2101 ( .A(n785), .B(n786), .S0(n1163), .Y(blockdata[127]) );
  MXI4X1 U2102 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n1123), .S1(n1156), .Y(n785) );
  MXI4X1 U2103 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n1123), .S1(n1156), .Y(n786) );
  OAI22XL U2104 ( .A0(n589), .A1(n1464), .B0(n17), .B1(n18), .Y(n608) );
  OAI22XL U2105 ( .A0(n590), .A1(n1463), .B0(n17), .B1(n20), .Y(n609) );
  OAI22XL U2106 ( .A0(n591), .A1(n1466), .B0(n17), .B1(n22), .Y(n610) );
  OAI22XL U2107 ( .A0(n592), .A1(n1465), .B0(n17), .B1(n24), .Y(n611) );
  OAI22XL U2108 ( .A0(n593), .A1(n1469), .B0(n17), .B1(n26), .Y(n612) );
  OAI22XL U2109 ( .A0(n594), .A1(n1468), .B0(n17), .B1(n28), .Y(n613) );
  OAI22XL U2110 ( .A0(n595), .A1(n1471), .B0(n17), .B1(n30), .Y(n614) );
  OAI22XL U2111 ( .A0(n597), .A1(n1470), .B0(n17), .B1(n32), .Y(n615) );
  OAI22XL U2112 ( .A0(n598), .A1(n1464), .B0(n35), .B1(n18), .Y(n616) );
  OAI22XL U2113 ( .A0(n599), .A1(n1463), .B0(n35), .B1(n20), .Y(n617) );
  OAI22XL U2114 ( .A0(n600), .A1(n1466), .B0(n35), .B1(n22), .Y(n618) );
  OAI22XL U2115 ( .A0(n601), .A1(n1465), .B0(n35), .B1(n24), .Y(n619) );
  OAI22XL U2116 ( .A0(n602), .A1(n1469), .B0(n35), .B1(n26), .Y(n620) );
  OAI22XL U2117 ( .A0(n603), .A1(n1468), .B0(n35), .B1(n28), .Y(n621) );
  OAI22XL U2118 ( .A0(n604), .A1(n1471), .B0(n35), .B1(n30), .Y(n622) );
  OAI22XL U2119 ( .A0(n605), .A1(n1470), .B0(n35), .B1(n32), .Y(n623) );
  NOR2X1 U2120 ( .A(state[1]), .B(state[2]), .Y(n503) );
  CLKINVX1 U2121 ( .A(mem_ready_r), .Y(n1508) );
  CLKINVX1 U2122 ( .A(wordIndex[0]), .Y(n1475) );
  CLKINVX1 U2123 ( .A(wordIndex[1]), .Y(n1474) );
  CLKINVX1 U2124 ( .A(mem_rdata_r[64]), .Y(n1575) );
  CLKINVX1 U2125 ( .A(mem_rdata_r[65]), .Y(n1574) );
  CLKINVX1 U2126 ( .A(mem_rdata_r[66]), .Y(n1573) );
  CLKINVX1 U2127 ( .A(mem_rdata_r[67]), .Y(n1572) );
  CLKINVX1 U2128 ( .A(mem_rdata_r[68]), .Y(n1571) );
  CLKINVX1 U2129 ( .A(mem_rdata_r[69]), .Y(n1570) );
  CLKINVX1 U2130 ( .A(mem_rdata_r[70]), .Y(n1569) );
  CLKINVX1 U2131 ( .A(mem_rdata_r[71]), .Y(n1568) );
  CLKINVX1 U2132 ( .A(mem_rdata_r[72]), .Y(n1567) );
  CLKINVX1 U2133 ( .A(mem_rdata_r[73]), .Y(n1566) );
  CLKINVX1 U2134 ( .A(mem_rdata_r[74]), .Y(n1565) );
  CLKINVX1 U2135 ( .A(mem_rdata_r[75]), .Y(n1564) );
  CLKINVX1 U2136 ( .A(mem_rdata_r[76]), .Y(n1563) );
  CLKINVX1 U2137 ( .A(mem_rdata_r[77]), .Y(n1562) );
  CLKINVX1 U2138 ( .A(mem_rdata_r[78]), .Y(n1561) );
  CLKINVX1 U2139 ( .A(mem_rdata_r[79]), .Y(n1560) );
  CLKINVX1 U2140 ( .A(mem_rdata_r[80]), .Y(n1559) );
  CLKINVX1 U2141 ( .A(mem_rdata_r[81]), .Y(n1558) );
  CLKINVX1 U2142 ( .A(mem_rdata_r[82]), .Y(n1557) );
  CLKINVX1 U2143 ( .A(mem_rdata_r[83]), .Y(n1556) );
  CLKINVX1 U2144 ( .A(mem_rdata_r[84]), .Y(n1555) );
  CLKINVX1 U2145 ( .A(mem_rdata_r[85]), .Y(n1554) );
  CLKINVX1 U2146 ( .A(mem_rdata_r[86]), .Y(n1553) );
  CLKINVX1 U2147 ( .A(mem_rdata_r[87]), .Y(n1552) );
  CLKINVX1 U2148 ( .A(mem_rdata_r[88]), .Y(n1551) );
  CLKINVX1 U2149 ( .A(mem_rdata_r[89]), .Y(n1550) );
  CLKINVX1 U2150 ( .A(mem_rdata_r[90]), .Y(n1549) );
  CLKINVX1 U2151 ( .A(mem_rdata_r[91]), .Y(n1548) );
  CLKINVX1 U2152 ( .A(mem_rdata_r[92]), .Y(n1547) );
  CLKINVX1 U2153 ( .A(mem_rdata_r[93]), .Y(n1546) );
  CLKINVX1 U2154 ( .A(mem_rdata_r[94]), .Y(n1545) );
  CLKINVX1 U2155 ( .A(mem_rdata_r[95]), .Y(n1544) );
  CLKINVX1 U2156 ( .A(mem_rdata_r[96]), .Y(n1543) );
  CLKINVX1 U2157 ( .A(mem_rdata_r[97]), .Y(n1542) );
  CLKINVX1 U2158 ( .A(mem_rdata_r[98]), .Y(n1541) );
  CLKINVX1 U2159 ( .A(mem_rdata_r[99]), .Y(n1540) );
  CLKINVX1 U2160 ( .A(mem_rdata_r[100]), .Y(n1539) );
  CLKINVX1 U2161 ( .A(mem_rdata_r[101]), .Y(n1538) );
  CLKINVX1 U2162 ( .A(mem_rdata_r[102]), .Y(n1537) );
  CLKINVX1 U2163 ( .A(mem_rdata_r[103]), .Y(n1536) );
  CLKINVX1 U2164 ( .A(mem_rdata_r[104]), .Y(n1535) );
  CLKINVX1 U2165 ( .A(mem_rdata_r[105]), .Y(n1534) );
  CLKINVX1 U2166 ( .A(mem_rdata_r[106]), .Y(n1533) );
  CLKINVX1 U2167 ( .A(mem_rdata_r[107]), .Y(n1532) );
  CLKINVX1 U2168 ( .A(mem_rdata_r[108]), .Y(n1531) );
  CLKINVX1 U2169 ( .A(mem_rdata_r[109]), .Y(n1530) );
  CLKINVX1 U2170 ( .A(mem_rdata_r[110]), .Y(n1529) );
  CLKINVX1 U2171 ( .A(mem_rdata_r[111]), .Y(n1528) );
  CLKINVX1 U2172 ( .A(mem_rdata_r[112]), .Y(n1527) );
  CLKINVX1 U2173 ( .A(mem_rdata_r[113]), .Y(n1526) );
  CLKINVX1 U2174 ( .A(mem_rdata_r[114]), .Y(n1525) );
  CLKINVX1 U2175 ( .A(mem_rdata_r[115]), .Y(n1524) );
  CLKINVX1 U2176 ( .A(mem_rdata_r[116]), .Y(n1523) );
  CLKINVX1 U2177 ( .A(mem_rdata_r[117]), .Y(n1522) );
  CLKINVX1 U2178 ( .A(mem_rdata_r[118]), .Y(n1521) );
  CLKINVX1 U2179 ( .A(mem_rdata_r[119]), .Y(n1520) );
  CLKINVX1 U2180 ( .A(mem_rdata_r[120]), .Y(n1519) );
  CLKINVX1 U2181 ( .A(mem_rdata_r[121]), .Y(n1518) );
  CLKINVX1 U2182 ( .A(mem_rdata_r[122]), .Y(n1517) );
  CLKINVX1 U2183 ( .A(mem_rdata_r[123]), .Y(n1516) );
  CLKINVX1 U2184 ( .A(mem_rdata_r[124]), .Y(n1515) );
  CLKINVX1 U2185 ( .A(mem_rdata_r[125]), .Y(n1514) );
  CLKINVX1 U2186 ( .A(mem_rdata_r[126]), .Y(n1513) );
  CLKINVX1 U2187 ( .A(mem_rdata_r[127]), .Y(n1512) );
  CLKINVX1 U2188 ( .A(mem_rdata_r[0]), .Y(n1639) );
  CLKINVX1 U2189 ( .A(mem_rdata_r[1]), .Y(n1638) );
  CLKINVX1 U2190 ( .A(mem_rdata_r[2]), .Y(n1637) );
  CLKINVX1 U2191 ( .A(mem_rdata_r[3]), .Y(n1636) );
  CLKINVX1 U2192 ( .A(mem_rdata_r[4]), .Y(n1635) );
  CLKINVX1 U2193 ( .A(mem_rdata_r[5]), .Y(n1634) );
  CLKINVX1 U2194 ( .A(mem_rdata_r[6]), .Y(n1633) );
  CLKINVX1 U2195 ( .A(mem_rdata_r[7]), .Y(n1632) );
  CLKINVX1 U2196 ( .A(mem_rdata_r[8]), .Y(n1631) );
  CLKINVX1 U2197 ( .A(mem_rdata_r[9]), .Y(n1630) );
  CLKINVX1 U2198 ( .A(mem_rdata_r[10]), .Y(n1629) );
  CLKINVX1 U2199 ( .A(mem_rdata_r[11]), .Y(n1628) );
  CLKINVX1 U2200 ( .A(mem_rdata_r[12]), .Y(n1627) );
  CLKINVX1 U2201 ( .A(mem_rdata_r[13]), .Y(n1626) );
  CLKINVX1 U2202 ( .A(mem_rdata_r[14]), .Y(n1625) );
  CLKINVX1 U2203 ( .A(mem_rdata_r[15]), .Y(n1624) );
  CLKINVX1 U2204 ( .A(mem_rdata_r[16]), .Y(n1623) );
  CLKINVX1 U2205 ( .A(mem_rdata_r[17]), .Y(n1622) );
  CLKINVX1 U2206 ( .A(mem_rdata_r[18]), .Y(n1621) );
  CLKINVX1 U2207 ( .A(mem_rdata_r[19]), .Y(n1620) );
  CLKINVX1 U2208 ( .A(mem_rdata_r[20]), .Y(n1619) );
  CLKINVX1 U2209 ( .A(mem_rdata_r[21]), .Y(n1618) );
  CLKINVX1 U2210 ( .A(mem_rdata_r[22]), .Y(n1617) );
  CLKINVX1 U2211 ( .A(mem_rdata_r[23]), .Y(n1616) );
  CLKINVX1 U2212 ( .A(mem_rdata_r[24]), .Y(n1615) );
  CLKINVX1 U2213 ( .A(mem_rdata_r[25]), .Y(n1614) );
  CLKINVX1 U2214 ( .A(mem_rdata_r[26]), .Y(n1613) );
  CLKINVX1 U2215 ( .A(mem_rdata_r[27]), .Y(n1612) );
  CLKINVX1 U2216 ( .A(mem_rdata_r[28]), .Y(n1611) );
  CLKINVX1 U2217 ( .A(mem_rdata_r[29]), .Y(n1610) );
  CLKINVX1 U2218 ( .A(mem_rdata_r[30]), .Y(n1609) );
  CLKINVX1 U2219 ( .A(mem_rdata_r[31]), .Y(n1608) );
  CLKINVX1 U2220 ( .A(mem_rdata_r[32]), .Y(n1607) );
  CLKINVX1 U2221 ( .A(mem_rdata_r[33]), .Y(n1606) );
  CLKINVX1 U2222 ( .A(mem_rdata_r[34]), .Y(n1605) );
  CLKINVX1 U2223 ( .A(mem_rdata_r[35]), .Y(n1604) );
  CLKINVX1 U2224 ( .A(mem_rdata_r[36]), .Y(n1603) );
  CLKINVX1 U2225 ( .A(mem_rdata_r[37]), .Y(n1602) );
  CLKINVX1 U2226 ( .A(mem_rdata_r[38]), .Y(n1601) );
  CLKINVX1 U2227 ( .A(mem_rdata_r[39]), .Y(n1600) );
  CLKINVX1 U2228 ( .A(mem_rdata_r[40]), .Y(n1599) );
  CLKINVX1 U2229 ( .A(mem_rdata_r[41]), .Y(n1598) );
  CLKINVX1 U2230 ( .A(mem_rdata_r[42]), .Y(n1597) );
  CLKINVX1 U2231 ( .A(mem_rdata_r[43]), .Y(n1596) );
  CLKINVX1 U2232 ( .A(mem_rdata_r[44]), .Y(n1595) );
  CLKINVX1 U2233 ( .A(mem_rdata_r[45]), .Y(n1594) );
  CLKINVX1 U2234 ( .A(mem_rdata_r[46]), .Y(n1593) );
  CLKINVX1 U2235 ( .A(mem_rdata_r[47]), .Y(n1592) );
  CLKINVX1 U2236 ( .A(mem_rdata_r[48]), .Y(n1591) );
  CLKINVX1 U2237 ( .A(mem_rdata_r[49]), .Y(n1590) );
  CLKINVX1 U2238 ( .A(mem_rdata_r[50]), .Y(n1589) );
  CLKINVX1 U2239 ( .A(mem_rdata_r[51]), .Y(n1588) );
  CLKINVX1 U2240 ( .A(mem_rdata_r[52]), .Y(n1587) );
  CLKINVX1 U2241 ( .A(mem_rdata_r[53]), .Y(n1586) );
  CLKINVX1 U2242 ( .A(mem_rdata_r[54]), .Y(n1585) );
  CLKINVX1 U2243 ( .A(mem_rdata_r[55]), .Y(n1584) );
  CLKINVX1 U2244 ( .A(mem_rdata_r[56]), .Y(n1583) );
  CLKINVX1 U2245 ( .A(mem_rdata_r[57]), .Y(n1582) );
  CLKINVX1 U2246 ( .A(mem_rdata_r[58]), .Y(n1581) );
  CLKINVX1 U2247 ( .A(mem_rdata_r[59]), .Y(n1580) );
  CLKINVX1 U2248 ( .A(mem_rdata_r[60]), .Y(n1579) );
  CLKINVX1 U2249 ( .A(mem_rdata_r[61]), .Y(n1578) );
  CLKINVX1 U2250 ( .A(mem_rdata_r[62]), .Y(n1577) );
  CLKINVX1 U2251 ( .A(mem_rdata_r[63]), .Y(n1576) );
  INVX4 U2252 ( .A(n703), .Y(n1305) );
endmodule

