
module cache ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1419, \blocktag[7][24] , \blocktag[7][22] ,
         \blocktag[7][20] , \blocktag[7][18] , \blocktag[7][17] ,
         \blocktag[7][16] , \blocktag[7][15] , \blocktag[7][14] ,
         \blocktag[7][13] , \blocktag[7][12] , \blocktag[7][11] ,
         \blocktag[7][10] , \blocktag[7][9] , \blocktag[7][8] ,
         \blocktag[7][7] , \blocktag[7][6] , \blocktag[7][5] ,
         \blocktag[7][4] , \blocktag[7][3] , \blocktag[7][2] ,
         \blocktag[7][1] , \blocktag[6][24] , \blocktag[6][22] ,
         \blocktag[6][20] , \blocktag[6][18] , \blocktag[6][17] ,
         \blocktag[6][16] , \blocktag[6][15] , \blocktag[6][14] ,
         \blocktag[6][13] , \blocktag[6][12] , \blocktag[6][11] ,
         \blocktag[6][10] , \blocktag[6][9] , \blocktag[6][8] ,
         \blocktag[6][7] , \blocktag[6][6] , \blocktag[6][5] ,
         \blocktag[6][4] , \blocktag[6][3] , \blocktag[6][2] ,
         \blocktag[6][1] , \blocktag[5][24] , \blocktag[5][22] ,
         \blocktag[5][20] , \blocktag[5][18] , \blocktag[5][17] ,
         \blocktag[5][16] , \blocktag[5][15] , \blocktag[5][14] ,
         \blocktag[5][13] , \blocktag[5][12] , \blocktag[5][11] ,
         \blocktag[5][10] , \blocktag[5][9] , \blocktag[5][8] ,
         \blocktag[5][7] , \blocktag[5][6] , \blocktag[5][5] ,
         \blocktag[5][4] , \blocktag[5][3] , \blocktag[5][2] ,
         \blocktag[5][1] , \blocktag[4][24] , \blocktag[4][22] ,
         \blocktag[4][20] , \blocktag[4][18] , \blocktag[4][17] ,
         \blocktag[4][16] , \blocktag[4][15] , \blocktag[4][14] ,
         \blocktag[4][13] , \blocktag[4][12] , \blocktag[4][11] ,
         \blocktag[4][10] , \blocktag[4][9] , \blocktag[4][8] ,
         \blocktag[4][7] , \blocktag[4][6] , \blocktag[4][5] ,
         \blocktag[4][4] , \blocktag[4][3] , \blocktag[4][2] ,
         \blocktag[4][1] , \blocktag[3][20] , \blocktag[3][19] ,
         \blocktag[3][18] , \blocktag[3][17] , \blocktag[3][16] ,
         \blocktag[3][15] , \blocktag[3][14] , \blocktag[3][13] ,
         \blocktag[3][12] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][9] , \blocktag[3][8] , \blocktag[3][7] ,
         \blocktag[3][6] , \blocktag[3][5] , \blocktag[3][4] ,
         \blocktag[3][3] , \blocktag[3][2] , \blocktag[3][1] ,
         \blocktag[3][0] , \blocktag[2][20] , \blocktag[2][19] ,
         \blocktag[2][18] , \blocktag[2][17] , \blocktag[2][16] ,
         \blocktag[2][15] , \blocktag[2][14] , \blocktag[2][13] ,
         \blocktag[2][12] , \blocktag[2][11] , \blocktag[2][10] ,
         \blocktag[2][9] , \blocktag[2][8] , \blocktag[2][7] ,
         \blocktag[2][6] , \blocktag[2][5] , \blocktag[2][4] ,
         \blocktag[2][3] , \blocktag[2][2] , \blocktag[2][1] ,
         \blocktag[2][0] , \blocktag[1][20] , \blocktag[1][19] ,
         \blocktag[1][18] , \blocktag[1][17] , \blocktag[1][16] ,
         \blocktag[1][15] , \blocktag[1][14] , \blocktag[1][13] ,
         \blocktag[1][12] , \blocktag[1][11] , \blocktag[1][10] ,
         \blocktag[1][9] , \blocktag[1][8] , \blocktag[1][7] ,
         \blocktag[1][6] , \blocktag[1][5] , \blocktag[1][4] ,
         \blocktag[1][3] , \blocktag[1][2] , \blocktag[1][1] ,
         \blocktag[1][0] , \blocktag[0][20] , \blocktag[0][19] ,
         \blocktag[0][18] , \blocktag[0][17] , \blocktag[0][16] ,
         \blocktag[0][15] , \blocktag[0][14] , \blocktag[0][13] ,
         \blocktag[0][12] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][9] , \blocktag[0][8] , \blocktag[0][7] ,
         \blocktag[0][6] , \blocktag[0][5] , \blocktag[0][4] ,
         \blocktag[0][3] , \blocktag[0][2] , \blocktag[0][1] ,
         \blocktag[0][0] , valid, dirty, \block[7][127] , \block[7][126] ,
         \block[7][125] , \block[7][124] , \block[7][123] , \block[7][122] ,
         \block[7][121] , \block[7][120] , \block[7][119] , \block[7][118] ,
         \block[7][117] , \block[7][116] , \block[7][115] , \block[7][114] ,
         \block[7][113] , \block[7][112] , \block[7][111] , \block[7][110] ,
         \block[7][109] , \block[7][108] , \block[7][107] , \block[7][106] ,
         \block[7][105] , \block[7][104] , \block[7][103] , \block[7][102] ,
         \block[7][101] , \block[7][100] , \block[7][99] , \block[7][98] ,
         \block[7][97] , \block[7][96] , \block[7][95] , \block[7][94] ,
         \block[7][93] , \block[7][92] , \block[7][91] , \block[7][90] ,
         \block[7][89] , \block[7][88] , \block[7][87] , \block[7][86] ,
         \block[7][85] , \block[7][84] , \block[7][83] , \block[7][82] ,
         \block[7][81] , \block[7][80] , \block[7][79] , \block[7][78] ,
         \block[7][77] , \block[7][76] , \block[7][75] , \block[7][74] ,
         \block[7][73] , \block[7][72] , \block[7][71] , \block[7][70] ,
         \block[7][69] , \block[7][68] , \block[7][67] , \block[7][66] ,
         \block[7][65] , \block[7][64] , \block[7][63] , \block[7][62] ,
         \block[7][61] , \block[7][60] , \block[7][59] , \block[7][58] ,
         \block[7][57] , \block[7][56] , \block[7][55] , \block[7][54] ,
         \block[7][53] , \block[7][52] , \block[7][51] , \block[7][50] ,
         \block[7][49] , \block[7][48] , \block[7][47] , \block[7][46] ,
         \block[7][45] , \block[7][44] , \block[7][43] , \block[7][42] ,
         \block[7][41] , \block[7][40] , \block[7][39] , \block[7][38] ,
         \block[7][37] , \block[7][36] , \block[7][35] , \block[7][34] ,
         \block[7][33] , \block[7][32] , \block[7][31] , \block[7][30] ,
         \block[7][29] , \block[7][28] , \block[7][27] , \block[7][26] ,
         \block[7][25] , \block[7][24] , \block[7][23] , \block[7][22] ,
         \block[7][21] , \block[7][20] , \block[7][19] , \block[7][18] ,
         \block[7][17] , \block[7][16] , \block[7][15] , \block[7][14] ,
         \block[7][13] , \block[7][12] , \block[7][11] , \block[7][10] ,
         \block[7][9] , \block[7][8] , \block[7][7] , \block[7][6] ,
         \block[7][5] , \block[7][4] , \block[7][3] , \block[7][2] ,
         \block[7][1] , \block[7][0] , \block[6][127] , \block[6][126] ,
         \block[6][125] , \block[6][124] , \block[6][123] , \block[6][122] ,
         \block[6][121] , \block[6][120] , \block[6][119] , \block[6][118] ,
         \block[6][117] , \block[6][116] , \block[6][115] , \block[6][114] ,
         \block[6][113] , \block[6][112] , \block[6][111] , \block[6][110] ,
         \block[6][109] , \block[6][108] , \block[6][107] , \block[6][106] ,
         \block[6][105] , \block[6][104] , \block[6][103] , \block[6][102] ,
         \block[6][101] , \block[6][100] , \block[6][99] , \block[6][98] ,
         \block[6][97] , \block[6][96] , \block[6][95] , \block[6][94] ,
         \block[6][93] , \block[6][92] , \block[6][91] , \block[6][90] ,
         \block[6][89] , \block[6][88] , \block[6][87] , \block[6][86] ,
         \block[6][85] , \block[6][84] , \block[6][83] , \block[6][82] ,
         \block[6][81] , \block[6][80] , \block[6][79] , \block[6][78] ,
         \block[6][77] , \block[6][76] , \block[6][75] , \block[6][74] ,
         \block[6][73] , \block[6][72] , \block[6][71] , \block[6][70] ,
         \block[6][69] , \block[6][68] , \block[6][67] , \block[6][66] ,
         \block[6][65] , \block[6][64] , \block[6][63] , \block[6][62] ,
         \block[6][61] , \block[6][60] , \block[6][59] , \block[6][58] ,
         \block[6][57] , \block[6][56] , \block[6][55] , \block[6][54] ,
         \block[6][53] , \block[6][52] , \block[6][51] , \block[6][50] ,
         \block[6][49] , \block[6][48] , \block[6][47] , \block[6][46] ,
         \block[6][45] , \block[6][44] , \block[6][43] , \block[6][42] ,
         \block[6][41] , \block[6][40] , \block[6][39] , \block[6][38] ,
         \block[6][37] , \block[6][36] , \block[6][35] , \block[6][34] ,
         \block[6][33] , \block[6][32] , \block[6][31] , \block[6][30] ,
         \block[6][29] , \block[6][28] , \block[6][27] , \block[6][26] ,
         \block[6][25] , \block[6][24] , \block[6][23] , \block[6][22] ,
         \block[6][21] , \block[6][20] , \block[6][19] , \block[6][18] ,
         \block[6][17] , \block[6][16] , \block[6][15] , \block[6][14] ,
         \block[6][13] , \block[6][12] , \block[6][11] , \block[6][10] ,
         \block[6][9] , \block[6][8] , \block[6][7] , \block[6][6] ,
         \block[6][5] , \block[6][4] , \block[6][3] , \block[6][2] ,
         \block[6][1] , \block[6][0] , \block[5][127] , \block[5][126] ,
         \block[5][125] , \block[5][124] , \block[5][123] , \block[5][122] ,
         \block[5][121] , \block[5][120] , \block[5][119] , \block[5][118] ,
         \block[5][117] , \block[5][116] , \block[5][115] , \block[5][114] ,
         \block[5][113] , \block[5][112] , \block[5][111] , \block[5][110] ,
         \block[5][109] , \block[5][108] , \block[5][107] , \block[5][106] ,
         \block[5][105] , \block[5][104] , \block[5][103] , \block[5][102] ,
         \block[5][101] , \block[5][100] , \block[5][99] , \block[5][98] ,
         \block[5][97] , \block[5][96] , \block[5][95] , \block[5][94] ,
         \block[5][93] , \block[5][92] , \block[5][91] , \block[5][90] ,
         \block[5][89] , \block[5][88] , \block[5][87] , \block[5][86] ,
         \block[5][85] , \block[5][84] , \block[5][83] , \block[5][82] ,
         \block[5][81] , \block[5][80] , \block[5][79] , \block[5][78] ,
         \block[5][77] , \block[5][76] , \block[5][75] , \block[5][74] ,
         \block[5][73] , \block[5][72] , \block[5][71] , \block[5][70] ,
         \block[5][69] , \block[5][68] , \block[5][67] , \block[5][66] ,
         \block[5][65] , \block[5][64] , \block[5][63] , \block[5][62] ,
         \block[5][61] , \block[5][60] , \block[5][59] , \block[5][58] ,
         \block[5][57] , \block[5][56] , \block[5][55] , \block[5][54] ,
         \block[5][53] , \block[5][52] , \block[5][51] , \block[5][50] ,
         \block[5][49] , \block[5][48] , \block[5][47] , \block[5][46] ,
         \block[5][45] , \block[5][44] , \block[5][43] , \block[5][42] ,
         \block[5][41] , \block[5][40] , \block[5][39] , \block[5][38] ,
         \block[5][37] , \block[5][36] , \block[5][35] , \block[5][34] ,
         \block[5][33] , \block[5][32] , \block[5][31] , \block[5][30] ,
         \block[5][29] , \block[5][28] , \block[5][27] , \block[5][26] ,
         \block[5][25] , \block[5][24] , \block[5][23] , \block[5][22] ,
         \block[5][21] , \block[5][20] , \block[5][19] , \block[5][18] ,
         \block[5][17] , \block[5][16] , \block[5][15] , \block[5][14] ,
         \block[5][13] , \block[5][12] , \block[5][11] , \block[5][10] ,
         \block[5][9] , \block[5][8] , \block[5][7] , \block[5][6] ,
         \block[5][5] , \block[5][4] , \block[5][3] , \block[5][2] ,
         \block[5][1] , \block[5][0] , \block[4][127] , \block[4][126] ,
         \block[4][125] , \block[4][124] , \block[4][123] , \block[4][122] ,
         \block[4][121] , \block[4][120] , \block[4][119] , \block[4][118] ,
         \block[4][117] , \block[4][116] , \block[4][115] , \block[4][114] ,
         \block[4][113] , \block[4][112] , \block[4][111] , \block[4][110] ,
         \block[4][109] , \block[4][108] , \block[4][107] , \block[4][106] ,
         \block[4][105] , \block[4][104] , \block[4][103] , \block[4][102] ,
         \block[4][101] , \block[4][100] , \block[4][99] , \block[4][98] ,
         \block[4][97] , \block[4][96] , \block[4][95] , \block[4][94] ,
         \block[4][93] , \block[4][92] , \block[4][91] , \block[4][90] ,
         \block[4][89] , \block[4][88] , \block[4][87] , \block[4][86] ,
         \block[4][85] , \block[4][84] , \block[4][83] , \block[4][82] ,
         \block[4][81] , \block[4][80] , \block[4][79] , \block[4][78] ,
         \block[4][77] , \block[4][76] , \block[4][75] , \block[4][74] ,
         \block[4][73] , \block[4][72] , \block[4][71] , \block[4][70] ,
         \block[4][69] , \block[4][68] , \block[4][67] , \block[4][66] ,
         \block[4][65] , \block[4][64] , \block[4][63] , \block[4][62] ,
         \block[4][61] , \block[4][60] , \block[4][59] , \block[4][58] ,
         \block[4][57] , \block[4][56] , \block[4][55] , \block[4][54] ,
         \block[4][53] , \block[4][52] , \block[4][51] , \block[4][50] ,
         \block[4][49] , \block[4][48] , \block[4][47] , \block[4][46] ,
         \block[4][45] , \block[4][44] , \block[4][43] , \block[4][42] ,
         \block[4][41] , \block[4][40] , \block[4][39] , \block[4][38] ,
         \block[4][37] , \block[4][36] , \block[4][35] , \block[4][34] ,
         \block[4][33] , \block[4][32] , \block[4][31] , \block[4][30] ,
         \block[4][29] , \block[4][28] , \block[4][27] , \block[4][26] ,
         \block[4][25] , \block[4][24] , \block[4][23] , \block[4][22] ,
         \block[4][21] , \block[4][20] , \block[4][19] , \block[4][18] ,
         \block[4][17] , \block[4][16] , \block[4][15] , \block[4][14] ,
         \block[4][13] , \block[4][12] , \block[4][11] , \block[4][10] ,
         \block[4][9] , \block[4][8] , \block[4][7] , \block[4][6] ,
         \block[4][5] , \block[4][4] , \block[4][3] , \block[4][2] ,
         \block[4][1] , \block[4][0] , \block[3][127] , \block[3][126] ,
         \block[3][125] , \block[3][124] , \block[3][123] , \block[3][122] ,
         \block[3][121] , \block[3][120] , \block[3][119] , \block[3][118] ,
         \block[3][117] , \block[3][116] , \block[3][115] , \block[3][114] ,
         \block[3][113] , \block[3][112] , \block[3][111] , \block[3][110] ,
         \block[3][109] , \block[3][108] , \block[3][107] , \block[3][106] ,
         \block[3][105] , \block[3][104] , \block[3][103] , \block[3][102] ,
         \block[3][101] , \block[3][100] , \block[3][99] , \block[3][98] ,
         \block[3][97] , \block[3][96] , \block[3][95] , \block[3][94] ,
         \block[3][93] , \block[3][92] , \block[3][91] , \block[3][90] ,
         \block[3][89] , \block[3][88] , \block[3][87] , \block[3][86] ,
         \block[3][85] , \block[3][84] , \block[3][83] , \block[3][82] ,
         \block[3][81] , \block[3][80] , \block[3][79] , \block[3][78] ,
         \block[3][77] , \block[3][76] , \block[3][75] , \block[3][74] ,
         \block[3][73] , \block[3][72] , \block[3][71] , \block[3][70] ,
         \block[3][69] , \block[3][68] , \block[3][67] , \block[3][66] ,
         \block[3][65] , \block[3][64] , \block[3][63] , \block[3][62] ,
         \block[3][61] , \block[3][60] , \block[3][59] , \block[3][58] ,
         \block[3][57] , \block[3][56] , \block[3][55] , \block[3][54] ,
         \block[3][53] , \block[3][52] , \block[3][51] , \block[3][50] ,
         \block[3][49] , \block[3][48] , \block[3][47] , \block[3][46] ,
         \block[3][45] , \block[3][44] , \block[3][43] , \block[3][42] ,
         \block[3][41] , \block[3][40] , \block[3][39] , \block[3][38] ,
         \block[3][37] , \block[3][36] , \block[3][35] , \block[3][34] ,
         \block[3][33] , \block[3][32] , \block[3][31] , \block[3][30] ,
         \block[3][29] , \block[3][28] , \block[3][27] , \block[3][26] ,
         \block[3][25] , \block[3][24] , \block[3][23] , \block[3][22] ,
         \block[3][21] , \block[3][20] , \block[3][19] , \block[3][18] ,
         \block[3][17] , \block[3][16] , \block[3][15] , \block[3][14] ,
         \block[3][13] , \block[3][12] , \block[3][11] , \block[3][10] ,
         \block[3][9] , \block[3][8] , \block[3][7] , \block[3][6] ,
         \block[3][5] , \block[3][4] , \block[3][3] , \block[3][2] ,
         \block[3][1] , \block[3][0] , \block[2][127] , \block[2][126] ,
         \block[2][125] , \block[2][124] , \block[2][123] , \block[2][122] ,
         \block[2][121] , \block[2][120] , \block[2][119] , \block[2][118] ,
         \block[2][117] , \block[2][116] , \block[2][115] , \block[2][114] ,
         \block[2][113] , \block[2][112] , \block[2][111] , \block[2][110] ,
         \block[2][109] , \block[2][108] , \block[2][107] , \block[2][106] ,
         \block[2][105] , \block[2][104] , \block[2][103] , \block[2][102] ,
         \block[2][101] , \block[2][100] , \block[2][99] , \block[2][98] ,
         \block[2][97] , \block[2][96] , \block[2][95] , \block[2][94] ,
         \block[2][93] , \block[2][92] , \block[2][91] , \block[2][90] ,
         \block[2][89] , \block[2][88] , \block[2][87] , \block[2][86] ,
         \block[2][85] , \block[2][84] , \block[2][83] , \block[2][82] ,
         \block[2][81] , \block[2][80] , \block[2][79] , \block[2][78] ,
         \block[2][77] , \block[2][76] , \block[2][75] , \block[2][74] ,
         \block[2][73] , \block[2][72] , \block[2][71] , \block[2][70] ,
         \block[2][69] , \block[2][68] , \block[2][67] , \block[2][66] ,
         \block[2][65] , \block[2][64] , \block[2][63] , \block[2][62] ,
         \block[2][61] , \block[2][60] , \block[2][59] , \block[2][58] ,
         \block[2][57] , \block[2][56] , \block[2][55] , \block[2][54] ,
         \block[2][53] , \block[2][52] , \block[2][51] , \block[2][50] ,
         \block[2][49] , \block[2][48] , \block[2][47] , \block[2][46] ,
         \block[2][45] , \block[2][44] , \block[2][43] , \block[2][42] ,
         \block[2][41] , \block[2][40] , \block[2][39] , \block[2][38] ,
         \block[2][37] , \block[2][36] , \block[2][35] , \block[2][34] ,
         \block[2][33] , \block[2][32] , \block[2][31] , \block[2][30] ,
         \block[2][29] , \block[2][28] , \block[2][27] , \block[2][26] ,
         \block[2][25] , \block[2][24] , \block[2][23] , \block[2][22] ,
         \block[2][21] , \block[2][20] , \block[2][19] , \block[2][18] ,
         \block[2][17] , \block[2][16] , \block[2][15] , \block[2][14] ,
         \block[2][13] , \block[2][12] , \block[2][11] , \block[2][10] ,
         \block[2][9] , \block[2][8] , \block[2][7] , \block[2][6] ,
         \block[2][5] , \block[2][4] , \block[2][3] , \block[2][2] ,
         \block[2][1] , \block[2][0] , \block[1][127] , \block[1][126] ,
         \block[1][125] , \block[1][124] , \block[1][123] , \block[1][122] ,
         \block[1][121] , \block[1][120] , \block[1][119] , \block[1][118] ,
         \block[1][117] , \block[1][116] , \block[1][115] , \block[1][114] ,
         \block[1][113] , \block[1][112] , \block[1][111] , \block[1][110] ,
         \block[1][109] , \block[1][108] , \block[1][107] , \block[1][106] ,
         \block[1][105] , \block[1][104] , \block[1][103] , \block[1][102] ,
         \block[1][101] , \block[1][100] , \block[1][99] , \block[1][98] ,
         \block[1][97] , \block[1][96] , \block[1][95] , \block[1][94] ,
         \block[1][93] , \block[1][92] , \block[1][91] , \block[1][90] ,
         \block[1][89] , \block[1][88] , \block[1][87] , \block[1][86] ,
         \block[1][85] , \block[1][84] , \block[1][83] , \block[1][82] ,
         \block[1][81] , \block[1][80] , \block[1][79] , \block[1][78] ,
         \block[1][77] , \block[1][76] , \block[1][75] , \block[1][74] ,
         \block[1][73] , \block[1][72] , \block[1][71] , \block[1][70] ,
         \block[1][69] , \block[1][68] , \block[1][67] , \block[1][66] ,
         \block[1][65] , \block[1][64] , \block[1][63] , \block[1][62] ,
         \block[1][61] , \block[1][60] , \block[1][59] , \block[1][58] ,
         \block[1][57] , \block[1][56] , \block[1][55] , \block[1][54] ,
         \block[1][53] , \block[1][52] , \block[1][51] , \block[1][50] ,
         \block[1][49] , \block[1][48] , \block[1][47] , \block[1][46] ,
         \block[1][45] , \block[1][44] , \block[1][43] , \block[1][42] ,
         \block[1][41] , \block[1][40] , \block[1][39] , \block[1][38] ,
         \block[1][37] , \block[1][36] , \block[1][35] , \block[1][34] ,
         \block[1][33] , \block[1][32] , \block[1][31] , \block[1][30] ,
         \block[1][29] , \block[1][28] , \block[1][27] , \block[1][26] ,
         \block[1][25] , \block[1][24] , \block[1][23] , \block[1][22] ,
         \block[1][21] , \block[1][20] , \block[1][19] , \block[1][18] ,
         \block[1][17] , \block[1][16] , \block[1][15] , \block[1][14] ,
         \block[1][13] , \block[1][12] , \block[1][11] , \block[1][10] ,
         \block[1][9] , \block[1][8] , \block[1][7] , \block[1][6] ,
         \block[1][5] , \block[1][4] , \block[1][3] , \block[1][2] ,
         \block[1][1] , \block[1][0] , \block[0][127] , \block[0][126] ,
         \block[0][125] , \block[0][124] , \block[0][123] , \block[0][122] ,
         \block[0][121] , \block[0][120] , \block[0][119] , \block[0][118] ,
         \block[0][117] , \block[0][116] , \block[0][115] , \block[0][114] ,
         \block[0][113] , \block[0][112] , \block[0][111] , \block[0][110] ,
         \block[0][109] , \block[0][108] , \block[0][107] , \block[0][106] ,
         \block[0][105] , \block[0][104] , \block[0][103] , \block[0][102] ,
         \block[0][101] , \block[0][100] , \block[0][99] , \block[0][98] ,
         \block[0][97] , \block[0][96] , \block[0][95] , \block[0][94] ,
         \block[0][93] , \block[0][92] , \block[0][91] , \block[0][90] ,
         \block[0][89] , \block[0][88] , \block[0][87] , \block[0][86] ,
         \block[0][85] , \block[0][84] , \block[0][83] , \block[0][82] ,
         \block[0][81] , \block[0][80] , \block[0][79] , \block[0][78] ,
         \block[0][77] , \block[0][76] , \block[0][75] , \block[0][74] ,
         \block[0][73] , \block[0][72] , \block[0][71] , \block[0][70] ,
         \block[0][69] , \block[0][68] , \block[0][67] , \block[0][66] ,
         \block[0][65] , \block[0][64] , \block[0][63] , \block[0][62] ,
         \block[0][61] , \block[0][60] , \block[0][59] , \block[0][58] ,
         \block[0][57] , \block[0][56] , \block[0][55] , \block[0][54] ,
         \block[0][53] , \block[0][52] , \block[0][51] , \block[0][50] ,
         \block[0][49] , \block[0][48] , \block[0][47] , \block[0][46] ,
         \block[0][45] , \block[0][44] , \block[0][43] , \block[0][42] ,
         \block[0][41] , \block[0][40] , \block[0][39] , \block[0][38] ,
         \block[0][37] , \block[0][36] , \block[0][35] , \block[0][34] ,
         \block[0][33] , \block[0][32] , \block[0][31] , \block[0][30] ,
         \block[0][29] , \block[0][28] , \block[0][27] , \block[0][26] ,
         \block[0][25] , \block[0][24] , \block[0][23] , \block[0][22] ,
         \block[0][21] , \block[0][20] , \block[0][19] , \block[0][18] ,
         \block[0][17] , \block[0][16] , \block[0][15] , \block[0][14] ,
         \block[0][13] , \block[0][12] , \block[0][11] , \block[0][10] ,
         \block[0][9] , \block[0][8] , \block[0][7] , \block[0][6] ,
         \block[0][5] , \block[0][4] , \block[0][3] , \block[0][2] ,
         \block[0][1] , \block[0][0] , N1768, N1769, N1771, N1772, N1773,
         N1774, N1776, N1777, n9, n11, n13, n14, n15, n19, n23, n27, n31, n35,
         n39, n43, n47, n51, n55, n59, n63, n67, n71, n75, n79, n83, n87, n91,
         n95, n99, n103, n107, n111, n115, n119, n123, n127, n131, n135, n139,
         n143, n144, n145, n147, n148, n150, n152, n154, n156, n158, n160,
         n162, n163, n164, n165, n166, n215, n255, n256, n257, n259, n260,
         n261, n262, n263, n266, n267, n276, n277, n340, n341, n342, n430,
         n431, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n503, n504, n505, n506, n508, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  EDFFX1 \block_reg[7][127]  ( .D(block_next[127]), .E(n1095), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFX1 \block_reg[7][126]  ( .D(block_next[126]), .E(n1095), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFX1 \block_reg[7][125]  ( .D(block_next[125]), .E(n1095), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFX1 \block_reg[7][124]  ( .D(block_next[124]), .E(n1099), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFX1 \block_reg[7][123]  ( .D(block_next[123]), .E(n1097), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFX1 \block_reg[7][122]  ( .D(block_next[122]), .E(n1096), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFX1 \block_reg[7][121]  ( .D(block_next[121]), .E(n1098), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFX1 \block_reg[7][120]  ( .D(block_next[120]), .E(n1098), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFX1 \block_reg[7][119]  ( .D(block_next[119]), .E(n1100), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFX1 \block_reg[7][118]  ( .D(block_next[118]), .E(n1101), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFX1 \block_reg[7][117]  ( .D(block_next[117]), .E(n1103), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFX1 \block_reg[7][116]  ( .D(block_next[116]), .E(n1101), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFX1 \block_reg[7][115]  ( .D(block_next[115]), .E(n1103), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFX1 \block_reg[7][114]  ( .D(block_next[114]), .E(n1102), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFX1 \block_reg[7][113]  ( .D(block_next[113]), .E(n1095), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFX1 \block_reg[7][112]  ( .D(block_next[112]), .E(n1095), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFX1 \block_reg[7][111]  ( .D(block_next[111]), .E(n1099), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFX1 \block_reg[7][110]  ( .D(block_next[110]), .E(n1097), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFX1 \block_reg[7][109]  ( .D(block_next[109]), .E(n1096), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFX1 \block_reg[7][108]  ( .D(block_next[108]), .E(n1098), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFX1 \block_reg[7][107]  ( .D(block_next[107]), .E(n1100), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFX1 \block_reg[7][106]  ( .D(block_next[106]), .E(n1100), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFX1 \block_reg[7][105]  ( .D(block_next[105]), .E(n1101), .CK(clk), .Q(
        \block[7][105] ) );
  EDFFX1 \block_reg[7][104]  ( .D(block_next[104]), .E(n1103), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFX1 \block_reg[7][103]  ( .D(block_next[103]), .E(n1102), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFX1 \block_reg[7][102]  ( .D(block_next[102]), .E(n1102), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFX1 \block_reg[7][101]  ( .D(block_next[101]), .E(n1102), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFX1 \block_reg[7][100]  ( .D(block_next[100]), .E(n1102), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFX1 \block_reg[7][99]  ( .D(block_next[99]), .E(n1102), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFX1 \block_reg[7][98]  ( .D(block_next[98]), .E(n1102), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFX1 \block_reg[7][97]  ( .D(block_next[97]), .E(n1102), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFX1 \block_reg[7][96]  ( .D(block_next[96]), .E(n1102), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFX1 \block_reg[7][95]  ( .D(block_next[95]), .E(n1102), .CK(clk), .Q(
        \block[7][95] ) );
  EDFFX1 \block_reg[7][94]  ( .D(block_next[94]), .E(n1102), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFX1 \block_reg[7][93]  ( .D(block_next[93]), .E(n1102), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFX1 \block_reg[7][92]  ( .D(block_next[92]), .E(n1102), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFX1 \block_reg[7][91]  ( .D(block_next[91]), .E(n1102), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFX1 \block_reg[7][90]  ( .D(block_next[90]), .E(n1101), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFX1 \block_reg[7][89]  ( .D(block_next[89]), .E(n1101), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFX1 \block_reg[7][88]  ( .D(block_next[88]), .E(n1101), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFX1 \block_reg[7][87]  ( .D(block_next[87]), .E(n1101), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFX1 \block_reg[7][86]  ( .D(block_next[86]), .E(n1101), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFX1 \block_reg[7][85]  ( .D(block_next[85]), .E(n1101), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFX1 \block_reg[7][84]  ( .D(block_next[84]), .E(n1101), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFX1 \block_reg[7][83]  ( .D(block_next[83]), .E(n1101), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFX1 \block_reg[7][82]  ( .D(block_next[82]), .E(n1101), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFX1 \block_reg[7][81]  ( .D(block_next[81]), .E(n1101), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFX1 \block_reg[7][80]  ( .D(block_next[80]), .E(n1101), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFX1 \block_reg[7][79]  ( .D(block_next[79]), .E(n1101), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFX1 \block_reg[7][78]  ( .D(block_next[78]), .E(n1101), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFX1 \block_reg[7][77]  ( .D(block_next[77]), .E(n1102), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFX1 \block_reg[7][76]  ( .D(block_next[76]), .E(n1099), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFX1 \block_reg[7][75]  ( .D(block_next[75]), .E(n1097), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFX1 \block_reg[7][74]  ( .D(block_next[74]), .E(n1096), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFX1 \block_reg[7][73]  ( .D(block_next[73]), .E(n1098), .CK(clk), .Q(
        \block[7][73] ) );
  EDFFX1 \block_reg[7][72]  ( .D(block_next[72]), .E(n1100), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFX1 \block_reg[7][71]  ( .D(block_next[71]), .E(n1101), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFX1 \block_reg[7][70]  ( .D(block_next[70]), .E(n1103), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFX1 \block_reg[7][69]  ( .D(block_next[69]), .E(n1102), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFX1 \block_reg[7][68]  ( .D(block_next[68]), .E(n1095), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFX1 \block_reg[7][67]  ( .D(block_next[67]), .E(n1099), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFX1 \block_reg[7][66]  ( .D(block_next[66]), .E(n1097), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFX1 \block_reg[7][65]  ( .D(block_next[65]), .E(n1096), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFX1 \block_reg[7][64]  ( .D(block_next[64]), .E(n1100), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFX1 \block_reg[7][63]  ( .D(block_next[63]), .E(n1100), .CK(clk), .Q(
        \block[7][63] ) );
  EDFFX1 \block_reg[7][62]  ( .D(block_next[62]), .E(n1100), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFX1 \block_reg[7][61]  ( .D(block_next[61]), .E(n1100), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFX1 \block_reg[7][60]  ( .D(block_next[60]), .E(n1100), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFX1 \block_reg[7][59]  ( .D(block_next[59]), .E(n1100), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFX1 \block_reg[7][58]  ( .D(block_next[58]), .E(n1100), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFX1 \block_reg[7][57]  ( .D(block_next[57]), .E(n1100), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFX1 \block_reg[7][56]  ( .D(block_next[56]), .E(n1100), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFX1 \block_reg[7][55]  ( .D(block_next[55]), .E(n1100), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFX1 \block_reg[7][54]  ( .D(block_next[54]), .E(n1100), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n1100), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n1100), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[7][51]  ( .D(block_next[51]), .E(n1099), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFX1 \block_reg[7][50]  ( .D(block_next[50]), .E(n1099), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n1099), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[7][48]  ( .D(block_next[48]), .E(n1099), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFX1 \block_reg[7][47]  ( .D(block_next[47]), .E(n1099), .CK(clk), .Q(
        \block[7][47] ) );
  EDFFX1 \block_reg[7][46]  ( .D(block_next[46]), .E(n1099), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFX1 \block_reg[7][45]  ( .D(block_next[45]), .E(n1099), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFX1 \block_reg[7][44]  ( .D(block_next[44]), .E(n1099), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFX1 \block_reg[7][43]  ( .D(block_next[43]), .E(n1099), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFX1 \block_reg[7][42]  ( .D(block_next[42]), .E(n1099), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n1099), .CK(clk), .Q(
        \block[7][41] ) );
  EDFFX1 \block_reg[7][40]  ( .D(block_next[40]), .E(n1099), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFX1 \block_reg[7][39]  ( .D(block_next[39]), .E(n1099), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n1098), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n1098), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n1098), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n1098), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n1098), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFX1 \block_reg[7][33]  ( .D(block_next[33]), .E(n1098), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n1098), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[7][31]  ( .D(block_next[31]), .E(n1098), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFX1 \block_reg[7][30]  ( .D(block_next[30]), .E(n1098), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFX1 \block_reg[7][29]  ( .D(block_next[29]), .E(n1098), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFX1 \block_reg[7][28]  ( .D(block_next[28]), .E(n1098), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFX1 \block_reg[7][27]  ( .D(block_next[27]), .E(n1098), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFX1 \block_reg[7][26]  ( .D(block_next[26]), .E(n1098), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFX1 \block_reg[7][25]  ( .D(block_next[25]), .E(n1097), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFX1 \block_reg[7][24]  ( .D(block_next[24]), .E(n1097), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFX1 \block_reg[7][23]  ( .D(block_next[23]), .E(n1097), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFX1 \block_reg[7][22]  ( .D(block_next[22]), .E(n1097), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFX1 \block_reg[7][21]  ( .D(block_next[21]), .E(n1097), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFX1 \block_reg[7][20]  ( .D(block_next[20]), .E(n1097), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFX1 \block_reg[7][19]  ( .D(block_next[19]), .E(n1097), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFX1 \block_reg[7][18]  ( .D(block_next[18]), .E(n1097), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFX1 \block_reg[7][17]  ( .D(block_next[17]), .E(n1097), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFX1 \block_reg[7][16]  ( .D(block_next[16]), .E(n1097), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFX1 \block_reg[7][15]  ( .D(block_next[15]), .E(n1097), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFX1 \block_reg[7][14]  ( .D(block_next[14]), .E(n1097), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFX1 \block_reg[7][13]  ( .D(block_next[13]), .E(n1097), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFX1 \block_reg[7][12]  ( .D(block_next[12]), .E(n1096), .CK(clk), .Q(
        \block[7][12] ) );
  EDFFX1 \block_reg[7][11]  ( .D(block_next[11]), .E(n1096), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFX1 \block_reg[7][10]  ( .D(block_next[10]), .E(n1096), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFX1 \block_reg[7][9]  ( .D(block_next[9]), .E(n1096), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFX1 \block_reg[7][8]  ( .D(block_next[8]), .E(n1096), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFX1 \block_reg[7][7]  ( .D(block_next[7]), .E(n1096), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFX1 \block_reg[7][6]  ( .D(block_next[6]), .E(n1096), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFX1 \block_reg[7][5]  ( .D(block_next[5]), .E(n1096), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFX1 \block_reg[7][4]  ( .D(block_next[4]), .E(n1096), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFX1 \block_reg[7][3]  ( .D(block_next[3]), .E(n1096), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFX1 \block_reg[7][2]  ( .D(block_next[2]), .E(n1096), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFX1 \block_reg[7][1]  ( .D(block_next[1]), .E(n1096), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFX1 \block_reg[7][0]  ( .D(block_next[0]), .E(n1096), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFX1 \block_reg[3][127]  ( .D(block_next[127]), .E(n1131), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFX1 \block_reg[3][126]  ( .D(block_next[126]), .E(n1131), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFX1 \block_reg[3][125]  ( .D(block_next[125]), .E(n1131), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFX1 \block_reg[3][124]  ( .D(block_next[124]), .E(n1135), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFX1 \block_reg[3][123]  ( .D(block_next[123]), .E(n1133), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFX1 \block_reg[3][122]  ( .D(block_next[122]), .E(n1132), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFX1 \block_reg[3][121]  ( .D(block_next[121]), .E(n1134), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFX1 \block_reg[3][120]  ( .D(block_next[120]), .E(n1134), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFX1 \block_reg[3][119]  ( .D(block_next[119]), .E(n1136), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFX1 \block_reg[3][118]  ( .D(block_next[118]), .E(n1137), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFX1 \block_reg[3][117]  ( .D(block_next[117]), .E(n1139), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFX1 \block_reg[3][116]  ( .D(block_next[116]), .E(n1137), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFX1 \block_reg[3][115]  ( .D(block_next[115]), .E(n1139), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFX1 \block_reg[3][114]  ( .D(block_next[114]), .E(n1138), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFX1 \block_reg[3][113]  ( .D(block_next[113]), .E(n1131), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFX1 \block_reg[3][112]  ( .D(block_next[112]), .E(n1131), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFX1 \block_reg[3][111]  ( .D(block_next[111]), .E(n1135), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFX1 \block_reg[3][110]  ( .D(block_next[110]), .E(n1133), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFX1 \block_reg[3][109]  ( .D(block_next[109]), .E(n1132), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFX1 \block_reg[3][108]  ( .D(block_next[108]), .E(n1134), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFX1 \block_reg[3][107]  ( .D(block_next[107]), .E(n1136), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFX1 \block_reg[3][106]  ( .D(block_next[106]), .E(n1136), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFX1 \block_reg[3][105]  ( .D(block_next[105]), .E(n1137), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFX1 \block_reg[3][104]  ( .D(block_next[104]), .E(n1139), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFX1 \block_reg[3][103]  ( .D(block_next[103]), .E(n1138), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFX1 \block_reg[3][102]  ( .D(block_next[102]), .E(n1138), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFX1 \block_reg[3][101]  ( .D(block_next[101]), .E(n1138), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFX1 \block_reg[3][100]  ( .D(block_next[100]), .E(n1138), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFX1 \block_reg[3][99]  ( .D(block_next[99]), .E(n1138), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFX1 \block_reg[3][98]  ( .D(block_next[98]), .E(n1138), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFX1 \block_reg[3][97]  ( .D(block_next[97]), .E(n1138), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFX1 \block_reg[3][96]  ( .D(block_next[96]), .E(n1138), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFX1 \block_reg[3][95]  ( .D(block_next[95]), .E(n1138), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFX1 \block_reg[3][94]  ( .D(block_next[94]), .E(n1138), .CK(clk), .Q(
        \block[3][94] ) );
  EDFFX1 \block_reg[3][93]  ( .D(block_next[93]), .E(n1138), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFX1 \block_reg[3][92]  ( .D(block_next[92]), .E(n1138), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFX1 \block_reg[3][91]  ( .D(block_next[91]), .E(n1138), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFX1 \block_reg[3][90]  ( .D(block_next[90]), .E(n1137), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFX1 \block_reg[3][89]  ( .D(block_next[89]), .E(n1137), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFX1 \block_reg[3][88]  ( .D(block_next[88]), .E(n1137), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFX1 \block_reg[3][87]  ( .D(block_next[87]), .E(n1137), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFX1 \block_reg[3][86]  ( .D(block_next[86]), .E(n1137), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFX1 \block_reg[3][85]  ( .D(block_next[85]), .E(n1137), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFX1 \block_reg[3][84]  ( .D(block_next[84]), .E(n1137), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFX1 \block_reg[3][83]  ( .D(block_next[83]), .E(n1137), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFX1 \block_reg[3][82]  ( .D(block_next[82]), .E(n1137), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFX1 \block_reg[3][81]  ( .D(block_next[81]), .E(n1137), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFX1 \block_reg[3][80]  ( .D(block_next[80]), .E(n1137), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFX1 \block_reg[3][79]  ( .D(block_next[79]), .E(n1137), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFX1 \block_reg[3][78]  ( .D(block_next[78]), .E(n1137), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFX1 \block_reg[3][77]  ( .D(block_next[77]), .E(n1138), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFX1 \block_reg[3][76]  ( .D(block_next[76]), .E(n1135), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFX1 \block_reg[3][75]  ( .D(block_next[75]), .E(n1133), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFX1 \block_reg[3][74]  ( .D(block_next[74]), .E(n1132), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFX1 \block_reg[3][73]  ( .D(block_next[73]), .E(n1134), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFX1 \block_reg[3][72]  ( .D(block_next[72]), .E(n1136), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFX1 \block_reg[3][71]  ( .D(block_next[71]), .E(n1137), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFX1 \block_reg[3][70]  ( .D(block_next[70]), .E(n1139), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFX1 \block_reg[3][69]  ( .D(block_next[69]), .E(n1138), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFX1 \block_reg[3][68]  ( .D(block_next[68]), .E(n1131), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFX1 \block_reg[3][67]  ( .D(block_next[67]), .E(n1135), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFX1 \block_reg[3][66]  ( .D(block_next[66]), .E(n1133), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFX1 \block_reg[3][65]  ( .D(block_next[65]), .E(n1132), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFX1 \block_reg[3][64]  ( .D(block_next[64]), .E(n1136), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[3][63]  ( .D(block_next[63]), .E(n1136), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFX1 \block_reg[3][62]  ( .D(block_next[62]), .E(n1136), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFX1 \block_reg[3][61]  ( .D(block_next[61]), .E(n1136), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFX1 \block_reg[3][60]  ( .D(block_next[60]), .E(n1136), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFX1 \block_reg[3][59]  ( .D(block_next[59]), .E(n1136), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFX1 \block_reg[3][58]  ( .D(block_next[58]), .E(n1136), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFX1 \block_reg[3][57]  ( .D(block_next[57]), .E(n1136), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFX1 \block_reg[3][56]  ( .D(block_next[56]), .E(n1136), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFX1 \block_reg[3][55]  ( .D(block_next[55]), .E(n1136), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFX1 \block_reg[3][54]  ( .D(block_next[54]), .E(n1136), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n1136), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n1136), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[3][51]  ( .D(block_next[51]), .E(n1135), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFX1 \block_reg[3][50]  ( .D(block_next[50]), .E(n1135), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n1135), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[3][48]  ( .D(block_next[48]), .E(n1135), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFX1 \block_reg[3][47]  ( .D(block_next[47]), .E(n1135), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFX1 \block_reg[3][46]  ( .D(block_next[46]), .E(n1135), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFX1 \block_reg[3][45]  ( .D(block_next[45]), .E(n1135), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFX1 \block_reg[3][44]  ( .D(block_next[44]), .E(n1135), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFX1 \block_reg[3][43]  ( .D(block_next[43]), .E(n1135), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFX1 \block_reg[3][42]  ( .D(block_next[42]), .E(n1135), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n1135), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[3][40]  ( .D(block_next[40]), .E(n1135), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFX1 \block_reg[3][39]  ( .D(block_next[39]), .E(n1135), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n1134), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n1134), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n1134), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n1134), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n1134), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[3][33]  ( .D(block_next[33]), .E(n1134), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n1134), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[3][31]  ( .D(block_next[31]), .E(n1134), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFX1 \block_reg[3][30]  ( .D(block_next[30]), .E(n1134), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFX1 \block_reg[3][29]  ( .D(block_next[29]), .E(n1134), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFX1 \block_reg[3][28]  ( .D(block_next[28]), .E(n1134), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFX1 \block_reg[3][27]  ( .D(block_next[27]), .E(n1134), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFX1 \block_reg[3][26]  ( .D(block_next[26]), .E(n1134), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFX1 \block_reg[3][25]  ( .D(block_next[25]), .E(n1133), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFX1 \block_reg[3][24]  ( .D(block_next[24]), .E(n1133), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFX1 \block_reg[3][23]  ( .D(block_next[23]), .E(n1133), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFX1 \block_reg[3][22]  ( .D(block_next[22]), .E(n1133), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFX1 \block_reg[3][21]  ( .D(block_next[21]), .E(n1133), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n1133), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFX1 \block_reg[3][19]  ( .D(block_next[19]), .E(n1133), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFX1 \block_reg[3][18]  ( .D(block_next[18]), .E(n1133), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFX1 \block_reg[3][17]  ( .D(block_next[17]), .E(n1133), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFX1 \block_reg[3][16]  ( .D(block_next[16]), .E(n1133), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFX1 \block_reg[3][15]  ( .D(block_next[15]), .E(n1133), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFX1 \block_reg[3][14]  ( .D(block_next[14]), .E(n1133), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFX1 \block_reg[3][13]  ( .D(block_next[13]), .E(n1133), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFX1 \block_reg[3][12]  ( .D(block_next[12]), .E(n1132), .CK(clk), .Q(
        \block[3][12] ) );
  EDFFX1 \block_reg[3][11]  ( .D(block_next[11]), .E(n1132), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFX1 \block_reg[3][10]  ( .D(block_next[10]), .E(n1132), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFX1 \block_reg[3][9]  ( .D(block_next[9]), .E(n1132), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFX1 \block_reg[3][8]  ( .D(block_next[8]), .E(n1132), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFX1 \block_reg[3][7]  ( .D(block_next[7]), .E(n1132), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFX1 \block_reg[3][6]  ( .D(block_next[6]), .E(n1132), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFX1 \block_reg[3][5]  ( .D(block_next[5]), .E(n1132), .CK(clk), .Q(
        \block[3][5] ) );
  EDFFX1 \block_reg[3][4]  ( .D(block_next[4]), .E(n1132), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFX1 \block_reg[3][3]  ( .D(block_next[3]), .E(n1132), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFX1 \block_reg[3][2]  ( .D(block_next[2]), .E(n1132), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFX1 \block_reg[3][1]  ( .D(block_next[1]), .E(n1132), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFX1 \block_reg[3][0]  ( .D(block_next[0]), .E(n1132), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFX1 \block_reg[5][127]  ( .D(block_next[127]), .E(n1113), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFX1 \block_reg[5][126]  ( .D(block_next[126]), .E(n1113), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFX1 \block_reg[5][125]  ( .D(block_next[125]), .E(n1113), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFX1 \block_reg[5][124]  ( .D(block_next[124]), .E(n1117), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFX1 \block_reg[5][123]  ( .D(block_next[123]), .E(n1115), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFX1 \block_reg[5][122]  ( .D(block_next[122]), .E(n1114), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFX1 \block_reg[5][121]  ( .D(block_next[121]), .E(n1116), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFX1 \block_reg[5][120]  ( .D(block_next[120]), .E(n1116), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFX1 \block_reg[5][119]  ( .D(block_next[119]), .E(n1118), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFX1 \block_reg[5][118]  ( .D(block_next[118]), .E(n1119), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFX1 \block_reg[5][117]  ( .D(block_next[117]), .E(n1121), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFX1 \block_reg[5][116]  ( .D(block_next[116]), .E(n1119), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFX1 \block_reg[5][115]  ( .D(block_next[115]), .E(n1121), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFX1 \block_reg[5][114]  ( .D(block_next[114]), .E(n1120), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFX1 \block_reg[5][113]  ( .D(block_next[113]), .E(n1113), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFX1 \block_reg[5][112]  ( .D(block_next[112]), .E(n1113), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFX1 \block_reg[5][111]  ( .D(block_next[111]), .E(n1117), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFX1 \block_reg[5][110]  ( .D(block_next[110]), .E(n1115), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFX1 \block_reg[5][109]  ( .D(block_next[109]), .E(n1114), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFX1 \block_reg[5][108]  ( .D(block_next[108]), .E(n1116), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFX1 \block_reg[5][107]  ( .D(block_next[107]), .E(n1118), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFX1 \block_reg[5][106]  ( .D(block_next[106]), .E(n1118), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFX1 \block_reg[5][105]  ( .D(block_next[105]), .E(n1119), .CK(clk), .Q(
        \block[5][105] ) );
  EDFFX1 \block_reg[5][104]  ( .D(block_next[104]), .E(n1121), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFX1 \block_reg[5][103]  ( .D(block_next[103]), .E(n1120), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFX1 \block_reg[5][102]  ( .D(block_next[102]), .E(n1120), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFX1 \block_reg[5][101]  ( .D(block_next[101]), .E(n1120), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFX1 \block_reg[5][100]  ( .D(block_next[100]), .E(n1120), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFX1 \block_reg[5][99]  ( .D(block_next[99]), .E(n1120), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFX1 \block_reg[5][98]  ( .D(block_next[98]), .E(n1120), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFX1 \block_reg[5][97]  ( .D(block_next[97]), .E(n1120), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFX1 \block_reg[5][96]  ( .D(block_next[96]), .E(n1120), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFX1 \block_reg[5][95]  ( .D(block_next[95]), .E(n1120), .CK(clk), .Q(
        \block[5][95] ) );
  EDFFX1 \block_reg[5][94]  ( .D(block_next[94]), .E(n1120), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFX1 \block_reg[5][93]  ( .D(block_next[93]), .E(n1120), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFX1 \block_reg[5][92]  ( .D(block_next[92]), .E(n1120), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFX1 \block_reg[5][91]  ( .D(block_next[91]), .E(n1120), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFX1 \block_reg[5][90]  ( .D(block_next[90]), .E(n1119), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFX1 \block_reg[5][89]  ( .D(block_next[89]), .E(n1119), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFX1 \block_reg[5][88]  ( .D(block_next[88]), .E(n1119), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFX1 \block_reg[5][87]  ( .D(block_next[87]), .E(n1119), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFX1 \block_reg[5][86]  ( .D(block_next[86]), .E(n1119), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFX1 \block_reg[5][85]  ( .D(block_next[85]), .E(n1119), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFX1 \block_reg[5][84]  ( .D(block_next[84]), .E(n1119), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFX1 \block_reg[5][83]  ( .D(block_next[83]), .E(n1119), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFX1 \block_reg[5][82]  ( .D(block_next[82]), .E(n1119), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFX1 \block_reg[5][81]  ( .D(block_next[81]), .E(n1119), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFX1 \block_reg[5][80]  ( .D(block_next[80]), .E(n1119), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFX1 \block_reg[5][79]  ( .D(block_next[79]), .E(n1119), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFX1 \block_reg[5][78]  ( .D(block_next[78]), .E(n1119), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFX1 \block_reg[5][77]  ( .D(block_next[77]), .E(n1120), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFX1 \block_reg[5][76]  ( .D(block_next[76]), .E(n1117), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFX1 \block_reg[5][75]  ( .D(block_next[75]), .E(n1115), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFX1 \block_reg[5][74]  ( .D(block_next[74]), .E(n1114), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFX1 \block_reg[5][73]  ( .D(block_next[73]), .E(n1116), .CK(clk), .Q(
        \block[5][73] ) );
  EDFFX1 \block_reg[5][72]  ( .D(block_next[72]), .E(n1118), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFX1 \block_reg[5][71]  ( .D(block_next[71]), .E(n1119), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFX1 \block_reg[5][70]  ( .D(block_next[70]), .E(n1121), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFX1 \block_reg[5][69]  ( .D(block_next[69]), .E(n1120), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFX1 \block_reg[5][68]  ( .D(block_next[68]), .E(n1113), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFX1 \block_reg[5][67]  ( .D(block_next[67]), .E(n1117), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFX1 \block_reg[5][66]  ( .D(block_next[66]), .E(n1115), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFX1 \block_reg[5][65]  ( .D(block_next[65]), .E(n1114), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFX1 \block_reg[5][64]  ( .D(block_next[64]), .E(n1118), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFX1 \block_reg[5][63]  ( .D(block_next[63]), .E(n1118), .CK(clk), .Q(
        \block[5][63] ) );
  EDFFX1 \block_reg[5][62]  ( .D(block_next[62]), .E(n1118), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFX1 \block_reg[5][61]  ( .D(block_next[61]), .E(n1118), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFX1 \block_reg[5][60]  ( .D(block_next[60]), .E(n1118), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFX1 \block_reg[5][59]  ( .D(block_next[59]), .E(n1118), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFX1 \block_reg[5][58]  ( .D(block_next[58]), .E(n1118), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFX1 \block_reg[5][57]  ( .D(block_next[57]), .E(n1118), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFX1 \block_reg[5][56]  ( .D(block_next[56]), .E(n1118), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFX1 \block_reg[5][55]  ( .D(block_next[55]), .E(n1118), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFX1 \block_reg[5][54]  ( .D(block_next[54]), .E(n1118), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFX1 \block_reg[5][53]  ( .D(block_next[53]), .E(n1118), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFX1 \block_reg[5][52]  ( .D(block_next[52]), .E(n1118), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFX1 \block_reg[5][51]  ( .D(block_next[51]), .E(n1117), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFX1 \block_reg[5][50]  ( .D(block_next[50]), .E(n1117), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFX1 \block_reg[5][49]  ( .D(block_next[49]), .E(n1117), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFX1 \block_reg[5][48]  ( .D(block_next[48]), .E(n1117), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFX1 \block_reg[5][47]  ( .D(block_next[47]), .E(n1117), .CK(clk), .Q(
        \block[5][47] ) );
  EDFFX1 \block_reg[5][46]  ( .D(block_next[46]), .E(n1117), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFX1 \block_reg[5][45]  ( .D(block_next[45]), .E(n1117), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFX1 \block_reg[5][44]  ( .D(block_next[44]), .E(n1117), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFX1 \block_reg[5][43]  ( .D(block_next[43]), .E(n1117), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFX1 \block_reg[5][42]  ( .D(block_next[42]), .E(n1117), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n1117), .CK(clk), .Q(
        \block[5][41] ) );
  EDFFX1 \block_reg[5][40]  ( .D(block_next[40]), .E(n1117), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFX1 \block_reg[5][39]  ( .D(block_next[39]), .E(n1117), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n1116), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n1116), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n1116), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFX1 \block_reg[5][35]  ( .D(block_next[35]), .E(n1116), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFX1 \block_reg[5][34]  ( .D(block_next[34]), .E(n1116), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFX1 \block_reg[5][33]  ( .D(block_next[33]), .E(n1116), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n1116), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFX1 \block_reg[5][31]  ( .D(block_next[31]), .E(n1116), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFX1 \block_reg[5][30]  ( .D(block_next[30]), .E(n1116), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFX1 \block_reg[5][29]  ( .D(block_next[29]), .E(n1116), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFX1 \block_reg[5][28]  ( .D(block_next[28]), .E(n1116), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFX1 \block_reg[5][27]  ( .D(block_next[27]), .E(n1116), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFX1 \block_reg[5][26]  ( .D(block_next[26]), .E(n1116), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFX1 \block_reg[5][25]  ( .D(block_next[25]), .E(n1115), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFX1 \block_reg[5][24]  ( .D(block_next[24]), .E(n1115), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFX1 \block_reg[5][23]  ( .D(block_next[23]), .E(n1115), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFX1 \block_reg[5][22]  ( .D(block_next[22]), .E(n1115), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFX1 \block_reg[5][21]  ( .D(block_next[21]), .E(n1115), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[5][20]  ( .D(block_next[20]), .E(n1115), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFX1 \block_reg[5][19]  ( .D(block_next[19]), .E(n1115), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFX1 \block_reg[5][18]  ( .D(block_next[18]), .E(n1115), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFX1 \block_reg[5][17]  ( .D(block_next[17]), .E(n1115), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFX1 \block_reg[5][16]  ( .D(block_next[16]), .E(n1115), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFX1 \block_reg[5][15]  ( .D(block_next[15]), .E(n1115), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[5][14]  ( .D(block_next[14]), .E(n1115), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFX1 \block_reg[5][13]  ( .D(block_next[13]), .E(n1115), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFX1 \block_reg[5][12]  ( .D(block_next[12]), .E(n1114), .CK(clk), .Q(
        \block[5][12] ) );
  EDFFX1 \block_reg[5][11]  ( .D(block_next[11]), .E(n1114), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFX1 \block_reg[5][10]  ( .D(block_next[10]), .E(n1114), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFX1 \block_reg[5][9]  ( .D(block_next[9]), .E(n1114), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFX1 \block_reg[5][8]  ( .D(block_next[8]), .E(n1114), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFX1 \block_reg[5][7]  ( .D(block_next[7]), .E(n1114), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFX1 \block_reg[5][6]  ( .D(block_next[6]), .E(n1114), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFX1 \block_reg[5][5]  ( .D(block_next[5]), .E(n1114), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFX1 \block_reg[5][4]  ( .D(block_next[4]), .E(n1114), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFX1 \block_reg[5][3]  ( .D(block_next[3]), .E(n1114), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFX1 \block_reg[5][2]  ( .D(block_next[2]), .E(n1114), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFX1 \block_reg[5][1]  ( .D(block_next[1]), .E(n1114), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFX1 \block_reg[5][0]  ( .D(block_next[0]), .E(n1114), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFX1 \block_reg[1][127]  ( .D(block_next[127]), .E(n1156), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFX1 \block_reg[1][126]  ( .D(block_next[126]), .E(n1156), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFX1 \block_reg[1][125]  ( .D(block_next[125]), .E(n1149), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFX1 \block_reg[1][124]  ( .D(block_next[124]), .E(n1151), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFX1 \block_reg[1][123]  ( .D(block_next[123]), .E(n1156), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFX1 \block_reg[1][122]  ( .D(block_next[122]), .E(n1149), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFX1 \block_reg[1][121]  ( .D(block_next[121]), .E(n1149), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFX1 \block_reg[1][120]  ( .D(block_next[120]), .E(n1155), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFX1 \block_reg[1][119]  ( .D(block_next[119]), .E(n1156), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFX1 \block_reg[1][118]  ( .D(block_next[118]), .E(n1150), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFX1 \block_reg[1][117]  ( .D(block_next[117]), .E(n1149), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFX1 \block_reg[1][116]  ( .D(block_next[116]), .E(n1155), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFX1 \block_reg[1][115]  ( .D(block_next[115]), .E(n1155), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFX1 \block_reg[1][114]  ( .D(block_next[114]), .E(n1155), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFX1 \block_reg[1][113]  ( .D(block_next[113]), .E(n1155), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFX1 \block_reg[1][112]  ( .D(block_next[112]), .E(n1155), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFX1 \block_reg[1][111]  ( .D(block_next[111]), .E(n1155), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFX1 \block_reg[1][110]  ( .D(block_next[110]), .E(n1155), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFX1 \block_reg[1][109]  ( .D(block_next[109]), .E(n1155), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFX1 \block_reg[1][108]  ( .D(block_next[108]), .E(n1155), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFX1 \block_reg[1][107]  ( .D(block_next[107]), .E(n1155), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFX1 \block_reg[1][106]  ( .D(block_next[106]), .E(n1155), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFX1 \block_reg[1][105]  ( .D(block_next[105]), .E(n1155), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFX1 \block_reg[1][104]  ( .D(block_next[104]), .E(n1155), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFX1 \block_reg[1][103]  ( .D(block_next[103]), .E(n1154), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFX1 \block_reg[1][102]  ( .D(block_next[102]), .E(n1154), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFX1 \block_reg[1][101]  ( .D(block_next[101]), .E(n1154), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFX1 \block_reg[1][100]  ( .D(block_next[100]), .E(n1154), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFX1 \block_reg[1][99]  ( .D(block_next[99]), .E(n1154), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFX1 \block_reg[1][98]  ( .D(block_next[98]), .E(n1154), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFX1 \block_reg[1][97]  ( .D(block_next[97]), .E(n1154), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFX1 \block_reg[1][96]  ( .D(block_next[96]), .E(n1154), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFX1 \block_reg[1][95]  ( .D(block_next[95]), .E(n1154), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFX1 \block_reg[1][94]  ( .D(block_next[94]), .E(n1154), .CK(clk), .Q(
        \block[1][94] ) );
  EDFFX1 \block_reg[1][93]  ( .D(block_next[93]), .E(n1154), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFX1 \block_reg[1][92]  ( .D(block_next[92]), .E(n1154), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFX1 \block_reg[1][91]  ( .D(block_next[91]), .E(n1154), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFX1 \block_reg[1][90]  ( .D(block_next[90]), .E(n1153), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFX1 \block_reg[1][89]  ( .D(block_next[89]), .E(n1153), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFX1 \block_reg[1][88]  ( .D(block_next[88]), .E(n1153), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFX1 \block_reg[1][87]  ( .D(block_next[87]), .E(n1153), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFX1 \block_reg[1][86]  ( .D(block_next[86]), .E(n1153), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFX1 \block_reg[1][85]  ( .D(block_next[85]), .E(n1153), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFX1 \block_reg[1][84]  ( .D(block_next[84]), .E(n1153), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFX1 \block_reg[1][83]  ( .D(block_next[83]), .E(n1153), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFX1 \block_reg[1][82]  ( .D(block_next[82]), .E(n1153), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFX1 \block_reg[1][81]  ( .D(block_next[81]), .E(n1153), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFX1 \block_reg[1][80]  ( .D(block_next[80]), .E(n1153), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFX1 \block_reg[1][79]  ( .D(block_next[79]), .E(n1153), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFX1 \block_reg[1][78]  ( .D(block_next[78]), .E(n1153), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFX1 \block_reg[1][77]  ( .D(block_next[77]), .E(n1152), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFX1 \block_reg[1][76]  ( .D(block_next[76]), .E(n1152), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFX1 \block_reg[1][75]  ( .D(block_next[75]), .E(n1152), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFX1 \block_reg[1][74]  ( .D(block_next[74]), .E(n1152), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFX1 \block_reg[1][73]  ( .D(block_next[73]), .E(n1152), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFX1 \block_reg[1][72]  ( .D(block_next[72]), .E(n1152), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFX1 \block_reg[1][71]  ( .D(block_next[71]), .E(n1152), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFX1 \block_reg[1][70]  ( .D(block_next[70]), .E(n1152), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFX1 \block_reg[1][69]  ( .D(block_next[69]), .E(n1152), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFX1 \block_reg[1][68]  ( .D(block_next[68]), .E(n1152), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFX1 \block_reg[1][67]  ( .D(block_next[67]), .E(n1152), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFX1 \block_reg[1][66]  ( .D(block_next[66]), .E(n1152), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFX1 \block_reg[1][65]  ( .D(block_next[65]), .E(n1152), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFX1 \block_reg[1][64]  ( .D(block_next[64]), .E(n1151), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[1][63]  ( .D(block_next[63]), .E(n1151), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFX1 \block_reg[1][62]  ( .D(block_next[62]), .E(n1151), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFX1 \block_reg[1][61]  ( .D(block_next[61]), .E(n1151), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFX1 \block_reg[1][60]  ( .D(block_next[60]), .E(n1151), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFX1 \block_reg[1][59]  ( .D(block_next[59]), .E(n1151), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFX1 \block_reg[1][58]  ( .D(block_next[58]), .E(n1151), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFX1 \block_reg[1][57]  ( .D(block_next[57]), .E(n1151), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFX1 \block_reg[1][56]  ( .D(block_next[56]), .E(n1151), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFX1 \block_reg[1][55]  ( .D(block_next[55]), .E(n1151), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFX1 \block_reg[1][54]  ( .D(block_next[54]), .E(n1151), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n1151), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n1151), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[1][51]  ( .D(block_next[51]), .E(n1152), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFX1 \block_reg[1][50]  ( .D(block_next[50]), .E(n1153), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n1151), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[1][48]  ( .D(block_next[48]), .E(n1155), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFX1 \block_reg[1][47]  ( .D(block_next[47]), .E(n1154), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFX1 \block_reg[1][46]  ( .D(block_next[46]), .E(n1157), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFX1 \block_reg[1][45]  ( .D(block_next[45]), .E(n1157), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFX1 \block_reg[1][44]  ( .D(block_next[44]), .E(n1157), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFX1 \block_reg[1][43]  ( .D(block_next[43]), .E(n1149), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFX1 \block_reg[1][42]  ( .D(block_next[42]), .E(N1769), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFX1 \block_reg[1][41]  ( .D(block_next[41]), .E(n1156), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[1][40]  ( .D(block_next[40]), .E(n1149), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFX1 \block_reg[1][39]  ( .D(block_next[39]), .E(n1157), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFX1 \block_reg[1][38]  ( .D(block_next[38]), .E(n1151), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFX1 \block_reg[1][37]  ( .D(block_next[37]), .E(n1155), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[1][36]  ( .D(block_next[36]), .E(n1154), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(N1769), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFX1 \block_reg[1][34]  ( .D(block_next[34]), .E(n1157), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFX1 \block_reg[1][33]  ( .D(block_next[33]), .E(n1152), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFX1 \block_reg[1][32]  ( .D(block_next[32]), .E(n1153), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[1][31]  ( .D(block_next[31]), .E(n1151), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFX1 \block_reg[1][30]  ( .D(block_next[30]), .E(n1155), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFX1 \block_reg[1][29]  ( .D(block_next[29]), .E(n1154), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFX1 \block_reg[1][28]  ( .D(block_next[28]), .E(n1157), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFX1 \block_reg[1][27]  ( .D(block_next[27]), .E(n1152), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFX1 \block_reg[1][26]  ( .D(block_next[26]), .E(n1153), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFX1 \block_reg[1][25]  ( .D(block_next[25]), .E(n1150), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFX1 \block_reg[1][24]  ( .D(block_next[24]), .E(n1150), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFX1 \block_reg[1][23]  ( .D(block_next[23]), .E(n1150), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFX1 \block_reg[1][22]  ( .D(block_next[22]), .E(n1150), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFX1 \block_reg[1][21]  ( .D(block_next[21]), .E(n1150), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n1150), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFX1 \block_reg[1][19]  ( .D(block_next[19]), .E(n1150), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFX1 \block_reg[1][18]  ( .D(block_next[18]), .E(n1150), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFX1 \block_reg[1][17]  ( .D(block_next[17]), .E(n1150), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFX1 \block_reg[1][16]  ( .D(block_next[16]), .E(n1150), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFX1 \block_reg[1][15]  ( .D(block_next[15]), .E(n1150), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFX1 \block_reg[1][14]  ( .D(block_next[14]), .E(n1150), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFX1 \block_reg[1][13]  ( .D(block_next[13]), .E(n1150), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFX1 \block_reg[1][12]  ( .D(block_next[12]), .E(n1149), .CK(clk), .Q(
        \block[1][12] ) );
  EDFFX1 \block_reg[1][11]  ( .D(block_next[11]), .E(n1149), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFX1 \block_reg[1][10]  ( .D(block_next[10]), .E(n1149), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFX1 \block_reg[1][9]  ( .D(block_next[9]), .E(n1149), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFX1 \block_reg[1][8]  ( .D(block_next[8]), .E(n1149), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFX1 \block_reg[1][7]  ( .D(block_next[7]), .E(n1149), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFX1 \block_reg[1][6]  ( .D(block_next[6]), .E(n1149), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFX1 \block_reg[1][5]  ( .D(block_next[5]), .E(n1149), .CK(clk), .Q(
        \block[1][5] ) );
  EDFFX1 \block_reg[1][4]  ( .D(block_next[4]), .E(n1149), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFX1 \block_reg[1][3]  ( .D(block_next[3]), .E(n1149), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFX1 \block_reg[1][2]  ( .D(block_next[2]), .E(n1149), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFX1 \block_reg[1][1]  ( .D(block_next[1]), .E(n1149), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFX1 \block_reg[1][0]  ( .D(block_next[0]), .E(n1149), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFX1 \block_reg[4][127]  ( .D(block_next[127]), .E(n1122), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFX1 \block_reg[4][126]  ( .D(block_next[126]), .E(n1122), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFX1 \block_reg[4][125]  ( .D(block_next[125]), .E(n1122), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFX1 \block_reg[4][124]  ( .D(block_next[124]), .E(n1126), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFX1 \block_reg[4][123]  ( .D(block_next[123]), .E(n1124), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFX1 \block_reg[4][122]  ( .D(block_next[122]), .E(n1123), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFX1 \block_reg[4][121]  ( .D(block_next[121]), .E(n1125), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFX1 \block_reg[4][120]  ( .D(block_next[120]), .E(n1125), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFX1 \block_reg[4][119]  ( .D(block_next[119]), .E(n1127), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFX1 \block_reg[4][118]  ( .D(block_next[118]), .E(n1128), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFX1 \block_reg[4][117]  ( .D(block_next[117]), .E(n1130), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFX1 \block_reg[4][116]  ( .D(block_next[116]), .E(n1128), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFX1 \block_reg[4][115]  ( .D(block_next[115]), .E(n1130), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFX1 \block_reg[4][114]  ( .D(block_next[114]), .E(n1129), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFX1 \block_reg[4][113]  ( .D(block_next[113]), .E(n1122), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFX1 \block_reg[4][112]  ( .D(block_next[112]), .E(n1122), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFX1 \block_reg[4][111]  ( .D(block_next[111]), .E(n1126), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFX1 \block_reg[4][110]  ( .D(block_next[110]), .E(n1124), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFX1 \block_reg[4][109]  ( .D(block_next[109]), .E(n1123), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFX1 \block_reg[4][108]  ( .D(block_next[108]), .E(n1125), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFX1 \block_reg[4][107]  ( .D(block_next[107]), .E(n1127), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFX1 \block_reg[4][106]  ( .D(block_next[106]), .E(n1127), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFX1 \block_reg[4][105]  ( .D(block_next[105]), .E(n1128), .CK(clk), .Q(
        \block[4][105] ) );
  EDFFX1 \block_reg[4][104]  ( .D(block_next[104]), .E(n1130), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFX1 \block_reg[4][103]  ( .D(block_next[103]), .E(n1129), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFX1 \block_reg[4][102]  ( .D(block_next[102]), .E(n1129), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFX1 \block_reg[4][101]  ( .D(block_next[101]), .E(n1129), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFX1 \block_reg[4][100]  ( .D(block_next[100]), .E(n1129), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFX1 \block_reg[4][99]  ( .D(block_next[99]), .E(n1129), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFX1 \block_reg[4][98]  ( .D(block_next[98]), .E(n1129), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFX1 \block_reg[4][97]  ( .D(block_next[97]), .E(n1129), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFX1 \block_reg[4][96]  ( .D(block_next[96]), .E(n1129), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFX1 \block_reg[4][95]  ( .D(block_next[95]), .E(n1129), .CK(clk), .Q(
        \block[4][95] ) );
  EDFFX1 \block_reg[4][94]  ( .D(block_next[94]), .E(n1129), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFX1 \block_reg[4][93]  ( .D(block_next[93]), .E(n1129), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFX1 \block_reg[4][92]  ( .D(block_next[92]), .E(n1129), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFX1 \block_reg[4][91]  ( .D(block_next[91]), .E(n1129), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFX1 \block_reg[4][90]  ( .D(block_next[90]), .E(n1128), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFX1 \block_reg[4][89]  ( .D(block_next[89]), .E(n1128), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFX1 \block_reg[4][88]  ( .D(block_next[88]), .E(n1128), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFX1 \block_reg[4][87]  ( .D(block_next[87]), .E(n1128), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFX1 \block_reg[4][86]  ( .D(block_next[86]), .E(n1128), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFX1 \block_reg[4][85]  ( .D(block_next[85]), .E(n1128), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFX1 \block_reg[4][84]  ( .D(block_next[84]), .E(n1128), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFX1 \block_reg[4][83]  ( .D(block_next[83]), .E(n1128), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFX1 \block_reg[4][82]  ( .D(block_next[82]), .E(n1128), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFX1 \block_reg[4][81]  ( .D(block_next[81]), .E(n1128), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFX1 \block_reg[4][80]  ( .D(block_next[80]), .E(n1128), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFX1 \block_reg[4][79]  ( .D(block_next[79]), .E(n1128), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFX1 \block_reg[4][78]  ( .D(block_next[78]), .E(n1128), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFX1 \block_reg[4][77]  ( .D(block_next[77]), .E(n1129), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFX1 \block_reg[4][76]  ( .D(block_next[76]), .E(n1126), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFX1 \block_reg[4][75]  ( .D(block_next[75]), .E(n1124), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFX1 \block_reg[4][74]  ( .D(block_next[74]), .E(n1123), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFX1 \block_reg[4][73]  ( .D(block_next[73]), .E(n1125), .CK(clk), .Q(
        \block[4][73] ) );
  EDFFX1 \block_reg[4][72]  ( .D(block_next[72]), .E(n1127), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFX1 \block_reg[4][71]  ( .D(block_next[71]), .E(n1128), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFX1 \block_reg[4][70]  ( .D(block_next[70]), .E(n1130), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFX1 \block_reg[4][69]  ( .D(block_next[69]), .E(n1129), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFX1 \block_reg[4][68]  ( .D(block_next[68]), .E(n1122), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFX1 \block_reg[4][67]  ( .D(block_next[67]), .E(n1126), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFX1 \block_reg[4][66]  ( .D(block_next[66]), .E(n1124), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFX1 \block_reg[4][65]  ( .D(block_next[65]), .E(n1123), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFX1 \block_reg[4][64]  ( .D(block_next[64]), .E(n1127), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFX1 \block_reg[4][63]  ( .D(block_next[63]), .E(n1127), .CK(clk), .Q(
        \block[4][63] ) );
  EDFFX1 \block_reg[4][62]  ( .D(block_next[62]), .E(n1127), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFX1 \block_reg[4][61]  ( .D(block_next[61]), .E(n1127), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFX1 \block_reg[4][60]  ( .D(block_next[60]), .E(n1127), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFX1 \block_reg[4][59]  ( .D(block_next[59]), .E(n1127), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFX1 \block_reg[4][58]  ( .D(block_next[58]), .E(n1127), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFX1 \block_reg[4][57]  ( .D(block_next[57]), .E(n1127), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFX1 \block_reg[4][56]  ( .D(block_next[56]), .E(n1127), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFX1 \block_reg[4][55]  ( .D(block_next[55]), .E(n1127), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFX1 \block_reg[4][54]  ( .D(block_next[54]), .E(n1127), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n1127), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n1127), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[4][51]  ( .D(block_next[51]), .E(n1126), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFX1 \block_reg[4][50]  ( .D(block_next[50]), .E(n1126), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n1126), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[4][48]  ( .D(block_next[48]), .E(n1126), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFX1 \block_reg[4][47]  ( .D(block_next[47]), .E(n1126), .CK(clk), .Q(
        \block[4][47] ) );
  EDFFX1 \block_reg[4][46]  ( .D(block_next[46]), .E(n1126), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFX1 \block_reg[4][45]  ( .D(block_next[45]), .E(n1126), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFX1 \block_reg[4][44]  ( .D(block_next[44]), .E(n1126), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFX1 \block_reg[4][43]  ( .D(block_next[43]), .E(n1126), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFX1 \block_reg[4][42]  ( .D(block_next[42]), .E(n1126), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n1126), .CK(clk), .Q(
        \block[4][41] ) );
  EDFFX1 \block_reg[4][40]  ( .D(block_next[40]), .E(n1126), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFX1 \block_reg[4][39]  ( .D(block_next[39]), .E(n1126), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n1125), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n1125), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n1125), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n1125), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFX1 \block_reg[4][34]  ( .D(block_next[34]), .E(n1125), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFX1 \block_reg[4][33]  ( .D(block_next[33]), .E(n1125), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n1125), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[4][31]  ( .D(block_next[31]), .E(n1125), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFX1 \block_reg[4][30]  ( .D(block_next[30]), .E(n1125), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFX1 \block_reg[4][29]  ( .D(block_next[29]), .E(n1125), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFX1 \block_reg[4][28]  ( .D(block_next[28]), .E(n1125), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFX1 \block_reg[4][27]  ( .D(block_next[27]), .E(n1125), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFX1 \block_reg[4][26]  ( .D(block_next[26]), .E(n1125), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFX1 \block_reg[4][25]  ( .D(block_next[25]), .E(n1124), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFX1 \block_reg[4][24]  ( .D(block_next[24]), .E(n1124), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFX1 \block_reg[4][23]  ( .D(block_next[23]), .E(n1124), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFX1 \block_reg[4][22]  ( .D(block_next[22]), .E(n1124), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFX1 \block_reg[4][21]  ( .D(block_next[21]), .E(n1124), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n1124), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFX1 \block_reg[4][19]  ( .D(block_next[19]), .E(n1124), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFX1 \block_reg[4][18]  ( .D(block_next[18]), .E(n1124), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFX1 \block_reg[4][17]  ( .D(block_next[17]), .E(n1124), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFX1 \block_reg[4][16]  ( .D(block_next[16]), .E(n1124), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFX1 \block_reg[4][15]  ( .D(block_next[15]), .E(n1124), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFX1 \block_reg[4][14]  ( .D(block_next[14]), .E(n1124), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFX1 \block_reg[4][13]  ( .D(block_next[13]), .E(n1124), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFX1 \block_reg[4][12]  ( .D(block_next[12]), .E(n1123), .CK(clk), .Q(
        \block[4][12] ) );
  EDFFX1 \block_reg[4][11]  ( .D(block_next[11]), .E(n1123), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFX1 \block_reg[4][10]  ( .D(block_next[10]), .E(n1123), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFX1 \block_reg[4][9]  ( .D(block_next[9]), .E(n1123), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFX1 \block_reg[4][8]  ( .D(block_next[8]), .E(n1123), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFX1 \block_reg[4][7]  ( .D(block_next[7]), .E(n1123), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFX1 \block_reg[4][6]  ( .D(block_next[6]), .E(n1123), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFX1 \block_reg[4][5]  ( .D(block_next[5]), .E(n1123), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFX1 \block_reg[4][4]  ( .D(block_next[4]), .E(n1123), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFX1 \block_reg[4][3]  ( .D(block_next[3]), .E(n1123), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFX1 \block_reg[4][2]  ( .D(block_next[2]), .E(n1123), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFX1 \block_reg[4][1]  ( .D(block_next[1]), .E(n1123), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFX1 \block_reg[4][0]  ( .D(block_next[0]), .E(n1123), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFX1 \block_reg[0][127]  ( .D(block_next[127]), .E(n1158), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFX1 \block_reg[0][126]  ( .D(block_next[126]), .E(n1158), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFX1 \block_reg[0][125]  ( .D(block_next[125]), .E(n1158), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFX1 \block_reg[0][124]  ( .D(block_next[124]), .E(n1162), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFX1 \block_reg[0][123]  ( .D(block_next[123]), .E(n1160), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFX1 \block_reg[0][122]  ( .D(block_next[122]), .E(n1159), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFX1 \block_reg[0][121]  ( .D(block_next[121]), .E(n1161), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFX1 \block_reg[0][120]  ( .D(block_next[120]), .E(n1161), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFX1 \block_reg[0][119]  ( .D(block_next[119]), .E(n1163), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFX1 \block_reg[0][118]  ( .D(block_next[118]), .E(n1164), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFX1 \block_reg[0][117]  ( .D(block_next[117]), .E(n1166), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFX1 \block_reg[0][116]  ( .D(block_next[116]), .E(n1164), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFX1 \block_reg[0][115]  ( .D(block_next[115]), .E(n1166), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFX1 \block_reg[0][114]  ( .D(block_next[114]), .E(n1165), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFX1 \block_reg[0][113]  ( .D(block_next[113]), .E(n1158), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFX1 \block_reg[0][112]  ( .D(block_next[112]), .E(n1158), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFX1 \block_reg[0][111]  ( .D(block_next[111]), .E(n1162), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFX1 \block_reg[0][110]  ( .D(block_next[110]), .E(n1160), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFX1 \block_reg[0][109]  ( .D(block_next[109]), .E(n1159), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFX1 \block_reg[0][108]  ( .D(block_next[108]), .E(n1161), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFX1 \block_reg[0][107]  ( .D(block_next[107]), .E(n1163), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFX1 \block_reg[0][106]  ( .D(block_next[106]), .E(n1163), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFX1 \block_reg[0][105]  ( .D(block_next[105]), .E(n1164), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFX1 \block_reg[0][104]  ( .D(block_next[104]), .E(n1166), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFX1 \block_reg[0][103]  ( .D(block_next[103]), .E(n1165), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFX1 \block_reg[0][102]  ( .D(block_next[102]), .E(n1165), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFX1 \block_reg[0][101]  ( .D(block_next[101]), .E(n1165), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFX1 \block_reg[0][100]  ( .D(block_next[100]), .E(n1165), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFX1 \block_reg[0][99]  ( .D(block_next[99]), .E(n1165), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFX1 \block_reg[0][98]  ( .D(block_next[98]), .E(n1165), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFX1 \block_reg[0][97]  ( .D(block_next[97]), .E(n1165), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFX1 \block_reg[0][96]  ( .D(block_next[96]), .E(n1165), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFX1 \block_reg[0][95]  ( .D(block_next[95]), .E(n1165), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFX1 \block_reg[0][94]  ( .D(block_next[94]), .E(n1165), .CK(clk), .Q(
        \block[0][94] ) );
  EDFFX1 \block_reg[0][93]  ( .D(block_next[93]), .E(n1165), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFX1 \block_reg[0][92]  ( .D(block_next[92]), .E(n1165), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFX1 \block_reg[0][91]  ( .D(block_next[91]), .E(n1165), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFX1 \block_reg[0][90]  ( .D(block_next[90]), .E(n1164), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFX1 \block_reg[0][89]  ( .D(block_next[89]), .E(n1164), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFX1 \block_reg[0][88]  ( .D(block_next[88]), .E(n1164), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFX1 \block_reg[0][87]  ( .D(block_next[87]), .E(n1164), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFX1 \block_reg[0][86]  ( .D(block_next[86]), .E(n1164), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFX1 \block_reg[0][85]  ( .D(block_next[85]), .E(n1164), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFX1 \block_reg[0][84]  ( .D(block_next[84]), .E(n1164), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFX1 \block_reg[0][83]  ( .D(block_next[83]), .E(n1164), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFX1 \block_reg[0][82]  ( .D(block_next[82]), .E(n1164), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFX1 \block_reg[0][81]  ( .D(block_next[81]), .E(n1164), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFX1 \block_reg[0][80]  ( .D(block_next[80]), .E(n1164), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFX1 \block_reg[0][79]  ( .D(block_next[79]), .E(n1164), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFX1 \block_reg[0][78]  ( .D(block_next[78]), .E(n1164), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFX1 \block_reg[0][77]  ( .D(block_next[77]), .E(n1165), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFX1 \block_reg[0][76]  ( .D(block_next[76]), .E(n1162), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFX1 \block_reg[0][75]  ( .D(block_next[75]), .E(n1160), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFX1 \block_reg[0][74]  ( .D(block_next[74]), .E(n1159), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFX1 \block_reg[0][73]  ( .D(block_next[73]), .E(n1161), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFX1 \block_reg[0][72]  ( .D(block_next[72]), .E(n1163), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFX1 \block_reg[0][71]  ( .D(block_next[71]), .E(n1164), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFX1 \block_reg[0][70]  ( .D(block_next[70]), .E(n1166), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFX1 \block_reg[0][69]  ( .D(block_next[69]), .E(n1165), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFX1 \block_reg[0][68]  ( .D(block_next[68]), .E(n1158), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFX1 \block_reg[0][67]  ( .D(block_next[67]), .E(n1162), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFX1 \block_reg[0][66]  ( .D(block_next[66]), .E(n1160), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFX1 \block_reg[0][65]  ( .D(block_next[65]), .E(n1159), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFX1 \block_reg[0][64]  ( .D(block_next[64]), .E(n1163), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[0][63]  ( .D(block_next[63]), .E(n1163), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFX1 \block_reg[0][62]  ( .D(block_next[62]), .E(n1163), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFX1 \block_reg[0][61]  ( .D(block_next[61]), .E(n1163), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFX1 \block_reg[0][60]  ( .D(block_next[60]), .E(n1163), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFX1 \block_reg[0][59]  ( .D(block_next[59]), .E(n1163), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFX1 \block_reg[0][58]  ( .D(block_next[58]), .E(n1163), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFX1 \block_reg[0][57]  ( .D(block_next[57]), .E(n1163), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFX1 \block_reg[0][56]  ( .D(block_next[56]), .E(n1163), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFX1 \block_reg[0][55]  ( .D(block_next[55]), .E(n1163), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFX1 \block_reg[0][54]  ( .D(block_next[54]), .E(n1163), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n1163), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n1163), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[0][51]  ( .D(block_next[51]), .E(n1162), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFX1 \block_reg[0][50]  ( .D(block_next[50]), .E(n1162), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n1162), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[0][48]  ( .D(block_next[48]), .E(n1162), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFX1 \block_reg[0][47]  ( .D(block_next[47]), .E(n1162), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFX1 \block_reg[0][46]  ( .D(block_next[46]), .E(n1162), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFX1 \block_reg[0][45]  ( .D(block_next[45]), .E(n1162), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFX1 \block_reg[0][44]  ( .D(block_next[44]), .E(n1162), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFX1 \block_reg[0][43]  ( .D(block_next[43]), .E(n1162), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFX1 \block_reg[0][42]  ( .D(block_next[42]), .E(n1162), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n1162), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[0][40]  ( .D(block_next[40]), .E(n1162), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFX1 \block_reg[0][39]  ( .D(block_next[39]), .E(n1162), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n1161), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n1161), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n1161), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n1161), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[0][34]  ( .D(block_next[34]), .E(n1161), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFX1 \block_reg[0][33]  ( .D(block_next[33]), .E(n1161), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n1161), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[0][31]  ( .D(block_next[31]), .E(n1161), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFX1 \block_reg[0][30]  ( .D(block_next[30]), .E(n1161), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFX1 \block_reg[0][29]  ( .D(block_next[29]), .E(n1161), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFX1 \block_reg[0][28]  ( .D(block_next[28]), .E(n1161), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFX1 \block_reg[0][27]  ( .D(block_next[27]), .E(n1161), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFX1 \block_reg[0][26]  ( .D(block_next[26]), .E(n1161), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFX1 \block_reg[0][25]  ( .D(block_next[25]), .E(n1160), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFX1 \block_reg[0][24]  ( .D(block_next[24]), .E(n1160), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFX1 \block_reg[0][23]  ( .D(block_next[23]), .E(n1160), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFX1 \block_reg[0][22]  ( .D(block_next[22]), .E(n1160), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFX1 \block_reg[0][21]  ( .D(block_next[21]), .E(n1160), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n1160), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFX1 \block_reg[0][19]  ( .D(block_next[19]), .E(n1160), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFX1 \block_reg[0][18]  ( .D(block_next[18]), .E(n1160), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFX1 \block_reg[0][17]  ( .D(block_next[17]), .E(n1160), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFX1 \block_reg[0][16]  ( .D(block_next[16]), .E(n1160), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFX1 \block_reg[0][15]  ( .D(block_next[15]), .E(n1160), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFX1 \block_reg[0][14]  ( .D(block_next[14]), .E(n1160), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFX1 \block_reg[0][13]  ( .D(block_next[13]), .E(n1160), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFX1 \block_reg[0][12]  ( .D(block_next[12]), .E(n1159), .CK(clk), .Q(
        \block[0][12] ) );
  EDFFX1 \block_reg[0][11]  ( .D(block_next[11]), .E(n1159), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFX1 \block_reg[0][10]  ( .D(block_next[10]), .E(n1159), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFX1 \block_reg[0][9]  ( .D(block_next[9]), .E(n1159), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFX1 \block_reg[0][8]  ( .D(block_next[8]), .E(n1159), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFX1 \block_reg[0][7]  ( .D(block_next[7]), .E(n1159), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFX1 \block_reg[0][6]  ( .D(block_next[6]), .E(n1159), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFX1 \block_reg[0][5]  ( .D(block_next[5]), .E(n1159), .CK(clk), .Q(
        \block[0][5] ) );
  EDFFX1 \block_reg[0][4]  ( .D(block_next[4]), .E(n1159), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFX1 \block_reg[0][3]  ( .D(block_next[3]), .E(n1159), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFX1 \block_reg[0][2]  ( .D(block_next[2]), .E(n1159), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFX1 \block_reg[0][1]  ( .D(block_next[1]), .E(n1159), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFX1 \block_reg[0][0]  ( .D(block_next[0]), .E(n1159), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFX1 \block_reg[6][127]  ( .D(block_next[127]), .E(n1109), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFX1 \block_reg[6][126]  ( .D(block_next[126]), .E(n1110), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFX1 \block_reg[6][125]  ( .D(block_next[125]), .E(n1112), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFX1 \block_reg[6][124]  ( .D(block_next[124]), .E(n1104), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFX1 \block_reg[6][123]  ( .D(block_next[123]), .E(n1106), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFX1 \block_reg[6][122]  ( .D(block_next[122]), .E(n1109), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFX1 \block_reg[6][121]  ( .D(block_next[121]), .E(n1110), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFX1 \block_reg[6][120]  ( .D(block_next[120]), .E(n1112), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFX1 \block_reg[6][119]  ( .D(block_next[119]), .E(n1104), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFX1 \block_reg[6][118]  ( .D(block_next[118]), .E(n1106), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFX1 \block_reg[6][117]  ( .D(block_next[117]), .E(n1109), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFX1 \block_reg[6][116]  ( .D(block_next[116]), .E(n1105), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFX1 \block_reg[6][115]  ( .D(block_next[115]), .E(n1105), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFX1 \block_reg[6][114]  ( .D(block_next[114]), .E(n1105), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFX1 \block_reg[6][113]  ( .D(block_next[113]), .E(n1108), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFX1 \block_reg[6][112]  ( .D(block_next[112]), .E(n1107), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFX1 \block_reg[6][111]  ( .D(block_next[111]), .E(n1111), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFX1 \block_reg[6][110]  ( .D(block_next[110]), .E(n1104), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFX1 \block_reg[6][109]  ( .D(block_next[109]), .E(n1106), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFX1 \block_reg[6][108]  ( .D(block_next[108]), .E(n1109), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFX1 \block_reg[6][107]  ( .D(block_next[107]), .E(n1110), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFX1 \block_reg[6][106]  ( .D(block_next[106]), .E(n1112), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFX1 \block_reg[6][105]  ( .D(block_next[105]), .E(n1104), .CK(clk), .Q(
        \block[6][105] ) );
  EDFFX1 \block_reg[6][104]  ( .D(block_next[104]), .E(n1106), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFX1 \block_reg[6][103]  ( .D(block_next[103]), .E(n1111), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFX1 \block_reg[6][102]  ( .D(block_next[102]), .E(n1111), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFX1 \block_reg[6][101]  ( .D(block_next[101]), .E(n1111), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFX1 \block_reg[6][100]  ( .D(block_next[100]), .E(n1111), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFX1 \block_reg[6][99]  ( .D(block_next[99]), .E(n1111), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFX1 \block_reg[6][98]  ( .D(block_next[98]), .E(n1111), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFX1 \block_reg[6][97]  ( .D(block_next[97]), .E(n1111), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFX1 \block_reg[6][96]  ( .D(block_next[96]), .E(n1111), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFX1 \block_reg[6][95]  ( .D(block_next[95]), .E(n1111), .CK(clk), .Q(
        \block[6][95] ) );
  EDFFX1 \block_reg[6][94]  ( .D(block_next[94]), .E(n1111), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFX1 \block_reg[6][93]  ( .D(block_next[93]), .E(n1111), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFX1 \block_reg[6][92]  ( .D(block_next[92]), .E(n1111), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFX1 \block_reg[6][91]  ( .D(block_next[91]), .E(n1111), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFX1 \block_reg[6][90]  ( .D(block_next[90]), .E(n1110), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFX1 \block_reg[6][89]  ( .D(block_next[89]), .E(n1110), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFX1 \block_reg[6][88]  ( .D(block_next[88]), .E(n1110), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFX1 \block_reg[6][87]  ( .D(block_next[87]), .E(n1110), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFX1 \block_reg[6][86]  ( .D(block_next[86]), .E(n1110), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFX1 \block_reg[6][85]  ( .D(block_next[85]), .E(n1110), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFX1 \block_reg[6][84]  ( .D(block_next[84]), .E(n1110), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFX1 \block_reg[6][83]  ( .D(block_next[83]), .E(n1110), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFX1 \block_reg[6][82]  ( .D(block_next[82]), .E(n1110), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFX1 \block_reg[6][81]  ( .D(block_next[81]), .E(n1110), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFX1 \block_reg[6][80]  ( .D(block_next[80]), .E(n1110), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFX1 \block_reg[6][79]  ( .D(block_next[79]), .E(n1110), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFX1 \block_reg[6][78]  ( .D(block_next[78]), .E(n1110), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFX1 \block_reg[6][77]  ( .D(block_next[77]), .E(n1109), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFX1 \block_reg[6][76]  ( .D(block_next[76]), .E(n1109), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFX1 \block_reg[6][75]  ( .D(block_next[75]), .E(n1109), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFX1 \block_reg[6][74]  ( .D(block_next[74]), .E(n1109), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFX1 \block_reg[6][73]  ( .D(block_next[73]), .E(n1109), .CK(clk), .Q(
        \block[6][73] ) );
  EDFFX1 \block_reg[6][72]  ( .D(block_next[72]), .E(n1109), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFX1 \block_reg[6][71]  ( .D(block_next[71]), .E(n1109), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFX1 \block_reg[6][70]  ( .D(block_next[70]), .E(n1109), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFX1 \block_reg[6][69]  ( .D(block_next[69]), .E(n1109), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFX1 \block_reg[6][68]  ( .D(block_next[68]), .E(n1109), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFX1 \block_reg[6][67]  ( .D(block_next[67]), .E(n1109), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFX1 \block_reg[6][66]  ( .D(block_next[66]), .E(n1109), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFX1 \block_reg[6][65]  ( .D(block_next[65]), .E(n1109), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFX1 \block_reg[6][64]  ( .D(block_next[64]), .E(n1108), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFX1 \block_reg[6][63]  ( .D(block_next[63]), .E(n1108), .CK(clk), .Q(
        \block[6][63] ) );
  EDFFX1 \block_reg[6][62]  ( .D(block_next[62]), .E(n1108), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFX1 \block_reg[6][61]  ( .D(block_next[61]), .E(n1108), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFX1 \block_reg[6][60]  ( .D(block_next[60]), .E(n1108), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFX1 \block_reg[6][59]  ( .D(block_next[59]), .E(n1108), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFX1 \block_reg[6][58]  ( .D(block_next[58]), .E(n1108), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFX1 \block_reg[6][57]  ( .D(block_next[57]), .E(n1108), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFX1 \block_reg[6][56]  ( .D(block_next[56]), .E(n1108), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFX1 \block_reg[6][55]  ( .D(block_next[55]), .E(n1108), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFX1 \block_reg[6][54]  ( .D(block_next[54]), .E(n1108), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n1108), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n1108), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[6][51]  ( .D(block_next[51]), .E(n1107), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFX1 \block_reg[6][50]  ( .D(block_next[50]), .E(n1107), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFX1 \block_reg[6][49]  ( .D(block_next[49]), .E(n1107), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFX1 \block_reg[6][48]  ( .D(block_next[48]), .E(n1107), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFX1 \block_reg[6][47]  ( .D(block_next[47]), .E(n1107), .CK(clk), .Q(
        \block[6][47] ) );
  EDFFX1 \block_reg[6][46]  ( .D(block_next[46]), .E(n1107), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFX1 \block_reg[6][45]  ( .D(block_next[45]), .E(n1107), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFX1 \block_reg[6][44]  ( .D(block_next[44]), .E(n1107), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFX1 \block_reg[6][43]  ( .D(block_next[43]), .E(n1107), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFX1 \block_reg[6][42]  ( .D(block_next[42]), .E(n1107), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n1107), .CK(clk), .Q(
        \block[6][41] ) );
  EDFFX1 \block_reg[6][40]  ( .D(block_next[40]), .E(n1107), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFX1 \block_reg[6][39]  ( .D(block_next[39]), .E(n1107), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n1106), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n1106), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n1106), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n1106), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFX1 \block_reg[6][34]  ( .D(block_next[34]), .E(n1106), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFX1 \block_reg[6][33]  ( .D(block_next[33]), .E(n1106), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n1106), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[6][31]  ( .D(block_next[31]), .E(n1106), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFX1 \block_reg[6][30]  ( .D(block_next[30]), .E(n1106), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFX1 \block_reg[6][29]  ( .D(block_next[29]), .E(n1106), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFX1 \block_reg[6][28]  ( .D(block_next[28]), .E(n1106), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFX1 \block_reg[6][27]  ( .D(block_next[27]), .E(n1106), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFX1 \block_reg[6][26]  ( .D(block_next[26]), .E(n1106), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFX1 \block_reg[6][25]  ( .D(block_next[25]), .E(n1105), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFX1 \block_reg[6][24]  ( .D(block_next[24]), .E(n1105), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFX1 \block_reg[6][23]  ( .D(block_next[23]), .E(n1105), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFX1 \block_reg[6][22]  ( .D(block_next[22]), .E(n1105), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFX1 \block_reg[6][21]  ( .D(block_next[21]), .E(n1105), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n1105), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFX1 \block_reg[6][19]  ( .D(block_next[19]), .E(n1105), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFX1 \block_reg[6][18]  ( .D(block_next[18]), .E(n1105), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFX1 \block_reg[6][17]  ( .D(block_next[17]), .E(n1105), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFX1 \block_reg[6][16]  ( .D(block_next[16]), .E(n1105), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFX1 \block_reg[6][15]  ( .D(block_next[15]), .E(n1105), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFX1 \block_reg[6][14]  ( .D(block_next[14]), .E(n1105), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFX1 \block_reg[6][13]  ( .D(block_next[13]), .E(n1105), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFX1 \block_reg[6][12]  ( .D(block_next[12]), .E(n1104), .CK(clk), .Q(
        \block[6][12] ) );
  EDFFX1 \block_reg[6][11]  ( .D(block_next[11]), .E(n1104), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFX1 \block_reg[6][10]  ( .D(block_next[10]), .E(n1104), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFX1 \block_reg[6][9]  ( .D(block_next[9]), .E(n1104), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFX1 \block_reg[6][8]  ( .D(block_next[8]), .E(n1104), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFX1 \block_reg[6][7]  ( .D(block_next[7]), .E(n1104), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFX1 \block_reg[6][6]  ( .D(block_next[6]), .E(n1104), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFX1 \block_reg[6][5]  ( .D(block_next[5]), .E(n1104), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFX1 \block_reg[6][4]  ( .D(block_next[4]), .E(n1104), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFX1 \block_reg[6][3]  ( .D(block_next[3]), .E(n1104), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFX1 \block_reg[6][2]  ( .D(block_next[2]), .E(n1104), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFX1 \block_reg[6][1]  ( .D(block_next[1]), .E(n1104), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFX1 \block_reg[6][0]  ( .D(block_next[0]), .E(n1104), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFX1 \block_reg[2][127]  ( .D(block_next[127]), .E(n1140), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFX1 \block_reg[2][126]  ( .D(block_next[126]), .E(n1140), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFX1 \block_reg[2][125]  ( .D(block_next[125]), .E(n1140), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFX1 \block_reg[2][124]  ( .D(block_next[124]), .E(n1144), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFX1 \block_reg[2][123]  ( .D(block_next[123]), .E(n1142), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFX1 \block_reg[2][122]  ( .D(block_next[122]), .E(n1141), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFX1 \block_reg[2][121]  ( .D(block_next[121]), .E(n1143), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFX1 \block_reg[2][120]  ( .D(block_next[120]), .E(n1143), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFX1 \block_reg[2][119]  ( .D(block_next[119]), .E(n1145), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFX1 \block_reg[2][118]  ( .D(block_next[118]), .E(n1146), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFX1 \block_reg[2][117]  ( .D(block_next[117]), .E(n1148), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFX1 \block_reg[2][116]  ( .D(block_next[116]), .E(n1146), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFX1 \block_reg[2][115]  ( .D(block_next[115]), .E(n1148), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFX1 \block_reg[2][114]  ( .D(block_next[114]), .E(n1147), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFX1 \block_reg[2][113]  ( .D(block_next[113]), .E(n1140), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFX1 \block_reg[2][112]  ( .D(block_next[112]), .E(n1140), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFX1 \block_reg[2][111]  ( .D(block_next[111]), .E(n1144), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFX1 \block_reg[2][110]  ( .D(block_next[110]), .E(n1142), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFX1 \block_reg[2][109]  ( .D(block_next[109]), .E(n1141), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFX1 \block_reg[2][108]  ( .D(block_next[108]), .E(n1143), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFX1 \block_reg[2][107]  ( .D(block_next[107]), .E(n1145), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFX1 \block_reg[2][106]  ( .D(block_next[106]), .E(n1145), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFX1 \block_reg[2][105]  ( .D(block_next[105]), .E(n1146), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFX1 \block_reg[2][104]  ( .D(block_next[104]), .E(n1148), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFX1 \block_reg[2][103]  ( .D(block_next[103]), .E(n1147), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFX1 \block_reg[2][102]  ( .D(block_next[102]), .E(n1147), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFX1 \block_reg[2][101]  ( .D(block_next[101]), .E(n1147), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFX1 \block_reg[2][100]  ( .D(block_next[100]), .E(n1147), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFX1 \block_reg[2][99]  ( .D(block_next[99]), .E(n1147), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFX1 \block_reg[2][98]  ( .D(block_next[98]), .E(n1147), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFX1 \block_reg[2][97]  ( .D(block_next[97]), .E(n1147), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFX1 \block_reg[2][96]  ( .D(block_next[96]), .E(n1147), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFX1 \block_reg[2][95]  ( .D(block_next[95]), .E(n1147), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFX1 \block_reg[2][94]  ( .D(block_next[94]), .E(n1147), .CK(clk), .Q(
        \block[2][94] ) );
  EDFFX1 \block_reg[2][93]  ( .D(block_next[93]), .E(n1147), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFX1 \block_reg[2][92]  ( .D(block_next[92]), .E(n1147), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFX1 \block_reg[2][91]  ( .D(block_next[91]), .E(n1147), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFX1 \block_reg[2][90]  ( .D(block_next[90]), .E(n1146), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFX1 \block_reg[2][89]  ( .D(block_next[89]), .E(n1146), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFX1 \block_reg[2][88]  ( .D(block_next[88]), .E(n1146), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFX1 \block_reg[2][87]  ( .D(block_next[87]), .E(n1146), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFX1 \block_reg[2][86]  ( .D(block_next[86]), .E(n1146), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFX1 \block_reg[2][85]  ( .D(block_next[85]), .E(n1146), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFX1 \block_reg[2][84]  ( .D(block_next[84]), .E(n1146), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFX1 \block_reg[2][83]  ( .D(block_next[83]), .E(n1146), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFX1 \block_reg[2][82]  ( .D(block_next[82]), .E(n1146), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFX1 \block_reg[2][81]  ( .D(block_next[81]), .E(n1146), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFX1 \block_reg[2][80]  ( .D(block_next[80]), .E(n1146), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFX1 \block_reg[2][79]  ( .D(block_next[79]), .E(n1146), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFX1 \block_reg[2][78]  ( .D(block_next[78]), .E(n1146), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFX1 \block_reg[2][77]  ( .D(block_next[77]), .E(n1147), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFX1 \block_reg[2][76]  ( .D(block_next[76]), .E(n1144), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFX1 \block_reg[2][75]  ( .D(block_next[75]), .E(n1142), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFX1 \block_reg[2][74]  ( .D(block_next[74]), .E(n1141), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFX1 \block_reg[2][73]  ( .D(block_next[73]), .E(n1143), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFX1 \block_reg[2][72]  ( .D(block_next[72]), .E(n1145), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFX1 \block_reg[2][71]  ( .D(block_next[71]), .E(n1146), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFX1 \block_reg[2][70]  ( .D(block_next[70]), .E(n1148), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFX1 \block_reg[2][69]  ( .D(block_next[69]), .E(n1147), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFX1 \block_reg[2][68]  ( .D(block_next[68]), .E(n1140), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFX1 \block_reg[2][67]  ( .D(block_next[67]), .E(n1144), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFX1 \block_reg[2][66]  ( .D(block_next[66]), .E(n1142), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFX1 \block_reg[2][65]  ( .D(block_next[65]), .E(n1141), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFX1 \block_reg[2][64]  ( .D(block_next[64]), .E(n1145), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFX1 \block_reg[2][63]  ( .D(block_next[63]), .E(n1145), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFX1 \block_reg[2][62]  ( .D(block_next[62]), .E(n1145), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFX1 \block_reg[2][61]  ( .D(block_next[61]), .E(n1145), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFX1 \block_reg[2][60]  ( .D(block_next[60]), .E(n1145), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFX1 \block_reg[2][59]  ( .D(block_next[59]), .E(n1145), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFX1 \block_reg[2][58]  ( .D(block_next[58]), .E(n1145), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFX1 \block_reg[2][57]  ( .D(block_next[57]), .E(n1145), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFX1 \block_reg[2][56]  ( .D(block_next[56]), .E(n1145), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFX1 \block_reg[2][55]  ( .D(block_next[55]), .E(n1145), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFX1 \block_reg[2][54]  ( .D(block_next[54]), .E(n1145), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFX1 \block_reg[2][53]  ( .D(block_next[53]), .E(n1145), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFX1 \block_reg[2][52]  ( .D(block_next[52]), .E(n1145), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFX1 \block_reg[2][51]  ( .D(block_next[51]), .E(n1144), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFX1 \block_reg[2][50]  ( .D(block_next[50]), .E(n1144), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFX1 \block_reg[2][49]  ( .D(block_next[49]), .E(n1144), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFX1 \block_reg[2][48]  ( .D(block_next[48]), .E(n1144), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFX1 \block_reg[2][47]  ( .D(block_next[47]), .E(n1144), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFX1 \block_reg[2][46]  ( .D(block_next[46]), .E(n1144), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFX1 \block_reg[2][45]  ( .D(block_next[45]), .E(n1144), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFX1 \block_reg[2][44]  ( .D(block_next[44]), .E(n1144), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFX1 \block_reg[2][43]  ( .D(block_next[43]), .E(n1144), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFX1 \block_reg[2][42]  ( .D(block_next[42]), .E(n1144), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFX1 \block_reg[2][41]  ( .D(block_next[41]), .E(n1144), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFX1 \block_reg[2][40]  ( .D(block_next[40]), .E(n1144), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFX1 \block_reg[2][39]  ( .D(block_next[39]), .E(n1144), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFX1 \block_reg[2][38]  ( .D(block_next[38]), .E(n1143), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFX1 \block_reg[2][37]  ( .D(block_next[37]), .E(n1143), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFX1 \block_reg[2][36]  ( .D(block_next[36]), .E(n1143), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFX1 \block_reg[2][35]  ( .D(block_next[35]), .E(n1143), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFX1 \block_reg[2][34]  ( .D(block_next[34]), .E(n1143), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFX1 \block_reg[2][33]  ( .D(block_next[33]), .E(n1143), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFX1 \block_reg[2][32]  ( .D(block_next[32]), .E(n1143), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFX1 \block_reg[2][31]  ( .D(block_next[31]), .E(n1143), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFX1 \block_reg[2][30]  ( .D(block_next[30]), .E(n1143), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFX1 \block_reg[2][29]  ( .D(block_next[29]), .E(n1143), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFX1 \block_reg[2][28]  ( .D(block_next[28]), .E(n1143), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFX1 \block_reg[2][27]  ( .D(block_next[27]), .E(n1143), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFX1 \block_reg[2][26]  ( .D(block_next[26]), .E(n1143), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFX1 \block_reg[2][25]  ( .D(block_next[25]), .E(n1142), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFX1 \block_reg[2][24]  ( .D(block_next[24]), .E(n1142), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFX1 \block_reg[2][23]  ( .D(block_next[23]), .E(n1142), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFX1 \block_reg[2][22]  ( .D(block_next[22]), .E(n1142), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFX1 \block_reg[2][21]  ( .D(block_next[21]), .E(n1142), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFX1 \block_reg[2][20]  ( .D(block_next[20]), .E(n1142), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFX1 \block_reg[2][19]  ( .D(block_next[19]), .E(n1142), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFX1 \block_reg[2][18]  ( .D(block_next[18]), .E(n1142), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFX1 \block_reg[2][17]  ( .D(block_next[17]), .E(n1142), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFX1 \block_reg[2][16]  ( .D(block_next[16]), .E(n1142), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFX1 \block_reg[2][15]  ( .D(block_next[15]), .E(n1142), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFX1 \block_reg[2][14]  ( .D(block_next[14]), .E(n1142), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFX1 \block_reg[2][13]  ( .D(block_next[13]), .E(n1142), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFX1 \block_reg[2][12]  ( .D(block_next[12]), .E(n1141), .CK(clk), .Q(
        \block[2][12] ) );
  EDFFX1 \block_reg[2][11]  ( .D(block_next[11]), .E(n1141), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFX1 \block_reg[2][10]  ( .D(block_next[10]), .E(n1141), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFX1 \block_reg[2][9]  ( .D(block_next[9]), .E(n1141), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFX1 \block_reg[2][8]  ( .D(block_next[8]), .E(n1141), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFX1 \block_reg[2][7]  ( .D(block_next[7]), .E(n1141), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFX1 \block_reg[2][6]  ( .D(block_next[6]), .E(n1141), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFX1 \block_reg[2][5]  ( .D(block_next[5]), .E(n1141), .CK(clk), .Q(
        \block[2][5] ) );
  EDFFX1 \block_reg[2][4]  ( .D(block_next[4]), .E(n1141), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFX1 \block_reg[2][3]  ( .D(block_next[3]), .E(n1141), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFX1 \block_reg[2][2]  ( .D(block_next[2]), .E(n1141), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFX1 \block_reg[2][1]  ( .D(block_next[1]), .E(n1141), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFX1 \block_reg[2][0]  ( .D(block_next[0]), .E(n1141), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n1095), .CK(clk), 
        .Q(\blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(blocktag_next[23]), .E(N1777), .CK(clk), 
        .QN(n646) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n1095), .CK(clk), 
        .Q(\blocktag[7][22] ) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n1095), .CK(clk), 
        .QN(n634) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n1095), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n1095), .CK(clk), 
        .QN(n626) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n1095), .CK(clk), 
        .Q(\blocktag[7][18] ) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(blocktag_next[17]), .E(N1777), .CK(clk), 
        .Q(\blocktag[7][17] ) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(N1777), .CK(clk), 
        .Q(\blocktag[7][16] ) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(N1777), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(blocktag_next[14]), .E(n1103), .CK(clk), 
        .Q(\blocktag[7][14] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n1103), .CK(clk), 
        .Q(\blocktag[7][13] ) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(blocktag_next[12]), .E(n1103), .CK(clk), 
        .Q(\blocktag[7][12] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n1103), .CK(clk), 
        .Q(\blocktag[7][11] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(blocktag_next[10]), .E(n1103), .CK(clk), 
        .Q(\blocktag[7][10] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(blocktag_next[7]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][7] ) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][6] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(blocktag_next[5]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][4] ) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n1103), .CK(clk), .Q(
        \blocktag[7][2] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n1102), .CK(clk), .Q(
        \blocktag[7][1] ) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n1102), .CK(clk), 
        .QN(n649) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n1131), .CK(clk), 
        .QN(n622) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(blocktag_next[23]), .E(n1131), .CK(clk), 
        .QN(n642) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n1131), .CK(clk), 
        .QN(n638) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n1131), .CK(clk), 
        .QN(n630) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n1131), .CK(clk), 
        .Q(\blocktag[3][20] ) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n1131), .CK(clk), 
        .Q(\blocktag[3][19] ) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(N1772), .CK(clk), 
        .Q(\blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(blocktag_next[17]), .E(N1772), .CK(clk), 
        .Q(\blocktag[3][17] ) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(N1772), .CK(clk), 
        .Q(\blocktag[3][16] ) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(N1772), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(blocktag_next[14]), .E(n1139), .CK(clk), 
        .Q(\blocktag[3][14] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n1139), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(blocktag_next[12]), .E(n1139), .CK(clk), 
        .Q(\blocktag[3][12] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n1139), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(blocktag_next[10]), .E(n1139), .CK(clk), 
        .Q(\blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][9] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][8] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(blocktag_next[7]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][7] ) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][6] ) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(blocktag_next[5]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][4] ) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n1139), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n1138), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n1138), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n1113), .CK(clk), 
        .Q(\blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(blocktag_next[23]), .E(N1774), .CK(clk), 
        .QN(n644) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n1113), .CK(clk), 
        .Q(\blocktag[5][22] ) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n1113), .CK(clk), 
        .QN(n632) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n1113), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n1113), .CK(clk), 
        .QN(n624) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n1113), .CK(clk), 
        .Q(\blocktag[5][18] ) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(blocktag_next[17]), .E(N1774), .CK(clk), 
        .Q(\blocktag[5][17] ) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(N1774), .CK(clk), 
        .Q(\blocktag[5][16] ) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(N1774), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(blocktag_next[14]), .E(n1121), .CK(clk), 
        .Q(\blocktag[5][14] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n1121), .CK(clk), 
        .Q(\blocktag[5][13] ) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(blocktag_next[12]), .E(n1121), .CK(clk), 
        .Q(\blocktag[5][12] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n1121), .CK(clk), 
        .Q(\blocktag[5][11] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(blocktag_next[10]), .E(n1121), .CK(clk), 
        .Q(\blocktag[5][10] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(blocktag_next[7]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][7] ) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][6] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(blocktag_next[5]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][4] ) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n1121), .CK(clk), .Q(
        \blocktag[5][2] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n1120), .CK(clk), .Q(
        \blocktag[5][1] ) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n1157), .CK(clk), 
        .QN(n620) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(blocktag_next[23]), .E(n1157), .CK(clk), 
        .QN(n640) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n1157), .CK(clk), 
        .QN(n636) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n1157), .CK(clk), 
        .QN(n628) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][20] ) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][19] ) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(blocktag_next[17]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][17] ) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][16] ) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n1157), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(blocktag_next[14]), .E(n1156), .CK(clk), 
        .Q(\blocktag[1][14] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n1156), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(blocktag_next[12]), .E(n1156), .CK(clk), 
        .Q(\blocktag[1][12] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n1156), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(blocktag_next[10]), .E(n1156), .CK(clk), 
        .Q(\blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][8] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(blocktag_next[7]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][7] ) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][6] ) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(blocktag_next[5]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][4] ) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n1154), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n1156), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n1122), .CK(clk), 
        .Q(\blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(blocktag_next[23]), .E(n1122), .CK(clk), 
        .QN(n643) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n1122), .CK(clk), 
        .Q(\blocktag[4][22] ) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n1122), .CK(clk), 
        .QN(n631) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n1122), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n1122), .CK(clk), 
        .QN(n623) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(N1773), .CK(clk), 
        .Q(\blocktag[4][18] ) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(blocktag_next[17]), .E(N1773), .CK(clk), 
        .Q(\blocktag[4][17] ) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(N1773), .CK(clk), 
        .Q(\blocktag[4][16] ) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(N1773), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(blocktag_next[14]), .E(n1130), .CK(clk), 
        .Q(\blocktag[4][14] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n1130), .CK(clk), 
        .Q(\blocktag[4][13] ) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(blocktag_next[12]), .E(n1130), .CK(clk), 
        .Q(\blocktag[4][12] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n1130), .CK(clk), 
        .Q(\blocktag[4][11] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(blocktag_next[10]), .E(n1130), .CK(clk), 
        .Q(\blocktag[4][10] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(blocktag_next[7]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][7] ) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][6] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(blocktag_next[5]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][4] ) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n1130), .CK(clk), .Q(
        \blocktag[4][2] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n1129), .CK(clk), .Q(
        \blocktag[4][1] ) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n1129), .CK(clk), 
        .QN(n647) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n1158), .CK(clk), 
        .QN(n619) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(blocktag_next[23]), .E(n1158), .CK(clk), 
        .QN(n639) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n1158), .CK(clk), 
        .QN(n635) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n1158), .CK(clk), 
        .QN(n627) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n1158), .CK(clk), 
        .Q(\blocktag[0][20] ) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n1158), .CK(clk), 
        .Q(\blocktag[0][19] ) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(N1768), .CK(clk), 
        .Q(\blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(blocktag_next[17]), .E(N1768), .CK(clk), 
        .Q(\blocktag[0][17] ) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(N1768), .CK(clk), 
        .Q(\blocktag[0][16] ) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(N1768), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(blocktag_next[14]), .E(n1166), .CK(clk), 
        .Q(\blocktag[0][14] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n1166), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(blocktag_next[12]), .E(n1166), .CK(clk), 
        .Q(\blocktag[0][12] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n1166), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(blocktag_next[10]), .E(n1166), .CK(clk), 
        .Q(\blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][8] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(blocktag_next[7]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][7] ) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][6] ) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(blocktag_next[5]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][4] ) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n1166), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n1165), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n1165), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(blocktag_next[23]), .E(n1109), .CK(clk), 
        .QN(n645) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n1110), .CK(clk), 
        .Q(\blocktag[6][22] ) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n1106), .CK(clk), 
        .QN(n633) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n1109), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n1104), .CK(clk), 
        .QN(n625) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n1106), .CK(clk), 
        .Q(\blocktag[6][18] ) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(blocktag_next[17]), .E(n1104), .CK(clk), 
        .Q(\blocktag[6][17] ) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][16] ) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n1110), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(blocktag_next[14]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][14] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][13] ) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(blocktag_next[12]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][12] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][11] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(blocktag_next[10]), .E(n1112), .CK(clk), 
        .Q(\blocktag[6][10] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(blocktag_next[7]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][7] ) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][6] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(blocktag_next[5]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][4] ) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][2] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n1112), .CK(clk), .Q(
        \blocktag[6][1] ) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n1110), .CK(clk), 
        .QN(n648) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n1140), .CK(clk), 
        .QN(n621) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(blocktag_next[23]), .E(n1140), .CK(clk), 
        .QN(n641) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n1140), .CK(clk), 
        .QN(n637) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n1140), .CK(clk), 
        .QN(n629) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n1140), .CK(clk), 
        .Q(\blocktag[2][20] ) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n1140), .CK(clk), 
        .Q(\blocktag[2][19] ) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(N1771), .CK(clk), 
        .Q(\blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(blocktag_next[17]), .E(N1771), .CK(clk), 
        .Q(\blocktag[2][17] ) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(N1771), .CK(clk), 
        .Q(\blocktag[2][16] ) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(N1771), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(blocktag_next[14]), .E(n1148), .CK(clk), 
        .Q(\blocktag[2][14] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n1148), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(blocktag_next[12]), .E(n1148), .CK(clk), 
        .Q(\blocktag[2][12] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n1148), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(blocktag_next[10]), .E(n1148), .CK(clk), 
        .Q(\blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][8] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(blocktag_next[7]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][7] ) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][6] ) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(blocktag_next[5]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][4] ) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n1148), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n1147), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n1147), .CK(clk), .Q(
        \blocktag[2][0] ) );
  DFFRX1 \blockvalid_reg[7]  ( .D(n503), .CK(clk), .RN(n1173), .Q(
        blockvalid[7]), .QN(n486) );
  DFFRX1 \blockvalid_reg[3]  ( .D(n498), .CK(clk), .RN(n1173), .Q(
        blockvalid[3]), .QN(n482) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n494), .CK(clk), .RN(n1173), .Q(
        blockdirty[7]), .QN(n478) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n490), .CK(clk), .RN(n1173), .Q(
        blockdirty[3]), .QN(n474) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n500), .CK(clk), .RN(n1173), .Q(
        blockvalid[5]), .QN(n484) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n496), .CK(clk), .RN(n1173), .Q(
        blockvalid[1]), .QN(n480) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n492), .CK(clk), .RN(n1173), .Q(
        blockdirty[5]), .QN(n476) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n488), .CK(clk), .RN(n1173), .Q(
        blockdirty[1]), .QN(n472) );
  DFFRX1 \blockvalid_reg[4]  ( .D(n499), .CK(clk), .RN(n1173), .Q(
        blockvalid[4]), .QN(n483) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n495), .CK(clk), .RN(n1173), .Q(
        blockvalid[0]), .QN(n479) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n491), .CK(clk), .RN(n1173), .Q(
        blockdirty[4]), .QN(n475) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n487), .CK(clk), .RN(n1173), .Q(
        blockdirty[0]), .QN(n471) );
  DFFRX1 \blockvalid_reg[6]  ( .D(n501), .CK(clk), .RN(n1173), .Q(
        blockvalid[6]), .QN(n485) );
  DFFRX1 \blockvalid_reg[2]  ( .D(n497), .CK(clk), .RN(n1173), .Q(
        blockvalid[2]), .QN(n481) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n493), .CK(clk), .RN(n1173), .Q(
        blockdirty[6]), .QN(n477) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n489), .CK(clk), .RN(n1173), .Q(
        blockdirty[2]), .QN(n473) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(n1120), .CK(clk), 
        .QN(n1172) );
  CLKBUFX2 U839 ( .A(n1029), .Y(n1031) );
  CLKBUFX2 U840 ( .A(n1029), .Y(n1030) );
  BUFX4 U841 ( .A(n267), .Y(n504) );
  CLKBUFX8 U842 ( .A(n277), .Y(n505) );
  NAND3XL U843 ( .A(proc_addr[1]), .B(n1258), .C(n164), .Y(n277) );
  NOR2X8 U844 ( .A(n145), .B(n611), .Y(n164) );
  INVX8 U845 ( .A(n1047), .Y(n506) );
  INVXL U846 ( .A(n1176), .Y(mem_write) );
  INVX4 U847 ( .A(n1419), .Y(n1176) );
  CLKBUFX6 U848 ( .A(n1053), .Y(n1049) );
  CLKBUFX6 U849 ( .A(n1053), .Y(n1052) );
  BUFX8 U850 ( .A(n1051), .Y(n1047) );
  BUFX8 U851 ( .A(n1050), .Y(n1045) );
  BUFX8 U852 ( .A(n1046), .Y(n1048) );
  NOR3X4 U853 ( .A(n1174), .B(proc_write), .C(n145), .Y(n143) );
  NAND2X2 U854 ( .A(valid), .B(n256), .Y(n145) );
  CLKBUFX3 U855 ( .A(n263), .Y(n508) );
  CLKBUFX3 U856 ( .A(n263), .Y(n1069) );
  AND4X4 U857 ( .A(n434), .B(n435), .C(n436), .D(n437), .Y(n256) );
  CLKINVX1 U858 ( .A(n1170), .Y(n1169) );
  NOR3X1 U859 ( .A(n446), .B(n555), .C(n449), .Y(n436) );
  AND4X1 U860 ( .A(n340), .B(n505), .C(n263), .D(n1175), .Y(n342) );
  AND4X1 U861 ( .A(n340), .B(n341), .C(n263), .D(n1175), .Y(n276) );
  INVX6 U862 ( .A(N32), .Y(n1170) );
  CLKINVX1 U863 ( .A(N33), .Y(n1168) );
  AND4X1 U864 ( .A(n340), .B(n505), .C(n341), .D(n1175), .Y(n262) );
  NOR2BX1 U865 ( .AN(n505), .B(n431), .Y(n430) );
  AND3X2 U866 ( .A(n255), .B(n612), .C(n165), .Y(mem_read) );
  NAND3X1 U867 ( .A(n433), .B(n1175), .C(n613), .Y(n260) );
  CLKMX2X2 U868 ( .A(n806), .B(n807), .S0(n1035), .Y(n510) );
  CLKMX2X2 U869 ( .A(n804), .B(n805), .S0(n1038), .Y(n511) );
  CLKMX2X2 U870 ( .A(n802), .B(n803), .S0(n1040), .Y(n512) );
  CLKMX2X2 U871 ( .A(n800), .B(n801), .S0(n1036), .Y(n513) );
  CLKMX2X2 U872 ( .A(n798), .B(n799), .S0(n1035), .Y(n514) );
  CLKMX2X2 U873 ( .A(n796), .B(n797), .S0(n1039), .Y(n515) );
  CLKMX2X2 U874 ( .A(n794), .B(n795), .S0(n1039), .Y(n516) );
  CLKMX2X2 U875 ( .A(n792), .B(n793), .S0(n1039), .Y(n517) );
  CLKMX2X2 U876 ( .A(n790), .B(n791), .S0(n1039), .Y(n518) );
  CLKMX2X2 U877 ( .A(n788), .B(n789), .S0(n1039), .Y(n519) );
  CLKMX2X2 U878 ( .A(n786), .B(n787), .S0(n1039), .Y(n520) );
  CLKMX2X2 U879 ( .A(n784), .B(n785), .S0(n1039), .Y(n521) );
  CLKMX2X2 U880 ( .A(n782), .B(n783), .S0(n1039), .Y(n522) );
  CLKMX2X2 U881 ( .A(n780), .B(n781), .S0(n1039), .Y(n523) );
  CLKMX2X2 U882 ( .A(n778), .B(n779), .S0(n1039), .Y(n524) );
  CLKMX2X2 U883 ( .A(n776), .B(n777), .S0(n1039), .Y(n525) );
  CLKMX2X2 U884 ( .A(n774), .B(n775), .S0(n1039), .Y(n526) );
  CLKMX2X2 U885 ( .A(n772), .B(n773), .S0(n1038), .Y(n527) );
  CLKMX2X2 U886 ( .A(n770), .B(n771), .S0(n1038), .Y(n528) );
  CLKMX2X2 U887 ( .A(n768), .B(n769), .S0(n1038), .Y(n529) );
  CLKMX2X2 U888 ( .A(n766), .B(n767), .S0(n1038), .Y(n530) );
  CLKMX2X2 U889 ( .A(n764), .B(n765), .S0(n1038), .Y(n531) );
  CLKMX2X2 U890 ( .A(n762), .B(n763), .S0(n1038), .Y(n532) );
  CLKMX2X2 U891 ( .A(n760), .B(n761), .S0(n1038), .Y(n533) );
  CLKMX2X2 U892 ( .A(n758), .B(n759), .S0(n1038), .Y(n534) );
  CLKMX2X2 U893 ( .A(n756), .B(n757), .S0(n1038), .Y(n535) );
  CLKMX2X2 U894 ( .A(n754), .B(n755), .S0(n1038), .Y(n536) );
  CLKMX2X2 U895 ( .A(n752), .B(n753), .S0(n1038), .Y(n537) );
  CLKMX2X2 U896 ( .A(n750), .B(n751), .S0(n1038), .Y(n538) );
  CLKMX2X2 U897 ( .A(n748), .B(n749), .S0(n1037), .Y(n539) );
  CLKMX2X2 U898 ( .A(n746), .B(n747), .S0(n1037), .Y(n540) );
  CLKMX2X2 U899 ( .A(n744), .B(n745), .S0(n1037), .Y(n541) );
  CLKMX2X2 U900 ( .A(n954), .B(n955), .S0(n1044), .Y(n542) );
  CLKMX2X2 U901 ( .A(n964), .B(n965), .S0(n1044), .Y(n543) );
  CLKMX2X2 U902 ( .A(n958), .B(n959), .S0(n1044), .Y(n544) );
  CLKMX2X2 U903 ( .A(n956), .B(n957), .S0(n1044), .Y(n545) );
  CLKMX2X2 U904 ( .A(n936), .B(n937), .S0(n1043), .Y(n546) );
  CLKMX2X2 U905 ( .A(n934), .B(n935), .S0(n1043), .Y(n547) );
  CLKMX2X2 U906 ( .A(n932), .B(n933), .S0(n1043), .Y(n548) );
  CLKMX2X2 U907 ( .A(n930), .B(n931), .S0(n1043), .Y(n549) );
  CLKMX2X2 U908 ( .A(n920), .B(n921), .S0(n1042), .Y(n550) );
  CLKMX2X2 U909 ( .A(n922), .B(n923), .S0(n1043), .Y(n551) );
  CLKMX2X2 U910 ( .A(n944), .B(n945), .S0(n1043), .Y(n552) );
  CLKMX2X2 U911 ( .A(n924), .B(n925), .S0(n1043), .Y(n553) );
  AND2X2 U912 ( .A(n617), .B(n618), .Y(n554) );
  OR2X1 U913 ( .A(n448), .B(n447), .Y(n555) );
  CLKMX2X2 U914 ( .A(n870), .B(n871), .S0(n1037), .Y(n556) );
  CLKMX2X2 U915 ( .A(n868), .B(n869), .S0(n1039), .Y(n557) );
  CLKMX2X2 U916 ( .A(n866), .B(n867), .S0(n1035), .Y(n558) );
  CLKMX2X2 U917 ( .A(n864), .B(n865), .S0(n1038), .Y(n559) );
  CLKMX2X2 U918 ( .A(n862), .B(n863), .S0(n1040), .Y(n560) );
  CLKMX2X2 U919 ( .A(n860), .B(n861), .S0(n1036), .Y(n561) );
  CLKMX2X2 U920 ( .A(n858), .B(n859), .S0(n1041), .Y(n562) );
  CLKMX2X2 U921 ( .A(n856), .B(n857), .S0(n1041), .Y(n563) );
  CLKMX2X2 U922 ( .A(n854), .B(n855), .S0(n1037), .Y(n564) );
  CLKMX2X2 U923 ( .A(n852), .B(n853), .S0(n1039), .Y(n565) );
  CLKMX2X2 U924 ( .A(n850), .B(n851), .S0(n1038), .Y(n566) );
  CLKMX2X2 U925 ( .A(n848), .B(n849), .S0(n1040), .Y(n567) );
  CLKMX2X2 U926 ( .A(n846), .B(n847), .S0(n1039), .Y(n568) );
  CLKMX2X2 U927 ( .A(n844), .B(n845), .S0(n1040), .Y(n569) );
  CLKMX2X2 U928 ( .A(n842), .B(n843), .S0(n1040), .Y(n570) );
  CLKMX2X2 U929 ( .A(n840), .B(n841), .S0(n1040), .Y(n571) );
  CLKMX2X2 U930 ( .A(n838), .B(n839), .S0(n1040), .Y(n572) );
  CLKMX2X2 U931 ( .A(n836), .B(n837), .S0(n1040), .Y(n573) );
  CLKMX2X2 U932 ( .A(n834), .B(n835), .S0(n1040), .Y(n574) );
  CLKMX2X2 U933 ( .A(n832), .B(n833), .S0(n1040), .Y(n575) );
  CLKMX2X2 U934 ( .A(n830), .B(n831), .S0(n1040), .Y(n576) );
  CLKMX2X2 U935 ( .A(n828), .B(n829), .S0(n1040), .Y(n577) );
  CLKMX2X2 U936 ( .A(n826), .B(n827), .S0(n1040), .Y(n578) );
  CLKMX2X2 U937 ( .A(n824), .B(n825), .S0(n1040), .Y(n579) );
  CLKMX2X2 U938 ( .A(n822), .B(n823), .S0(n1040), .Y(n580) );
  CLKMX2X2 U939 ( .A(n820), .B(n821), .S0(n1041), .Y(n581) );
  CLKMX2X2 U940 ( .A(n818), .B(n819), .S0(n1038), .Y(n582) );
  CLKMX2X2 U941 ( .A(n816), .B(n817), .S0(n1037), .Y(n583) );
  CLKMX2X2 U942 ( .A(n814), .B(n815), .S0(n1035), .Y(n584) );
  CLKMX2X2 U943 ( .A(n812), .B(n813), .S0(n1036), .Y(n585) );
  CLKMX2X2 U944 ( .A(n810), .B(n811), .S0(n1037), .Y(n586) );
  CLKMX2X2 U945 ( .A(n808), .B(n809), .S0(n1035), .Y(n587) );
  CLKMX2X2 U946 ( .A(n916), .B(n917), .S0(n1041), .Y(n588) );
  CLKMX2X2 U947 ( .A(n914), .B(n915), .S0(n1041), .Y(n589) );
  CLKMX2X2 U948 ( .A(n912), .B(n913), .S0(n1041), .Y(n590) );
  CLKMX2X2 U949 ( .A(n910), .B(n911), .S0(n1041), .Y(n591) );
  CLKMX2X2 U950 ( .A(n908), .B(n909), .S0(n1041), .Y(n592) );
  CLKMX2X2 U951 ( .A(n906), .B(n907), .S0(n1041), .Y(n593) );
  CLKMX2X2 U952 ( .A(n904), .B(n905), .S0(n1041), .Y(n594) );
  CLKMX2X2 U953 ( .A(n902), .B(n903), .S0(n1041), .Y(n595) );
  CLKMX2X2 U954 ( .A(n900), .B(n901), .S0(n1041), .Y(n596) );
  CLKMX2X2 U955 ( .A(n898), .B(n899), .S0(n1041), .Y(n597) );
  CLKMX2X2 U956 ( .A(n896), .B(n897), .S0(n1041), .Y(n598) );
  CLKMX2X2 U957 ( .A(n894), .B(n895), .S0(n1041), .Y(n599) );
  CLKMX2X2 U958 ( .A(n892), .B(n893), .S0(n1040), .Y(n600) );
  CLKMX2X2 U959 ( .A(n890), .B(n891), .S0(n1041), .Y(n601) );
  CLKMX2X2 U960 ( .A(n888), .B(n889), .S0(n1039), .Y(n602) );
  CLKMX2X2 U961 ( .A(n886), .B(n887), .S0(n1042), .Y(n603) );
  CLKMX2X2 U962 ( .A(n884), .B(n885), .S0(n1042), .Y(n604) );
  CLKMX2X2 U963 ( .A(n882), .B(n883), .S0(n1042), .Y(n605) );
  CLKMX2X2 U964 ( .A(n880), .B(n881), .S0(n1044), .Y(n606) );
  CLKMX2X2 U965 ( .A(n878), .B(n879), .S0(N33), .Y(n607) );
  CLKMX2X2 U966 ( .A(n876), .B(n877), .S0(N33), .Y(n608) );
  CLKMX2X2 U967 ( .A(n874), .B(n875), .S0(N33), .Y(n609) );
  CLKMX2X2 U968 ( .A(n872), .B(n873), .S0(N33), .Y(n610) );
  OR2X1 U969 ( .A(n1177), .B(proc_read), .Y(n611) );
  CLKINVX1 U970 ( .A(n612), .Y(n613) );
  CLKINVX1 U971 ( .A(mem_ready), .Y(n612) );
  CLKINVX1 U972 ( .A(proc_reset), .Y(n614) );
  INVX3 U973 ( .A(n614), .Y(n615) );
  BUFX4 U974 ( .A(n1032), .Y(n1004) );
  CLKBUFX6 U975 ( .A(n262), .Y(n1070) );
  BUFX2 U976 ( .A(n1006), .Y(n1027) );
  CLKBUFX3 U977 ( .A(n1169), .Y(n1029) );
  CLKBUFX2 U978 ( .A(n1167), .Y(n1034) );
  CLKINVX1 U979 ( .A(N31), .Y(n1171) );
  CLKINVX1 U980 ( .A(n1171), .Y(n677) );
  NAND2XL U981 ( .A(n164), .B(n144), .Y(n267) );
  CLKBUFX3 U982 ( .A(n1033), .Y(n1044) );
  XNOR2X1 U983 ( .A(proc_addr[13]), .B(n554), .Y(n450) );
  NAND2X1 U984 ( .A(n952), .B(n616), .Y(n617) );
  NAND2X1 U985 ( .A(n953), .B(n1044), .Y(n618) );
  INVXL U986 ( .A(n1044), .Y(n616) );
  MXI4XL U987 ( .A(\blocktag[0][8] ), .B(\blocktag[1][8] ), .C(
        \blocktag[2][8] ), .D(\blocktag[3][8] ), .S0(n998), .S1(n1002), .Y(
        n952) );
  MXI4XL U988 ( .A(\blocktag[4][8] ), .B(\blocktag[5][8] ), .C(
        \blocktag[6][8] ), .D(\blocktag[7][8] ), .S0(n998), .S1(n1031), .Y(
        n953) );
  INVXL U989 ( .A(n554), .Y(n1208) );
  CLKBUFX2 U990 ( .A(n1167), .Y(n1033) );
  NOR2BX4 U991 ( .AN(n504), .B(n431), .Y(n340) );
  CLKBUFX3 U992 ( .A(n974), .Y(n999) );
  CLKBUFX3 U993 ( .A(n974), .Y(n998) );
  CLKBUFX3 U994 ( .A(N31), .Y(n1000) );
  AND2X2 U995 ( .A(n261), .B(n165), .Y(n259) );
  XNOR2X1 U996 ( .A(n547), .B(proc_addr[22]), .Y(n448) );
  XNOR2X1 U997 ( .A(n550), .B(proc_addr[29]), .Y(n455) );
  XNOR2X1 U998 ( .A(n545), .B(proc_addr[11]), .Y(n462) );
  XNOR2X1 U999 ( .A(n549), .B(proc_addr[24]), .Y(n447) );
  XNOR2X1 U1000 ( .A(n548), .B(proc_addr[23]), .Y(n454) );
  XNOR2X1 U1001 ( .A(n543), .B(proc_addr[7]), .Y(n461) );
  XNOR2X1 U1002 ( .A(n546), .B(proc_addr[21]), .Y(n449) );
  XNOR2X1 U1003 ( .A(n544), .B(proc_addr[10]), .Y(n456) );
  XNOR2X1 U1004 ( .A(n542), .B(proc_addr[12]), .Y(n463) );
  NAND3X1 U1005 ( .A(n450), .B(n451), .C(n452), .Y(n446) );
  XNOR2X1 U1006 ( .A(proc_addr[18]), .B(tag[13]), .Y(n452) );
  XNOR2X1 U1007 ( .A(proc_addr[9]), .B(tag[4]), .Y(n451) );
  NAND3X1 U1008 ( .A(n457), .B(n458), .C(n459), .Y(n453) );
  XNOR2X1 U1009 ( .A(proc_addr[14]), .B(tag[9]), .Y(n457) );
  XNOR2X1 U1010 ( .A(proc_addr[20]), .B(tag[15]), .Y(n459) );
  XNOR2X1 U1011 ( .A(proc_addr[19]), .B(tag[14]), .Y(n458) );
  NAND3X1 U1012 ( .A(n464), .B(n465), .C(n466), .Y(n460) );
  XNOR2X1 U1013 ( .A(proc_addr[16]), .B(tag[11]), .Y(n464) );
  XNOR2X1 U1014 ( .A(proc_addr[26]), .B(tag[21]), .Y(n466) );
  XNOR2X1 U1015 ( .A(proc_addr[15]), .B(tag[10]), .Y(n465) );
  BUFX2 U1016 ( .A(n1005), .Y(n1028) );
  CLKBUFX2 U1017 ( .A(n1032), .Y(n1003) );
  BUFX2 U1018 ( .A(n973), .Y(n975) );
  CLKBUFX2 U1019 ( .A(n1032), .Y(n1002) );
  CLKBUFX2 U1020 ( .A(n342), .Y(n1057) );
  CLKBUFX2 U1021 ( .A(n276), .Y(n1064) );
  CLKBUFX2 U1022 ( .A(n14), .Y(n1089) );
  NOR2XL U1023 ( .A(n1167), .B(n1169), .Y(n470) );
  OAI211XL U1024 ( .A0(n1174), .A1(n1177), .B0(n1175), .C0(n1179), .Y(
        proc_stall) );
  NAND3X1 U1025 ( .A(n1258), .B(n1257), .C(n143), .Y(n15) );
  AND4X4 U1026 ( .A(n263), .B(n1175), .C(n341), .D(n430), .Y(n266) );
  BUFX2 U1027 ( .A(n260), .Y(n1071) );
  INVXL U1028 ( .A(tag[0]), .Y(n1204) );
  INVXL U1029 ( .A(tag[1]), .Y(n1205) );
  INVXL U1030 ( .A(tag[3]), .Y(n1206) );
  INVXL U1031 ( .A(tag[20]), .Y(n1215) );
  NOR2XL U1032 ( .A(n1170), .B(n1167), .Y(n469) );
  NOR2XL U1033 ( .A(n1168), .B(n1169), .Y(n468) );
  MXI4XL U1034 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n996), .S1(n1027), .Y(n918) );
  MXI4XL U1035 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n996), .S1(n1027), .Y(n919) );
  OAI2BB1XL U1036 ( .A0N(n165), .A1N(n613), .B0(dirty), .Y(n163) );
  NOR4X1 U1037 ( .A(n255), .B(n256), .C(n257), .D(n613), .Y(n1419) );
  MX2X1 U1038 ( .A(n678), .B(n679), .S0(n1042), .Y(valid) );
  MX4XL U1039 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n995), .S1(n1027), .Y(n678) );
  MX4XL U1040 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n995), .S1(n1027), .Y(n679) );
  NAND3X1 U1041 ( .A(n143), .B(n1258), .C(proc_addr[1]), .Y(n11) );
  NAND3X1 U1042 ( .A(n143), .B(n1257), .C(proc_addr[0]), .Y(n9) );
  MX4XL U1043 ( .A(n619), .B(n620), .C(n621), .D(n622), .S0(n996), .S1(n1031), 
        .Y(n920) );
  MX4XL U1044 ( .A(n623), .B(n624), .C(n625), .D(n626), .S0(n996), .S1(n1030), 
        .Y(n931) );
  MX4XL U1045 ( .A(n627), .B(n628), .C(n629), .D(n630), .S0(n996), .S1(n1030), 
        .Y(n926) );
  MX4XL U1046 ( .A(n631), .B(n632), .C(n633), .D(n634), .S0(n996), .S1(n1030), 
        .Y(n927) );
  MX4XL U1047 ( .A(n635), .B(n636), .C(n637), .D(n638), .S0(n996), .S1(n1030), 
        .Y(n924) );
  MX4XL U1048 ( .A(n639), .B(n640), .C(n641), .D(n642), .S0(n996), .S1(n1031), 
        .Y(n922) );
  MX4XL U1049 ( .A(n643), .B(n644), .C(n645), .D(n646), .S0(n996), .S1(n1031), 
        .Y(n923) );
  MX4X1 U1050 ( .A(n647), .B(n1172), .C(n648), .D(n649), .S0(n999), .S1(n1028), 
        .Y(n969) );
  MXI2X1 U1051 ( .A(n651), .B(n652), .S0(n1042), .Y(n650) );
  MX4X1 U1052 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n995), .S1(n1026), .Y(n651) );
  MX4X1 U1053 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n995), .S1(n1026), .Y(n652) );
  MXI2X1 U1054 ( .A(n654), .B(n655), .S0(n1042), .Y(n653) );
  MX4X1 U1055 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n995), .S1(n1026), .Y(n654) );
  MX4X1 U1056 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n995), .S1(n1026), .Y(n655) );
  MXI2X1 U1057 ( .A(n657), .B(n658), .S0(n1042), .Y(n656) );
  MX4X1 U1058 ( .A(\block[0][5] ), .B(\block[1][5] ), .C(\block[2][5] ), .D(
        \block[3][5] ), .S0(n995), .S1(n1026), .Y(n657) );
  MX4X1 U1059 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n994), .S1(n1026), .Y(n658) );
  MXI2X1 U1060 ( .A(n660), .B(n661), .S0(n1042), .Y(n659) );
  MX4X1 U1061 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n994), .S1(n1026), .Y(n660) );
  MX4X1 U1062 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n994), .S1(n1026), .Y(n661) );
  MXI2X1 U1063 ( .A(n663), .B(n664), .S0(n1042), .Y(n662) );
  MX4X1 U1064 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n994), .S1(n1026), .Y(n663) );
  MX4X1 U1065 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n994), .S1(n1026), .Y(n664) );
  MXI2X1 U1066 ( .A(n666), .B(n667), .S0(n1042), .Y(n665) );
  MX4X1 U1067 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n994), .S1(n1026), .Y(n666) );
  MX4X1 U1068 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n994), .S1(n1026), .Y(n667) );
  MXI2X1 U1069 ( .A(n669), .B(n670), .S0(n1042), .Y(n668) );
  MX4XL U1070 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n995), .S1(n1027), .Y(n669) );
  MX4XL U1071 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n995), .S1(n1027), .Y(n670) );
  MXI2X1 U1072 ( .A(n672), .B(n673), .S0(n1042), .Y(n671) );
  MX4XL U1073 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n995), .S1(n1027), .Y(n672) );
  MX4XL U1074 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n995), .S1(n1027), .Y(n673) );
  MXI2X1 U1075 ( .A(n675), .B(n676), .S0(n1042), .Y(n674) );
  MX4XL U1076 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n995), .S1(n1027), .Y(n675) );
  MX4XL U1077 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n995), .S1(n1027), .Y(n676) );
  NOR2X1 U1078 ( .A(proc_read), .B(proc_write), .Y(n257) );
  CLKINVX1 U1079 ( .A(proc_addr[1]), .Y(n1257) );
  CLKINVX1 U1080 ( .A(proc_addr[0]), .Y(n1258) );
  INVX1 U1081 ( .A(proc_write), .Y(n1177) );
  NAND3X1 U1082 ( .A(proc_addr[0]), .B(n1257), .C(n164), .Y(n341) );
  NAND3X1 U1083 ( .A(n1258), .B(n1257), .C(n164), .Y(n263) );
  CLKBUFX3 U1084 ( .A(n1006), .Y(n1026) );
  CLKBUFX3 U1085 ( .A(n1001), .Y(n1025) );
  CLKBUFX3 U1086 ( .A(n1026), .Y(n1024) );
  CLKBUFX3 U1087 ( .A(n1026), .Y(n1023) );
  CLKBUFX3 U1088 ( .A(n1001), .Y(n1022) );
  CLKBUFX3 U1089 ( .A(n1001), .Y(n1021) );
  CLKBUFX3 U1090 ( .A(n1001), .Y(n1020) );
  CLKBUFX3 U1091 ( .A(n1001), .Y(n1019) );
  CLKBUFX3 U1092 ( .A(n1001), .Y(n1018) );
  CLKBUFX3 U1093 ( .A(n1001), .Y(n1017) );
  CLKBUFX3 U1094 ( .A(n1001), .Y(n1016) );
  CLKBUFX3 U1095 ( .A(n1001), .Y(n1015) );
  CLKBUFX3 U1096 ( .A(n1001), .Y(n1014) );
  CLKBUFX3 U1097 ( .A(n1001), .Y(n1013) );
  CLKBUFX3 U1098 ( .A(n1001), .Y(n1012) );
  CLKBUFX3 U1099 ( .A(n1001), .Y(n1011) );
  CLKBUFX3 U1100 ( .A(n1001), .Y(n1010) );
  CLKBUFX3 U1101 ( .A(n1001), .Y(n1009) );
  CLKBUFX3 U1102 ( .A(n1001), .Y(n1008) );
  CLKBUFX3 U1103 ( .A(n1034), .Y(n1043) );
  CLKBUFX3 U1104 ( .A(n1034), .Y(n1042) );
  CLKBUFX3 U1105 ( .A(n976), .Y(n995) );
  CLKBUFX3 U1106 ( .A(n975), .Y(n997) );
  CLKBUFX3 U1107 ( .A(n975), .Y(n996) );
  CLKBUFX3 U1108 ( .A(n1004), .Y(n1005) );
  CLKBUFX3 U1109 ( .A(n1003), .Y(n1006) );
  CLKBUFX3 U1110 ( .A(n1037), .Y(n1041) );
  CLKBUFX3 U1111 ( .A(n1036), .Y(n1040) );
  CLKBUFX3 U1112 ( .A(n1035), .Y(n1039) );
  CLKBUFX3 U1113 ( .A(n1036), .Y(n1038) );
  CLKBUFX3 U1114 ( .A(n1042), .Y(n1037) );
  CLKBUFX3 U1115 ( .A(n976), .Y(n994) );
  CLKBUFX3 U1116 ( .A(n971), .Y(n993) );
  CLKBUFX3 U1117 ( .A(n971), .Y(n992) );
  CLKBUFX3 U1118 ( .A(n971), .Y(n991) );
  CLKBUFX3 U1119 ( .A(n971), .Y(n990) );
  CLKBUFX3 U1120 ( .A(n971), .Y(n989) );
  CLKBUFX3 U1121 ( .A(n971), .Y(n988) );
  CLKBUFX3 U1122 ( .A(n977), .Y(n987) );
  CLKBUFX3 U1123 ( .A(n971), .Y(n986) );
  CLKBUFX3 U1124 ( .A(n971), .Y(n985) );
  CLKBUFX3 U1125 ( .A(n977), .Y(n984) );
  CLKBUFX3 U1126 ( .A(n977), .Y(n983) );
  CLKBUFX3 U1127 ( .A(n970), .Y(n982) );
  CLKBUFX3 U1128 ( .A(n970), .Y(n981) );
  CLKBUFX3 U1129 ( .A(n977), .Y(n980) );
  CLKBUFX3 U1130 ( .A(n977), .Y(n979) );
  CLKBUFX3 U1131 ( .A(n970), .Y(n978) );
  CLKBUFX3 U1132 ( .A(n972), .Y(n976) );
  CLKBUFX3 U1133 ( .A(n973), .Y(n974) );
  CLKBUFX3 U1134 ( .A(n1176), .Y(n1053) );
  CLKBUFX3 U1135 ( .A(n1176), .Y(n1054) );
  CLKBUFX3 U1136 ( .A(n1176), .Y(n1050) );
  CLKBUFX3 U1137 ( .A(n1176), .Y(n1051) );
  CLKBUFX3 U1138 ( .A(n1042), .Y(n1036) );
  CLKBUFX3 U1139 ( .A(n1042), .Y(n1035) );
  CLKBUFX3 U1140 ( .A(n1001), .Y(n1007) );
  CLKBUFX3 U1141 ( .A(n1031), .Y(n1001) );
  CLKBUFX3 U1142 ( .A(n971), .Y(n977) );
  CLKBUFX3 U1143 ( .A(n342), .Y(n1056) );
  CLKBUFX3 U1144 ( .A(n342), .Y(n1055) );
  CLKBUFX3 U1145 ( .A(n276), .Y(n1063) );
  CLKBUFX3 U1146 ( .A(n276), .Y(n1062) );
  CLKBUFX3 U1147 ( .A(n1000), .Y(n972) );
  CLKBUFX3 U1148 ( .A(n1000), .Y(n973) );
  CLKBUFX3 U1149 ( .A(n1029), .Y(n1032) );
  CLKBUFX3 U1150 ( .A(n1176), .Y(n1046) );
  CLKBUFX3 U1151 ( .A(n1158), .Y(n1159) );
  CLKBUFX3 U1152 ( .A(n1158), .Y(n1160) );
  CLKBUFX3 U1153 ( .A(n1158), .Y(n1161) );
  CLKBUFX3 U1154 ( .A(n1158), .Y(n1162) );
  CLKBUFX3 U1155 ( .A(n1158), .Y(n1163) );
  CLKBUFX3 U1156 ( .A(n1158), .Y(n1164) );
  CLKBUFX3 U1157 ( .A(n1158), .Y(n1165) );
  CLKBUFX3 U1158 ( .A(N1769), .Y(n1149) );
  CLKBUFX3 U1159 ( .A(N1769), .Y(n1150) );
  CLKBUFX3 U1160 ( .A(n1150), .Y(n1151) );
  CLKBUFX3 U1161 ( .A(n1150), .Y(n1152) );
  CLKBUFX3 U1162 ( .A(n1150), .Y(n1153) );
  CLKBUFX3 U1163 ( .A(n1150), .Y(n1154) );
  CLKBUFX3 U1164 ( .A(n1150), .Y(n1155) );
  CLKBUFX3 U1165 ( .A(n1140), .Y(n1141) );
  CLKBUFX3 U1166 ( .A(n1140), .Y(n1142) );
  CLKBUFX3 U1167 ( .A(n1140), .Y(n1143) );
  CLKBUFX3 U1168 ( .A(n1140), .Y(n1144) );
  CLKBUFX3 U1169 ( .A(n1140), .Y(n1145) );
  CLKBUFX3 U1170 ( .A(n1140), .Y(n1146) );
  CLKBUFX3 U1171 ( .A(n1140), .Y(n1147) );
  CLKBUFX3 U1172 ( .A(n1131), .Y(n1132) );
  CLKBUFX3 U1173 ( .A(n1131), .Y(n1133) );
  CLKBUFX3 U1174 ( .A(n1131), .Y(n1134) );
  CLKBUFX3 U1175 ( .A(n1131), .Y(n1135) );
  CLKBUFX3 U1176 ( .A(n1131), .Y(n1136) );
  CLKBUFX3 U1177 ( .A(n1131), .Y(n1137) );
  CLKBUFX3 U1178 ( .A(n1131), .Y(n1138) );
  CLKBUFX3 U1179 ( .A(n1122), .Y(n1123) );
  CLKBUFX3 U1180 ( .A(n1122), .Y(n1124) );
  CLKBUFX3 U1181 ( .A(n1122), .Y(n1125) );
  CLKBUFX3 U1182 ( .A(n1122), .Y(n1126) );
  CLKBUFX3 U1183 ( .A(n1122), .Y(n1127) );
  CLKBUFX3 U1184 ( .A(n1122), .Y(n1128) );
  CLKBUFX3 U1185 ( .A(n1122), .Y(n1129) );
  CLKBUFX3 U1186 ( .A(n1113), .Y(n1114) );
  CLKBUFX3 U1187 ( .A(n1113), .Y(n1115) );
  CLKBUFX3 U1188 ( .A(n1113), .Y(n1116) );
  CLKBUFX3 U1189 ( .A(n1113), .Y(n1117) );
  CLKBUFX3 U1190 ( .A(n1113), .Y(n1118) );
  CLKBUFX3 U1191 ( .A(n1113), .Y(n1119) );
  CLKBUFX3 U1192 ( .A(n1113), .Y(n1120) );
  CLKBUFX3 U1193 ( .A(N1776), .Y(n1104) );
  CLKBUFX3 U1194 ( .A(N1776), .Y(n1105) );
  CLKBUFX3 U1195 ( .A(N1776), .Y(n1106) );
  CLKBUFX3 U1196 ( .A(n1105), .Y(n1107) );
  CLKBUFX3 U1197 ( .A(n1105), .Y(n1108) );
  CLKBUFX3 U1198 ( .A(N1776), .Y(n1109) );
  CLKBUFX3 U1199 ( .A(N1776), .Y(n1110) );
  CLKBUFX3 U1200 ( .A(n1105), .Y(n1111) );
  CLKBUFX3 U1201 ( .A(n1095), .Y(n1096) );
  CLKBUFX3 U1202 ( .A(n1095), .Y(n1097) );
  CLKBUFX3 U1203 ( .A(n1095), .Y(n1098) );
  CLKBUFX3 U1204 ( .A(n1095), .Y(n1099) );
  CLKBUFX3 U1205 ( .A(n1095), .Y(n1100) );
  CLKBUFX3 U1206 ( .A(n1095), .Y(n1101) );
  CLKBUFX3 U1207 ( .A(n1095), .Y(n1102) );
  CLKBUFX3 U1208 ( .A(n1158), .Y(n1166) );
  CLKBUFX3 U1209 ( .A(N1769), .Y(n1156) );
  CLKBUFX3 U1210 ( .A(n1140), .Y(n1148) );
  CLKBUFX3 U1211 ( .A(n1131), .Y(n1139) );
  CLKBUFX3 U1212 ( .A(n1122), .Y(n1130) );
  CLKBUFX3 U1213 ( .A(n1113), .Y(n1121) );
  CLKBUFX3 U1214 ( .A(N1776), .Y(n1112) );
  CLKBUFX3 U1215 ( .A(n1095), .Y(n1103) );
  CLKBUFX3 U1216 ( .A(n1150), .Y(n1157) );
  CLKBUFX3 U1217 ( .A(n1000), .Y(n971) );
  CLKBUFX3 U1218 ( .A(n971), .Y(n970) );
  CLKINVX1 U1219 ( .A(n150), .Y(n1256) );
  CLKINVX1 U1220 ( .A(n154), .Y(n1254) );
  CLKINVX1 U1221 ( .A(n158), .Y(n1252) );
  CLKINVX1 U1222 ( .A(n162), .Y(n1250) );
  CLKBUFX3 U1223 ( .A(n504), .Y(n1065) );
  CLKBUFX3 U1224 ( .A(n504), .Y(n1066) );
  CLKBUFX3 U1225 ( .A(n266), .Y(n1068) );
  CLKBUFX3 U1226 ( .A(n266), .Y(n1067) );
  CLKINVX1 U1227 ( .A(n145), .Y(n1179) );
  CLKBUFX3 U1228 ( .A(n1071), .Y(n1073) );
  CLKBUFX3 U1229 ( .A(n259), .Y(n1082) );
  CLKBUFX3 U1230 ( .A(n259), .Y(n1081) );
  CLKBUFX3 U1231 ( .A(n260), .Y(n1078) );
  CLKBUFX3 U1232 ( .A(n260), .Y(n1077) );
  CLKBUFX3 U1233 ( .A(n1071), .Y(n1076) );
  CLKBUFX3 U1234 ( .A(n1071), .Y(n1075) );
  CLKBUFX3 U1235 ( .A(n1071), .Y(n1074) );
  CLKBUFX3 U1236 ( .A(n260), .Y(n1080) );
  CLKBUFX3 U1237 ( .A(n1071), .Y(n1079) );
  CLKBUFX3 U1238 ( .A(n1071), .Y(n1072) );
  CLKBUFX3 U1239 ( .A(n14), .Y(n1088) );
  INVX3 U1240 ( .A(mem_read), .Y(n1083) );
  INVX3 U1241 ( .A(mem_read), .Y(n1084) );
  CLKBUFX3 U1242 ( .A(n15), .Y(n1085) );
  CLKBUFX3 U1243 ( .A(n15), .Y(n1086) );
  NOR2X1 U1244 ( .A(n1217), .B(n1045), .Y(mem_wdata[96]) );
  NOR2X1 U1245 ( .A(n1218), .B(n1048), .Y(mem_wdata[97]) );
  NOR2X1 U1246 ( .A(n1219), .B(n1176), .Y(mem_wdata[98]) );
  NOR2X1 U1247 ( .A(n1220), .B(n1045), .Y(mem_wdata[99]) );
  NOR2X1 U1248 ( .A(n1221), .B(n1054), .Y(mem_wdata[100]) );
  NOR2X1 U1249 ( .A(n1222), .B(n1054), .Y(mem_wdata[101]) );
  NOR2X1 U1250 ( .A(n1223), .B(n1045), .Y(mem_wdata[102]) );
  NOR2X1 U1251 ( .A(n1224), .B(n1048), .Y(mem_wdata[103]) );
  NOR2X1 U1252 ( .A(n1225), .B(n1054), .Y(mem_wdata[104]) );
  NOR2X1 U1253 ( .A(n1226), .B(n1049), .Y(mem_wdata[105]) );
  NOR2X1 U1254 ( .A(n1227), .B(n1052), .Y(mem_wdata[106]) );
  NOR2X1 U1255 ( .A(n1228), .B(n1053), .Y(mem_wdata[107]) );
  NOR2X1 U1256 ( .A(n1229), .B(n1051), .Y(mem_wdata[108]) );
  NOR2X1 U1257 ( .A(n1230), .B(n1049), .Y(mem_wdata[109]) );
  NOR2X1 U1258 ( .A(n1231), .B(n1051), .Y(mem_wdata[110]) );
  NOR2X1 U1259 ( .A(n1232), .B(n1052), .Y(mem_wdata[111]) );
  NOR2X1 U1260 ( .A(n1233), .B(n1047), .Y(mem_wdata[112]) );
  NOR2X1 U1261 ( .A(n1234), .B(n1050), .Y(mem_wdata[113]) );
  NOR2X1 U1262 ( .A(n1235), .B(n1046), .Y(mem_wdata[114]) );
  NOR2X1 U1263 ( .A(n1236), .B(n1047), .Y(mem_wdata[115]) );
  NOR2X1 U1264 ( .A(n1237), .B(n1049), .Y(mem_wdata[116]) );
  NOR2X1 U1265 ( .A(n1238), .B(n1049), .Y(mem_wdata[117]) );
  NOR2X1 U1266 ( .A(n1239), .B(n1050), .Y(mem_wdata[118]) );
  NOR2X1 U1267 ( .A(n1240), .B(n1048), .Y(mem_wdata[119]) );
  NOR2X1 U1268 ( .A(n1241), .B(n1053), .Y(mem_wdata[120]) );
  NOR2X1 U1269 ( .A(n1242), .B(n1051), .Y(mem_wdata[121]) );
  NOR2X1 U1270 ( .A(n1243), .B(n1046), .Y(mem_wdata[122]) );
  NOR2X1 U1271 ( .A(n1244), .B(n1046), .Y(mem_wdata[123]) );
  NOR2X1 U1272 ( .A(n1245), .B(n1052), .Y(mem_wdata[124]) );
  NOR2X1 U1273 ( .A(n1246), .B(n1047), .Y(mem_wdata[125]) );
  NOR2X1 U1274 ( .A(n1247), .B(n1050), .Y(mem_wdata[126]) );
  NOR2X1 U1275 ( .A(n1248), .B(n1046), .Y(mem_wdata[127]) );
  CLKBUFX3 U1276 ( .A(n15), .Y(n1087) );
  NAND2X1 U1277 ( .A(n677), .B(n470), .Y(n150) );
  NAND2X1 U1278 ( .A(n469), .B(N31), .Y(n154) );
  NAND2X1 U1279 ( .A(n468), .B(N31), .Y(n158) );
  NAND2X1 U1280 ( .A(n467), .B(N31), .Y(n162) );
  CLKINVX1 U1281 ( .A(n148), .Y(n1255) );
  CLKINVX1 U1282 ( .A(n152), .Y(n1253) );
  CLKINVX1 U1283 ( .A(n156), .Y(n1251) );
  CLKINVX1 U1284 ( .A(n160), .Y(n1249) );
  NOR4X1 U1285 ( .A(n460), .B(n461), .C(n462), .D(n463), .Y(n434) );
  NOR4X1 U1286 ( .A(n453), .B(n454), .C(n455), .D(n456), .Y(n435) );
  CLKBUFX3 U1287 ( .A(n505), .Y(n1060) );
  CLKBUFX3 U1288 ( .A(n505), .Y(n1061) );
  CLKBUFX3 U1289 ( .A(n341), .Y(n1058) );
  CLKBUFX3 U1290 ( .A(n341), .Y(n1059) );
  CLKINVX1 U1291 ( .A(n1168), .Y(n1167) );
  OAI22X2 U1292 ( .A0(n1082), .A1(n1204), .B0(n1203), .B1(n1073), .Y(
        blocktag_next[0]) );
  OAI22X2 U1293 ( .A0(n1082), .A1(n1205), .B0(n1202), .B1(n1072), .Y(
        blocktag_next[1]) );
  OAI22X2 U1294 ( .A0(n1081), .A1(n543), .B0(n1201), .B1(n1080), .Y(
        blocktag_next[2]) );
  OAI22X2 U1295 ( .A0(n1081), .A1(n1206), .B0(n1200), .B1(n1078), .Y(
        blocktag_next[3]) );
  OAI22X2 U1296 ( .A0(n1081), .A1(n1207), .B0(n1199), .B1(n1077), .Y(
        blocktag_next[4]) );
  OAI22X2 U1297 ( .A0(n1081), .A1(n544), .B0(n1198), .B1(n1080), .Y(
        blocktag_next[5]) );
  OAI22X2 U1298 ( .A0(n1081), .A1(n545), .B0(n1197), .B1(n1078), .Y(
        blocktag_next[6]) );
  OAI22X2 U1299 ( .A0(n1081), .A1(n542), .B0(n1196), .B1(n1077), .Y(
        blocktag_next[7]) );
  OAI22X2 U1300 ( .A0(n1081), .A1(n1208), .B0(n1195), .B1(n1080), .Y(
        blocktag_next[8]) );
  OAI22X2 U1301 ( .A0(n1081), .A1(n1209), .B0(n1194), .B1(n1078), .Y(
        blocktag_next[9]) );
  OAI22X2 U1302 ( .A0(n1082), .A1(n1210), .B0(n1193), .B1(n1072), .Y(
        blocktag_next[10]) );
  OAI22X2 U1303 ( .A0(n1082), .A1(n1211), .B0(n1192), .B1(n1072), .Y(
        blocktag_next[11]) );
  OAI22X2 U1304 ( .A0(n1082), .A1(n552), .B0(n1191), .B1(n1072), .Y(
        blocktag_next[12]) );
  OAI22X2 U1305 ( .A0(n1082), .A1(n1212), .B0(n1190), .B1(n1072), .Y(
        blocktag_next[13]) );
  OAI22X2 U1306 ( .A0(n1082), .A1(n1213), .B0(n1189), .B1(n1072), .Y(
        blocktag_next[14]) );
  OAI22X2 U1307 ( .A0(n1082), .A1(n1214), .B0(n1188), .B1(n1072), .Y(
        blocktag_next[15]) );
  OAI22X2 U1308 ( .A0(n1082), .A1(n546), .B0(n1187), .B1(n1072), .Y(
        blocktag_next[16]) );
  OAI22X2 U1309 ( .A0(n1082), .A1(n547), .B0(n1186), .B1(n1072), .Y(
        blocktag_next[17]) );
  OAI22X2 U1310 ( .A0(n1082), .A1(n548), .B0(n1185), .B1(n1072), .Y(
        blocktag_next[18]) );
  OAI22X2 U1311 ( .A0(n1082), .A1(n549), .B0(n1184), .B1(n1072), .Y(
        blocktag_next[19]) );
  OAI22X2 U1312 ( .A0(n1082), .A1(n1215), .B0(n1183), .B1(n1072), .Y(
        blocktag_next[20]) );
  OAI22X2 U1313 ( .A0(n1081), .A1(n1216), .B0(n1182), .B1(n1077), .Y(
        blocktag_next[21]) );
  OAI22X2 U1314 ( .A0(n1081), .A1(n553), .B0(n1181), .B1(n1079), .Y(
        blocktag_next[22]) );
  OAI22X2 U1315 ( .A0(n1081), .A1(n551), .B0(n1180), .B1(n1075), .Y(
        blocktag_next[23]) );
  OAI22X2 U1316 ( .A0(n1081), .A1(n550), .B0(n1178), .B1(n1076), .Y(
        blocktag_next[24]) );
  OAI221XL U1317 ( .A0(n1094), .A1(n557), .B0(n1091), .B1(n511), .C0(n95), .Y(
        proc_rdata[1]) );
  AOI2BB2X1 U1318 ( .B0(blockdata[97]), .B1(n1088), .A0N(n1085), .A1N(n671), 
        .Y(n95) );
  OAI221XL U1319 ( .A0(n1093), .A1(n558), .B0(n1090), .B1(n512), .C0(n51), .Y(
        proc_rdata[2]) );
  AOI2BB2X1 U1320 ( .B0(blockdata[98]), .B1(n1088), .A0N(n1086), .A1N(n674), 
        .Y(n51) );
  OAI221XL U1321 ( .A0(n1093), .A1(n559), .B0(n1090), .B1(n513), .C0(n39), .Y(
        proc_rdata[3]) );
  AOI2BB2X1 U1322 ( .B0(blockdata[99]), .B1(n14), .A0N(n1087), .A1N(n650), .Y(
        n39) );
  OAI221XL U1323 ( .A0(n1093), .A1(n560), .B0(n1090), .B1(n514), .C0(n35), .Y(
        proc_rdata[4]) );
  AOI2BB2X1 U1324 ( .B0(blockdata[100]), .B1(n14), .A0N(n1087), .A1N(n653), 
        .Y(n35) );
  OAI221XL U1325 ( .A0(n1093), .A1(n561), .B0(n1090), .B1(n515), .C0(n31), .Y(
        proc_rdata[5]) );
  AOI2BB2X1 U1326 ( .B0(blockdata[101]), .B1(n14), .A0N(n1087), .A1N(n656), 
        .Y(n31) );
  OAI221XL U1327 ( .A0(n1093), .A1(n562), .B0(n1090), .B1(n516), .C0(n27), .Y(
        proc_rdata[6]) );
  AOI2BB2X1 U1328 ( .B0(blockdata[102]), .B1(n14), .A0N(n1087), .A1N(n659), 
        .Y(n27) );
  OAI221XL U1329 ( .A0(n1093), .A1(n563), .B0(n1090), .B1(n517), .C0(n23), .Y(
        proc_rdata[7]) );
  AOI2BB2X1 U1330 ( .B0(blockdata[103]), .B1(n14), .A0N(n1087), .A1N(n662), 
        .Y(n23) );
  OAI221XL U1331 ( .A0(n1093), .A1(n564), .B0(n1090), .B1(n518), .C0(n19), .Y(
        proc_rdata[8]) );
  AOI2BB2X1 U1332 ( .B0(blockdata[104]), .B1(n14), .A0N(n1087), .A1N(n665), 
        .Y(n19) );
  OAI221XL U1333 ( .A0(n1093), .A1(n565), .B0(n1090), .B1(n519), .C0(n13), .Y(
        proc_rdata[9]) );
  AOI2BB2X1 U1334 ( .B0(blockdata[105]), .B1(n14), .A0N(n1087), .A1N(n588), 
        .Y(n13) );
  OAI221XL U1335 ( .A0(n1094), .A1(n573), .B0(n1091), .B1(n527), .C0(n107), 
        .Y(proc_rdata[17]) );
  AOI2BB2X1 U1336 ( .B0(blockdata[113]), .B1(n1088), .A0N(n1085), .A1N(n596), 
        .Y(n107) );
  OAI221XL U1337 ( .A0(n1094), .A1(n574), .B0(n1091), .B1(n528), .C0(n103), 
        .Y(proc_rdata[18]) );
  AOI2BB2X1 U1338 ( .B0(blockdata[114]), .B1(n1088), .A0N(n1085), .A1N(n597), 
        .Y(n103) );
  OAI221XL U1339 ( .A0(n1094), .A1(n575), .B0(n1091), .B1(n529), .C0(n99), .Y(
        proc_rdata[19]) );
  AOI2BB2X1 U1340 ( .B0(blockdata[115]), .B1(n1088), .A0N(n1085), .A1N(n598), 
        .Y(n99) );
  OAI221XL U1341 ( .A0(n1094), .A1(n576), .B0(n1091), .B1(n530), .C0(n91), .Y(
        proc_rdata[20]) );
  AOI2BB2X1 U1342 ( .B0(blockdata[116]), .B1(n1088), .A0N(n1086), .A1N(n599), 
        .Y(n91) );
  OAI221XL U1343 ( .A0(n1094), .A1(n577), .B0(n1091), .B1(n531), .C0(n87), .Y(
        proc_rdata[21]) );
  AOI2BB2X1 U1344 ( .B0(blockdata[117]), .B1(n1088), .A0N(n1086), .A1N(n600), 
        .Y(n87) );
  OAI221XL U1345 ( .A0(n1094), .A1(n578), .B0(n1091), .B1(n532), .C0(n83), .Y(
        proc_rdata[22]) );
  AOI2BB2X1 U1346 ( .B0(blockdata[118]), .B1(n1088), .A0N(n1086), .A1N(n601), 
        .Y(n83) );
  OAI221XL U1347 ( .A0(n1094), .A1(n579), .B0(n1091), .B1(n533), .C0(n79), .Y(
        proc_rdata[23]) );
  AOI2BB2X1 U1348 ( .B0(blockdata[119]), .B1(n1088), .A0N(n1086), .A1N(n602), 
        .Y(n79) );
  OAI221XL U1349 ( .A0(n1094), .A1(n580), .B0(n1091), .B1(n534), .C0(n75), .Y(
        proc_rdata[24]) );
  AOI2BB2X1 U1350 ( .B0(blockdata[120]), .B1(n1088), .A0N(n1086), .A1N(n603), 
        .Y(n75) );
  OAI221XL U1351 ( .A0(n1094), .A1(n581), .B0(n1091), .B1(n535), .C0(n71), .Y(
        proc_rdata[25]) );
  AOI2BB2X1 U1352 ( .B0(blockdata[121]), .B1(n1088), .A0N(n1086), .A1N(n604), 
        .Y(n71) );
  OAI221XL U1353 ( .A0(n1094), .A1(n582), .B0(n1091), .B1(n536), .C0(n67), .Y(
        proc_rdata[26]) );
  AOI2BB2X1 U1354 ( .B0(blockdata[122]), .B1(n1088), .A0N(n1086), .A1N(n605), 
        .Y(n67) );
  OAI221XL U1355 ( .A0(n1094), .A1(n583), .B0(n1091), .B1(n537), .C0(n63), .Y(
        proc_rdata[27]) );
  AOI2BB2X1 U1356 ( .B0(blockdata[123]), .B1(n1088), .A0N(n1086), .A1N(n606), 
        .Y(n63) );
  OAI221XL U1357 ( .A0(n1093), .A1(n584), .B0(n1090), .B1(n538), .C0(n59), .Y(
        proc_rdata[28]) );
  AOI2BB2X1 U1358 ( .B0(blockdata[124]), .B1(n14), .A0N(n1086), .A1N(n607), 
        .Y(n59) );
  OAI221XL U1359 ( .A0(n1093), .A1(n585), .B0(n1090), .B1(n539), .C0(n55), .Y(
        proc_rdata[29]) );
  AOI2BB2X1 U1360 ( .B0(blockdata[125]), .B1(n14), .A0N(n1086), .A1N(n608), 
        .Y(n55) );
  OAI221XL U1361 ( .A0(n1093), .A1(n586), .B0(n1090), .B1(n540), .C0(n47), .Y(
        proc_rdata[30]) );
  AOI2BB2X1 U1362 ( .B0(blockdata[126]), .B1(n14), .A0N(n1086), .A1N(n609), 
        .Y(n47) );
  OAI221XL U1363 ( .A0(n1093), .A1(n587), .B0(n1090), .B1(n541), .C0(n43), .Y(
        proc_rdata[31]) );
  AOI2BB2X1 U1364 ( .B0(blockdata[127]), .B1(n14), .A0N(n1087), .A1N(n610), 
        .Y(n43) );
  OAI221XL U1365 ( .A0(n1094), .A1(n556), .B0(n1092), .B1(n510), .C0(n139), 
        .Y(proc_rdata[0]) );
  AOI2BB2X1 U1366 ( .B0(blockdata[96]), .B1(n1089), .A0N(n1085), .A1N(n668), 
        .Y(n139) );
  OAI221XL U1367 ( .A0(n1093), .A1(n566), .B0(n1092), .B1(n520), .C0(n135), 
        .Y(proc_rdata[10]) );
  AOI2BB2X1 U1368 ( .B0(blockdata[106]), .B1(n1089), .A0N(n1085), .A1N(n589), 
        .Y(n135) );
  OAI221XL U1369 ( .A0(n1094), .A1(n567), .B0(n1092), .B1(n521), .C0(n131), 
        .Y(proc_rdata[11]) );
  AOI2BB2X1 U1370 ( .B0(blockdata[107]), .B1(n1089), .A0N(n1085), .A1N(n590), 
        .Y(n131) );
  OAI221XL U1371 ( .A0(n1093), .A1(n568), .B0(n1092), .B1(n522), .C0(n127), 
        .Y(proc_rdata[12]) );
  AOI2BB2X1 U1372 ( .B0(blockdata[108]), .B1(n1089), .A0N(n1085), .A1N(n591), 
        .Y(n127) );
  OAI221XL U1373 ( .A0(n1094), .A1(n569), .B0(n1092), .B1(n523), .C0(n123), 
        .Y(proc_rdata[13]) );
  AOI2BB2X1 U1374 ( .B0(blockdata[109]), .B1(n1089), .A0N(n1085), .A1N(n592), 
        .Y(n123) );
  OAI221XL U1375 ( .A0(n1093), .A1(n570), .B0(n1092), .B1(n524), .C0(n119), 
        .Y(proc_rdata[14]) );
  AOI2BB2X1 U1376 ( .B0(blockdata[110]), .B1(n1089), .A0N(n1085), .A1N(n593), 
        .Y(n119) );
  OAI221XL U1377 ( .A0(n9), .A1(n571), .B0(n1092), .B1(n525), .C0(n115), .Y(
        proc_rdata[15]) );
  AOI2BB2X1 U1378 ( .B0(blockdata[111]), .B1(n1089), .A0N(n1085), .A1N(n594), 
        .Y(n115) );
  OAI221XL U1379 ( .A0(n9), .A1(n572), .B0(n1092), .B1(n526), .C0(n111), .Y(
        proc_rdata[16]) );
  AOI2BB2X1 U1380 ( .B0(blockdata[112]), .B1(n1089), .A0N(n1085), .A1N(n595), 
        .Y(n111) );
  NOR2X1 U1381 ( .A(mem_read), .B(n506), .Y(n215) );
  NAND2X1 U1382 ( .A(dirty), .B(valid), .Y(n255) );
  NOR2X1 U1383 ( .A(n257), .B(n1179), .Y(n165) );
  AND2X2 U1384 ( .A(n144), .B(n143), .Y(n14) );
  OAI22XL U1385 ( .A0(n542), .A1(n1052), .B0(n1196), .B1(n1083), .Y(
        mem_addr[10]) );
  OAI22XL U1386 ( .A0(n1204), .A1(n1046), .B0(n1203), .B1(n1083), .Y(
        mem_addr[3]) );
  OAI22XL U1387 ( .A0(n1205), .A1(n1047), .B0(n1202), .B1(n1083), .Y(
        mem_addr[4]) );
  OAI22XL U1388 ( .A0(n543), .A1(n1045), .B0(n1201), .B1(n1083), .Y(
        mem_addr[5]) );
  OAI22XL U1389 ( .A0(n1206), .A1(n1048), .B0(n1200), .B1(n1083), .Y(
        mem_addr[6]) );
  OAI22XL U1390 ( .A0(n1207), .A1(n1049), .B0(n1199), .B1(n1083), .Y(
        mem_addr[7]) );
  OAI22XL U1391 ( .A0(n544), .A1(n1051), .B0(n1198), .B1(n1083), .Y(
        mem_addr[8]) );
  OAI22XL U1392 ( .A0(n545), .A1(n1050), .B0(n1197), .B1(n1083), .Y(
        mem_addr[9]) );
  OAI22XL U1393 ( .A0(n1208), .A1(n1051), .B0(n1195), .B1(n1084), .Y(
        mem_addr[11]) );
  OAI22XL U1394 ( .A0(n1209), .A1(n1054), .B0(n1194), .B1(n1084), .Y(
        mem_addr[12]) );
  OAI22XL U1395 ( .A0(n1210), .A1(n1053), .B0(n1193), .B1(n1084), .Y(
        mem_addr[13]) );
  OAI22XL U1396 ( .A0(n1211), .A1(n1047), .B0(n1192), .B1(n1084), .Y(
        mem_addr[14]) );
  OAI22XL U1397 ( .A0(n552), .A1(n1050), .B0(n1191), .B1(n1084), .Y(
        mem_addr[15]) );
  OAI22XL U1398 ( .A0(n1212), .A1(n1045), .B0(n1190), .B1(n1084), .Y(
        mem_addr[16]) );
  OAI22XL U1399 ( .A0(n1213), .A1(n1052), .B0(n1189), .B1(n1084), .Y(
        mem_addr[17]) );
  OAI22XL U1400 ( .A0(n1214), .A1(n1046), .B0(n1188), .B1(n1084), .Y(
        mem_addr[18]) );
  OAI22XL U1401 ( .A0(n546), .A1(n1176), .B0(n1187), .B1(n1084), .Y(
        mem_addr[19]) );
  OAI22XL U1402 ( .A0(n547), .A1(n1053), .B0(n1186), .B1(n1084), .Y(
        mem_addr[20]) );
  OAI22XL U1403 ( .A0(n548), .A1(n1054), .B0(n1185), .B1(n1084), .Y(
        mem_addr[21]) );
  OAI22XL U1404 ( .A0(n549), .A1(n1049), .B0(n1184), .B1(n1084), .Y(
        mem_addr[22]) );
  OAI22XL U1405 ( .A0(n1215), .A1(n1046), .B0(n1183), .B1(n1083), .Y(
        mem_addr[23]) );
  OAI22XL U1406 ( .A0(n1216), .A1(n1045), .B0(n1182), .B1(n1083), .Y(
        mem_addr[24]) );
  OAI22XL U1407 ( .A0(n553), .A1(n1054), .B0(n1181), .B1(n1083), .Y(
        mem_addr[25]) );
  OAI22XL U1408 ( .A0(n551), .A1(n1048), .B0(n1180), .B1(n1083), .Y(
        mem_addr[26]) );
  OAI22XL U1409 ( .A0(n550), .A1(n1176), .B0(n1178), .B1(n1083), .Y(
        mem_addr[27]) );
  CLKBUFX3 U1410 ( .A(n11), .Y(n1091) );
  CLKBUFX3 U1411 ( .A(n11), .Y(n1090) );
  CLKBUFX3 U1412 ( .A(n9), .Y(n1094) );
  CLKBUFX3 U1413 ( .A(n9), .Y(n1093) );
  NOR2X1 U1414 ( .A(n215), .B(n1171), .Y(mem_addr[0]) );
  NOR2X1 U1415 ( .A(n215), .B(n1170), .Y(mem_addr[1]) );
  NOR2X1 U1416 ( .A(n215), .B(n1168), .Y(mem_addr[2]) );
  NOR2X1 U1417 ( .A(n510), .B(n1176), .Y(mem_wdata[64]) );
  NOR2X1 U1418 ( .A(n511), .B(n1051), .Y(mem_wdata[65]) );
  NOR2X1 U1419 ( .A(n512), .B(n1046), .Y(mem_wdata[66]) );
  NOR2X1 U1420 ( .A(n513), .B(n1054), .Y(mem_wdata[67]) );
  NOR2X1 U1421 ( .A(n514), .B(n1053), .Y(mem_wdata[68]) );
  NOR2X1 U1422 ( .A(n515), .B(n1048), .Y(mem_wdata[69]) );
  NOR2X1 U1423 ( .A(n516), .B(n1048), .Y(mem_wdata[70]) );
  NOR2X1 U1424 ( .A(n517), .B(n1176), .Y(mem_wdata[71]) );
  NOR2X1 U1425 ( .A(n518), .B(n1053), .Y(mem_wdata[72]) );
  NOR2X1 U1426 ( .A(n519), .B(n1176), .Y(mem_wdata[73]) );
  NOR2X1 U1427 ( .A(n520), .B(n1052), .Y(mem_wdata[74]) );
  NOR2X1 U1428 ( .A(n521), .B(n1049), .Y(mem_wdata[75]) );
  NOR2X1 U1429 ( .A(n522), .B(n1052), .Y(mem_wdata[76]) );
  NOR2X1 U1430 ( .A(n523), .B(n1051), .Y(mem_wdata[77]) );
  NOR2X1 U1431 ( .A(n524), .B(n1050), .Y(mem_wdata[78]) );
  NOR2X1 U1432 ( .A(n525), .B(n1052), .Y(mem_wdata[79]) );
  NOR2X1 U1433 ( .A(n526), .B(n1053), .Y(mem_wdata[80]) );
  NOR2X1 U1434 ( .A(n527), .B(n1053), .Y(mem_wdata[81]) );
  NOR2X1 U1435 ( .A(n528), .B(n1053), .Y(mem_wdata[82]) );
  NOR2X1 U1436 ( .A(n529), .B(n1051), .Y(mem_wdata[83]) );
  NOR2X1 U1437 ( .A(n530), .B(n1047), .Y(mem_wdata[84]) );
  NOR2X1 U1438 ( .A(n531), .B(n1045), .Y(mem_wdata[85]) );
  NOR2X1 U1439 ( .A(n532), .B(n1050), .Y(mem_wdata[86]) );
  NOR2X1 U1440 ( .A(n533), .B(n1053), .Y(mem_wdata[87]) );
  NOR2X1 U1441 ( .A(n534), .B(n1047), .Y(mem_wdata[88]) );
  NOR2X1 U1442 ( .A(n535), .B(n1047), .Y(mem_wdata[89]) );
  NOR2X1 U1443 ( .A(n536), .B(n1045), .Y(mem_wdata[90]) );
  NOR2X1 U1444 ( .A(n537), .B(n1045), .Y(mem_wdata[91]) );
  NOR2X1 U1445 ( .A(n538), .B(n1048), .Y(mem_wdata[92]) );
  NOR2X1 U1446 ( .A(n539), .B(n1048), .Y(mem_wdata[93]) );
  NOR2X1 U1447 ( .A(n540), .B(n1049), .Y(mem_wdata[94]) );
  NOR2X1 U1448 ( .A(n541), .B(n1046), .Y(mem_wdata[95]) );
  NOR2X1 U1449 ( .A(n556), .B(n1046), .Y(mem_wdata[32]) );
  NOR2X1 U1450 ( .A(n557), .B(n1048), .Y(mem_wdata[33]) );
  NOR2X1 U1451 ( .A(n558), .B(n1176), .Y(mem_wdata[34]) );
  NOR2X1 U1452 ( .A(n559), .B(n1052), .Y(mem_wdata[35]) );
  NOR2X1 U1453 ( .A(n560), .B(n1050), .Y(mem_wdata[36]) );
  NOR2X1 U1454 ( .A(n561), .B(n1045), .Y(mem_wdata[37]) );
  NOR2X1 U1455 ( .A(n562), .B(n1048), .Y(mem_wdata[38]) );
  NOR2X1 U1456 ( .A(n563), .B(n1054), .Y(mem_wdata[39]) );
  NOR2X1 U1457 ( .A(n564), .B(n1049), .Y(mem_wdata[40]) );
  NOR2X1 U1458 ( .A(n565), .B(n1045), .Y(mem_wdata[41]) );
  NOR2X1 U1459 ( .A(n566), .B(n1052), .Y(mem_wdata[42]) );
  NOR2X1 U1460 ( .A(n567), .B(n1052), .Y(mem_wdata[43]) );
  NOR2X1 U1461 ( .A(n568), .B(n1054), .Y(mem_wdata[44]) );
  NOR2X1 U1462 ( .A(n569), .B(n1049), .Y(mem_wdata[45]) );
  NOR2X1 U1463 ( .A(n570), .B(n1176), .Y(mem_wdata[46]) );
  NOR2X1 U1464 ( .A(n571), .B(n1053), .Y(mem_wdata[47]) );
  NOR2X1 U1465 ( .A(n572), .B(n1052), .Y(mem_wdata[48]) );
  NOR2X1 U1466 ( .A(n573), .B(n1047), .Y(mem_wdata[49]) );
  NOR2X1 U1467 ( .A(n574), .B(n1048), .Y(mem_wdata[50]) );
  NOR2X1 U1468 ( .A(n575), .B(n1047), .Y(mem_wdata[51]) );
  NOR2X1 U1469 ( .A(n576), .B(n1047), .Y(mem_wdata[52]) );
  NOR2X1 U1470 ( .A(n577), .B(n1052), .Y(mem_wdata[53]) );
  NOR2X1 U1471 ( .A(n578), .B(n1047), .Y(mem_wdata[54]) );
  NOR2X1 U1472 ( .A(n579), .B(n1045), .Y(mem_wdata[55]) );
  NOR2X1 U1473 ( .A(n580), .B(n1054), .Y(mem_wdata[56]) );
  NOR2X1 U1474 ( .A(n581), .B(n1046), .Y(mem_wdata[57]) );
  NOR2X1 U1475 ( .A(n582), .B(n1053), .Y(mem_wdata[58]) );
  NOR2X1 U1476 ( .A(n583), .B(n1050), .Y(mem_wdata[59]) );
  NOR2X1 U1477 ( .A(n584), .B(n1046), .Y(mem_wdata[60]) );
  NOR2X1 U1478 ( .A(n585), .B(n1049), .Y(mem_wdata[61]) );
  NOR2X1 U1479 ( .A(n586), .B(n1054), .Y(mem_wdata[62]) );
  NOR2X1 U1480 ( .A(n587), .B(n1050), .Y(mem_wdata[63]) );
  NOR2X1 U1481 ( .A(n668), .B(n1054), .Y(mem_wdata[0]) );
  NOR2X1 U1482 ( .A(n671), .B(n1048), .Y(mem_wdata[1]) );
  NOR2X1 U1483 ( .A(n674), .B(n1046), .Y(mem_wdata[2]) );
  NOR2X1 U1484 ( .A(n650), .B(n1047), .Y(mem_wdata[3]) );
  NOR2X1 U1485 ( .A(n653), .B(n1051), .Y(mem_wdata[4]) );
  NOR2X1 U1486 ( .A(n656), .B(n1176), .Y(mem_wdata[5]) );
  NOR2X1 U1487 ( .A(n659), .B(n1051), .Y(mem_wdata[6]) );
  NOR2X1 U1488 ( .A(n662), .B(n1045), .Y(mem_wdata[7]) );
  NOR2X1 U1489 ( .A(n665), .B(n1054), .Y(mem_wdata[8]) );
  NOR2X1 U1490 ( .A(n588), .B(n1176), .Y(mem_wdata[9]) );
  NOR2X1 U1491 ( .A(n589), .B(n1050), .Y(mem_wdata[10]) );
  NOR2X1 U1492 ( .A(n590), .B(n1049), .Y(mem_wdata[11]) );
  NOR2X1 U1493 ( .A(n591), .B(n1046), .Y(mem_wdata[12]) );
  NOR2X1 U1494 ( .A(n592), .B(n1176), .Y(mem_wdata[13]) );
  NOR2X1 U1495 ( .A(n593), .B(n1053), .Y(mem_wdata[14]) );
  NOR2X1 U1496 ( .A(n594), .B(n1176), .Y(mem_wdata[15]) );
  NOR2X1 U1497 ( .A(n595), .B(n1053), .Y(mem_wdata[16]) );
  NOR2X1 U1498 ( .A(n596), .B(n1051), .Y(mem_wdata[17]) );
  NOR2X1 U1499 ( .A(n597), .B(n1176), .Y(mem_wdata[18]) );
  NOR2X1 U1500 ( .A(n598), .B(n1050), .Y(mem_wdata[19]) );
  NOR2X1 U1501 ( .A(n599), .B(n1051), .Y(mem_wdata[20]) );
  NOR2X1 U1502 ( .A(n600), .B(n1051), .Y(mem_wdata[21]) );
  NOR2X1 U1503 ( .A(n601), .B(n1052), .Y(mem_wdata[22]) );
  NOR2X1 U1504 ( .A(n602), .B(n1049), .Y(mem_wdata[23]) );
  NOR2X1 U1505 ( .A(n603), .B(n1051), .Y(mem_wdata[24]) );
  NOR2X1 U1506 ( .A(n604), .B(n1045), .Y(mem_wdata[25]) );
  NOR2X1 U1507 ( .A(n605), .B(n1048), .Y(mem_wdata[26]) );
  NOR2X1 U1508 ( .A(n606), .B(n1176), .Y(mem_wdata[27]) );
  NOR2X1 U1509 ( .A(n607), .B(n1050), .Y(mem_wdata[28]) );
  NOR2X1 U1510 ( .A(n608), .B(n1050), .Y(mem_wdata[29]) );
  NOR2X1 U1511 ( .A(n609), .B(n1054), .Y(mem_wdata[30]) );
  NOR2X1 U1512 ( .A(n610), .B(n1049), .Y(mem_wdata[31]) );
  CLKBUFX3 U1513 ( .A(n11), .Y(n1092) );
  NAND2X1 U1514 ( .A(n470), .B(n1171), .Y(n148) );
  NAND2X1 U1515 ( .A(n469), .B(n1171), .Y(n152) );
  NAND2X1 U1516 ( .A(n468), .B(n1171), .Y(n156) );
  NAND2X1 U1517 ( .A(n467), .B(n1171), .Y(n160) );
  INVX3 U1518 ( .A(n257), .Y(n1175) );
  NOR2X1 U1519 ( .A(n1168), .B(n1170), .Y(n467) );
  NOR2X1 U1520 ( .A(n1257), .B(n1258), .Y(n144) );
  CLKINVX1 U1521 ( .A(tag[4]), .Y(n1207) );
  CLKINVX1 U1522 ( .A(tag[9]), .Y(n1209) );
  CLKINVX1 U1523 ( .A(tag[10]), .Y(n1210) );
  CLKINVX1 U1524 ( .A(tag[11]), .Y(n1211) );
  CLKINVX1 U1525 ( .A(tag[13]), .Y(n1212) );
  CLKINVX1 U1526 ( .A(tag[14]), .Y(n1213) );
  CLKINVX1 U1527 ( .A(tag[15]), .Y(n1214) );
  CLKINVX1 U1528 ( .A(tag[21]), .Y(n1216) );
  CLKINVX1 U1529 ( .A(blockdata[96]), .Y(n1217) );
  CLKINVX1 U1530 ( .A(blockdata[97]), .Y(n1218) );
  CLKINVX1 U1531 ( .A(blockdata[98]), .Y(n1219) );
  CLKINVX1 U1532 ( .A(blockdata[99]), .Y(n1220) );
  CLKINVX1 U1533 ( .A(blockdata[100]), .Y(n1221) );
  CLKINVX1 U1534 ( .A(blockdata[101]), .Y(n1222) );
  CLKINVX1 U1535 ( .A(blockdata[102]), .Y(n1223) );
  CLKINVX1 U1536 ( .A(blockdata[103]), .Y(n1224) );
  CLKINVX1 U1537 ( .A(blockdata[104]), .Y(n1225) );
  CLKINVX1 U1538 ( .A(blockdata[105]), .Y(n1226) );
  CLKINVX1 U1539 ( .A(blockdata[106]), .Y(n1227) );
  CLKINVX1 U1540 ( .A(blockdata[107]), .Y(n1228) );
  CLKINVX1 U1541 ( .A(blockdata[108]), .Y(n1229) );
  CLKINVX1 U1542 ( .A(blockdata[109]), .Y(n1230) );
  CLKINVX1 U1543 ( .A(blockdata[110]), .Y(n1231) );
  CLKINVX1 U1544 ( .A(blockdata[111]), .Y(n1232) );
  CLKINVX1 U1545 ( .A(blockdata[112]), .Y(n1233) );
  CLKINVX1 U1546 ( .A(blockdata[113]), .Y(n1234) );
  CLKINVX1 U1547 ( .A(blockdata[114]), .Y(n1235) );
  CLKINVX1 U1548 ( .A(blockdata[115]), .Y(n1236) );
  CLKINVX1 U1549 ( .A(blockdata[116]), .Y(n1237) );
  CLKINVX1 U1550 ( .A(blockdata[117]), .Y(n1238) );
  CLKINVX1 U1551 ( .A(blockdata[118]), .Y(n1239) );
  CLKINVX1 U1552 ( .A(blockdata[119]), .Y(n1240) );
  CLKINVX1 U1553 ( .A(blockdata[120]), .Y(n1241) );
  CLKINVX1 U1554 ( .A(blockdata[121]), .Y(n1242) );
  CLKINVX1 U1555 ( .A(blockdata[122]), .Y(n1243) );
  CLKINVX1 U1556 ( .A(blockdata[123]), .Y(n1244) );
  CLKINVX1 U1557 ( .A(blockdata[124]), .Y(n1245) );
  CLKINVX1 U1558 ( .A(blockdata[125]), .Y(n1246) );
  CLKINVX1 U1559 ( .A(blockdata[126]), .Y(n1247) );
  CLKINVX1 U1560 ( .A(blockdata[127]), .Y(n1248) );
  CLKBUFX3 U1561 ( .A(N1768), .Y(n1158) );
  CLKBUFX3 U1562 ( .A(N1771), .Y(n1140) );
  CLKBUFX3 U1563 ( .A(N1772), .Y(n1131) );
  CLKBUFX3 U1564 ( .A(N1773), .Y(n1122) );
  CLKBUFX3 U1565 ( .A(N1774), .Y(n1113) );
  CLKBUFX3 U1566 ( .A(N1777), .Y(n1095) );
  OAI222X4 U1567 ( .A0(n1070), .A1(n668), .B0(n508), .B1(n1290), .C0(n1074), 
        .C1(n1418), .Y(block_next[0]) );
  CLKINVX1 U1568 ( .A(mem_rdata[0]), .Y(n1418) );
  OAI222X4 U1569 ( .A0(n1070), .A1(n671), .B0(n508), .B1(n1289), .C0(n1078), 
        .C1(n1417), .Y(block_next[1]) );
  CLKINVX1 U1570 ( .A(mem_rdata[1]), .Y(n1417) );
  OAI222X4 U1571 ( .A0(n1070), .A1(n674), .B0(n1069), .B1(n1288), .C0(n1077), 
        .C1(n1416), .Y(block_next[2]) );
  CLKINVX1 U1572 ( .A(mem_rdata[2]), .Y(n1416) );
  OAI222X4 U1573 ( .A0(n1070), .A1(n650), .B0(n508), .B1(n1287), .C0(n1077), 
        .C1(n1415), .Y(block_next[3]) );
  CLKINVX1 U1574 ( .A(mem_rdata[3]), .Y(n1415) );
  OAI222X4 U1575 ( .A0(n1070), .A1(n653), .B0(n1069), .B1(n1286), .C0(n1076), 
        .C1(n1414), .Y(block_next[4]) );
  CLKINVX1 U1576 ( .A(mem_rdata[4]), .Y(n1414) );
  OAI222X4 U1577 ( .A0(n1070), .A1(n656), .B0(n508), .B1(n1285), .C0(n1075), 
        .C1(n1413), .Y(block_next[5]) );
  CLKINVX1 U1578 ( .A(mem_rdata[5]), .Y(n1413) );
  OAI222X4 U1579 ( .A0(n1070), .A1(n659), .B0(n1069), .B1(n1284), .C0(n1075), 
        .C1(n1412), .Y(block_next[6]) );
  CLKINVX1 U1580 ( .A(mem_rdata[6]), .Y(n1412) );
  OAI222X4 U1581 ( .A0(n1070), .A1(n662), .B0(n508), .B1(n1283), .C0(n1074), 
        .C1(n1411), .Y(block_next[7]) );
  CLKINVX1 U1582 ( .A(mem_rdata[7]), .Y(n1411) );
  OAI222X4 U1583 ( .A0(n1070), .A1(n665), .B0(n1069), .B1(n1282), .C0(n1073), 
        .C1(n1410), .Y(block_next[8]) );
  CLKINVX1 U1584 ( .A(mem_rdata[8]), .Y(n1410) );
  OAI222X4 U1585 ( .A0(n1070), .A1(n588), .B0(n1069), .B1(n1281), .C0(n1073), 
        .C1(n1409), .Y(block_next[9]) );
  CLKINVX1 U1586 ( .A(mem_rdata[9]), .Y(n1409) );
  OAI222X4 U1587 ( .A0(n1070), .A1(n589), .B0(n1069), .B1(n1280), .C0(n1080), 
        .C1(n1408), .Y(block_next[10]) );
  CLKINVX1 U1588 ( .A(mem_rdata[10]), .Y(n1408) );
  OAI222X4 U1589 ( .A0(n1070), .A1(n590), .B0(n508), .B1(n1279), .C0(n1079), 
        .C1(n1407), .Y(block_next[11]) );
  CLKINVX1 U1590 ( .A(mem_rdata[11]), .Y(n1407) );
  OAI222X4 U1591 ( .A0(n1070), .A1(n591), .B0(n1069), .B1(n1278), .C0(n1079), 
        .C1(n1406), .Y(block_next[12]) );
  CLKINVX1 U1592 ( .A(mem_rdata[12]), .Y(n1406) );
  OAI222X4 U1593 ( .A0(n1070), .A1(n592), .B0(n508), .B1(n1277), .C0(n1079), 
        .C1(n1405), .Y(block_next[13]) );
  CLKINVX1 U1594 ( .A(mem_rdata[13]), .Y(n1405) );
  OAI222X4 U1595 ( .A0(n1070), .A1(n593), .B0(n508), .B1(n1276), .C0(n1078), 
        .C1(n1404), .Y(block_next[14]) );
  CLKINVX1 U1596 ( .A(mem_rdata[14]), .Y(n1404) );
  OAI222X4 U1597 ( .A0(n1070), .A1(n594), .B0(n1069), .B1(n1275), .C0(n1078), 
        .C1(n1403), .Y(block_next[15]) );
  CLKINVX1 U1598 ( .A(mem_rdata[15]), .Y(n1403) );
  OAI222X4 U1599 ( .A0(n1070), .A1(n595), .B0(n508), .B1(n1274), .C0(n1078), 
        .C1(n1402), .Y(block_next[16]) );
  CLKINVX1 U1600 ( .A(mem_rdata[16]), .Y(n1402) );
  OAI222X4 U1601 ( .A0(n1070), .A1(n596), .B0(n1069), .B1(n1273), .C0(n1078), 
        .C1(n1401), .Y(block_next[17]) );
  CLKINVX1 U1602 ( .A(mem_rdata[17]), .Y(n1401) );
  OAI222X4 U1603 ( .A0(n1070), .A1(n597), .B0(n1069), .B1(n1272), .C0(n1078), 
        .C1(n1400), .Y(block_next[18]) );
  CLKINVX1 U1604 ( .A(mem_rdata[18]), .Y(n1400) );
  OAI222X4 U1605 ( .A0(n1070), .A1(n598), .B0(n508), .B1(n1271), .C0(n1078), 
        .C1(n1399), .Y(block_next[19]) );
  CLKINVX1 U1606 ( .A(mem_rdata[19]), .Y(n1399) );
  OAI222X4 U1607 ( .A0(n1070), .A1(n599), .B0(n508), .B1(n1270), .C0(n1078), 
        .C1(n1398), .Y(block_next[20]) );
  CLKINVX1 U1608 ( .A(mem_rdata[20]), .Y(n1398) );
  OAI222X4 U1609 ( .A0(n1070), .A1(n600), .B0(n1069), .B1(n1269), .C0(n1078), 
        .C1(n1397), .Y(block_next[21]) );
  CLKINVX1 U1610 ( .A(mem_rdata[21]), .Y(n1397) );
  OAI222X4 U1611 ( .A0(n1070), .A1(n601), .B0(n1069), .B1(n1268), .C0(n1078), 
        .C1(n1396), .Y(block_next[22]) );
  CLKINVX1 U1612 ( .A(mem_rdata[22]), .Y(n1396) );
  OAI222X4 U1613 ( .A0(n1070), .A1(n602), .B0(n508), .B1(n1267), .C0(n1078), 
        .C1(n1395), .Y(block_next[23]) );
  CLKINVX1 U1614 ( .A(mem_rdata[23]), .Y(n1395) );
  OAI222X4 U1615 ( .A0(n1070), .A1(n603), .B0(n1069), .B1(n1266), .C0(n1078), 
        .C1(n1394), .Y(block_next[24]) );
  CLKINVX1 U1616 ( .A(mem_rdata[24]), .Y(n1394) );
  OAI222X4 U1617 ( .A0(n1070), .A1(n604), .B0(n508), .B1(n1265), .C0(n1078), 
        .C1(n1393), .Y(block_next[25]) );
  CLKINVX1 U1618 ( .A(mem_rdata[25]), .Y(n1393) );
  OAI222X4 U1619 ( .A0(n1070), .A1(n605), .B0(n508), .B1(n1264), .C0(n1078), 
        .C1(n1392), .Y(block_next[26]) );
  CLKINVX1 U1620 ( .A(mem_rdata[26]), .Y(n1392) );
  OAI222X4 U1621 ( .A0(n1070), .A1(n606), .B0(n1069), .B1(n1263), .C0(n1078), 
        .C1(n1391), .Y(block_next[27]) );
  CLKINVX1 U1622 ( .A(mem_rdata[27]), .Y(n1391) );
  OAI222X4 U1623 ( .A0(n1070), .A1(n607), .B0(n508), .B1(n1262), .C0(n1078), 
        .C1(n1390), .Y(block_next[28]) );
  CLKINVX1 U1624 ( .A(mem_rdata[28]), .Y(n1390) );
  OAI222X4 U1625 ( .A0(n1070), .A1(n608), .B0(n1069), .B1(n1261), .C0(n1077), 
        .C1(n1389), .Y(block_next[29]) );
  CLKINVX1 U1626 ( .A(mem_rdata[29]), .Y(n1389) );
  OAI222X4 U1627 ( .A0(n1070), .A1(n609), .B0(n508), .B1(n1260), .C0(n1077), 
        .C1(n1388), .Y(block_next[30]) );
  CLKINVX1 U1628 ( .A(mem_rdata[30]), .Y(n1388) );
  OAI222X4 U1629 ( .A0(n1070), .A1(n610), .B0(n1069), .B1(n1259), .C0(n1077), 
        .C1(n1387), .Y(block_next[31]) );
  CLKINVX1 U1630 ( .A(mem_rdata[31]), .Y(n1387) );
  OAI222X4 U1631 ( .A0(n1057), .A1(n556), .B0(n1290), .B1(n1058), .C0(n1077), 
        .C1(n1386), .Y(block_next[32]) );
  CLKINVX1 U1632 ( .A(mem_rdata[32]), .Y(n1386) );
  OAI222X4 U1633 ( .A0(n1057), .A1(n557), .B0(n1289), .B1(n1058), .C0(n1077), 
        .C1(n1385), .Y(block_next[33]) );
  CLKINVX1 U1634 ( .A(mem_rdata[33]), .Y(n1385) );
  OAI222X4 U1635 ( .A0(n1057), .A1(n558), .B0(n1288), .B1(n1058), .C0(n1077), 
        .C1(n1384), .Y(block_next[34]) );
  CLKINVX1 U1636 ( .A(mem_rdata[34]), .Y(n1384) );
  OAI222X4 U1637 ( .A0(n1057), .A1(n559), .B0(n1287), .B1(n1058), .C0(n1077), 
        .C1(n1383), .Y(block_next[35]) );
  CLKINVX1 U1638 ( .A(mem_rdata[35]), .Y(n1383) );
  OAI222X4 U1639 ( .A0(n1057), .A1(n560), .B0(n1286), .B1(n1058), .C0(n1077), 
        .C1(n1382), .Y(block_next[36]) );
  CLKINVX1 U1640 ( .A(mem_rdata[36]), .Y(n1382) );
  OAI222X4 U1641 ( .A0(n1057), .A1(n561), .B0(n1285), .B1(n1058), .C0(n1077), 
        .C1(n1381), .Y(block_next[37]) );
  CLKINVX1 U1642 ( .A(mem_rdata[37]), .Y(n1381) );
  OAI222X4 U1643 ( .A0(n1057), .A1(n562), .B0(n1284), .B1(n1059), .C0(n1077), 
        .C1(n1380), .Y(block_next[38]) );
  CLKINVX1 U1644 ( .A(mem_rdata[38]), .Y(n1380) );
  OAI222X4 U1645 ( .A0(n1057), .A1(n563), .B0(n1283), .B1(n1058), .C0(n1077), 
        .C1(n1379), .Y(block_next[39]) );
  CLKINVX1 U1646 ( .A(mem_rdata[39]), .Y(n1379) );
  OAI222X4 U1647 ( .A0(n1056), .A1(n564), .B0(n1282), .B1(n1058), .C0(n1077), 
        .C1(n1378), .Y(block_next[40]) );
  CLKINVX1 U1648 ( .A(mem_rdata[40]), .Y(n1378) );
  OAI222X4 U1649 ( .A0(n1056), .A1(n565), .B0(n1281), .B1(n1058), .C0(n1077), 
        .C1(n1377), .Y(block_next[41]) );
  CLKINVX1 U1650 ( .A(mem_rdata[41]), .Y(n1377) );
  OAI222X4 U1651 ( .A0(n1056), .A1(n566), .B0(n1280), .B1(n1058), .C0(n1077), 
        .C1(n1376), .Y(block_next[42]) );
  CLKINVX1 U1652 ( .A(mem_rdata[42]), .Y(n1376) );
  OAI222X4 U1653 ( .A0(n1056), .A1(n567), .B0(n1279), .B1(n1058), .C0(n1076), 
        .C1(n1375), .Y(block_next[43]) );
  CLKINVX1 U1654 ( .A(mem_rdata[43]), .Y(n1375) );
  OAI222X4 U1655 ( .A0(n1056), .A1(n568), .B0(n1278), .B1(n1058), .C0(n1076), 
        .C1(n1374), .Y(block_next[44]) );
  CLKINVX1 U1656 ( .A(mem_rdata[44]), .Y(n1374) );
  OAI222X4 U1657 ( .A0(n1056), .A1(n569), .B0(n1277), .B1(n1059), .C0(n1076), 
        .C1(n1373), .Y(block_next[45]) );
  CLKINVX1 U1658 ( .A(mem_rdata[45]), .Y(n1373) );
  OAI222X4 U1659 ( .A0(n1056), .A1(n570), .B0(n1276), .B1(n1059), .C0(n1076), 
        .C1(n1372), .Y(block_next[46]) );
  CLKINVX1 U1660 ( .A(mem_rdata[46]), .Y(n1372) );
  OAI222X4 U1661 ( .A0(n1056), .A1(n571), .B0(n1275), .B1(n1059), .C0(n1076), 
        .C1(n1371), .Y(block_next[47]) );
  CLKINVX1 U1662 ( .A(mem_rdata[47]), .Y(n1371) );
  OAI222X4 U1663 ( .A0(n1056), .A1(n572), .B0(n1274), .B1(n1059), .C0(n1076), 
        .C1(n1370), .Y(block_next[48]) );
  CLKINVX1 U1664 ( .A(mem_rdata[48]), .Y(n1370) );
  OAI222X4 U1665 ( .A0(n1056), .A1(n573), .B0(n1273), .B1(n1059), .C0(n1076), 
        .C1(n1369), .Y(block_next[49]) );
  CLKINVX1 U1666 ( .A(mem_rdata[49]), .Y(n1369) );
  OAI222X4 U1667 ( .A0(n1056), .A1(n574), .B0(n1272), .B1(n1059), .C0(n1076), 
        .C1(n1368), .Y(block_next[50]) );
  CLKINVX1 U1668 ( .A(mem_rdata[50]), .Y(n1368) );
  OAI222X4 U1669 ( .A0(n1056), .A1(n575), .B0(n1271), .B1(n1059), .C0(n1076), 
        .C1(n1367), .Y(block_next[51]) );
  CLKINVX1 U1670 ( .A(mem_rdata[51]), .Y(n1367) );
  OAI222X4 U1671 ( .A0(n1055), .A1(n576), .B0(n1270), .B1(n1059), .C0(n1076), 
        .C1(n1366), .Y(block_next[52]) );
  CLKINVX1 U1672 ( .A(mem_rdata[52]), .Y(n1366) );
  OAI222X4 U1673 ( .A0(n1055), .A1(n577), .B0(n1269), .B1(n1059), .C0(n1076), 
        .C1(n1365), .Y(block_next[53]) );
  CLKINVX1 U1674 ( .A(mem_rdata[53]), .Y(n1365) );
  OAI222X4 U1675 ( .A0(n1055), .A1(n578), .B0(n1268), .B1(n1059), .C0(n1076), 
        .C1(n1364), .Y(block_next[54]) );
  CLKINVX1 U1676 ( .A(mem_rdata[54]), .Y(n1364) );
  OAI222X4 U1677 ( .A0(n1055), .A1(n579), .B0(n1267), .B1(n1059), .C0(n1076), 
        .C1(n1363), .Y(block_next[55]) );
  CLKINVX1 U1678 ( .A(mem_rdata[55]), .Y(n1363) );
  OAI222X4 U1679 ( .A0(n1055), .A1(n580), .B0(n1266), .B1(n1058), .C0(n1076), 
        .C1(n1362), .Y(block_next[56]) );
  CLKINVX1 U1680 ( .A(mem_rdata[56]), .Y(n1362) );
  OAI222X4 U1681 ( .A0(n1055), .A1(n581), .B0(n1265), .B1(n1059), .C0(n1076), 
        .C1(n1361), .Y(block_next[57]) );
  CLKINVX1 U1682 ( .A(mem_rdata[57]), .Y(n1361) );
  OAI222X4 U1683 ( .A0(n1055), .A1(n582), .B0(n1264), .B1(n1058), .C0(n1075), 
        .C1(n1360), .Y(block_next[58]) );
  CLKINVX1 U1684 ( .A(mem_rdata[58]), .Y(n1360) );
  OAI222X4 U1685 ( .A0(n1055), .A1(n583), .B0(n1263), .B1(n1059), .C0(n1075), 
        .C1(n1359), .Y(block_next[59]) );
  CLKINVX1 U1686 ( .A(mem_rdata[59]), .Y(n1359) );
  OAI222X4 U1687 ( .A0(n1055), .A1(n584), .B0(n1262), .B1(n1058), .C0(n1075), 
        .C1(n1358), .Y(block_next[60]) );
  CLKINVX1 U1688 ( .A(mem_rdata[60]), .Y(n1358) );
  OAI222X4 U1689 ( .A0(n1055), .A1(n585), .B0(n1261), .B1(n1059), .C0(n1075), 
        .C1(n1357), .Y(block_next[61]) );
  CLKINVX1 U1690 ( .A(mem_rdata[61]), .Y(n1357) );
  OAI222X4 U1691 ( .A0(n1055), .A1(n586), .B0(n1260), .B1(n1058), .C0(n1075), 
        .C1(n1356), .Y(block_next[62]) );
  CLKINVX1 U1692 ( .A(mem_rdata[62]), .Y(n1356) );
  OAI222X4 U1693 ( .A0(n1055), .A1(n587), .B0(n1259), .B1(n1059), .C0(n1075), 
        .C1(n1355), .Y(block_next[63]) );
  CLKINVX1 U1694 ( .A(mem_rdata[63]), .Y(n1355) );
  OAI222X4 U1695 ( .A0(n1064), .A1(n510), .B0(n1290), .B1(n1060), .C0(n1075), 
        .C1(n1354), .Y(block_next[64]) );
  CLKINVX1 U1696 ( .A(mem_rdata[64]), .Y(n1354) );
  OAI222X4 U1697 ( .A0(n1064), .A1(n511), .B0(n1289), .B1(n1060), .C0(n1075), 
        .C1(n1353), .Y(block_next[65]) );
  CLKINVX1 U1698 ( .A(mem_rdata[65]), .Y(n1353) );
  OAI222X4 U1699 ( .A0(n1064), .A1(n512), .B0(n1288), .B1(n1060), .C0(n1075), 
        .C1(n1352), .Y(block_next[66]) );
  CLKINVX1 U1700 ( .A(mem_rdata[66]), .Y(n1352) );
  OAI222X4 U1701 ( .A0(n1064), .A1(n513), .B0(n1287), .B1(n1060), .C0(n1075), 
        .C1(n1351), .Y(block_next[67]) );
  CLKINVX1 U1702 ( .A(mem_rdata[67]), .Y(n1351) );
  OAI222X4 U1703 ( .A0(n1064), .A1(n514), .B0(n1060), .B1(n1286), .C0(n1075), 
        .C1(n1350), .Y(block_next[68]) );
  CLKINVX1 U1704 ( .A(mem_rdata[68]), .Y(n1350) );
  OAI222X4 U1705 ( .A0(n1064), .A1(n515), .B0(n1061), .B1(n1285), .C0(n1075), 
        .C1(n1349), .Y(block_next[69]) );
  CLKINVX1 U1706 ( .A(mem_rdata[69]), .Y(n1349) );
  OAI222X4 U1707 ( .A0(n1064), .A1(n516), .B0(n1060), .B1(n1284), .C0(n1075), 
        .C1(n1348), .Y(block_next[70]) );
  CLKINVX1 U1708 ( .A(mem_rdata[70]), .Y(n1348) );
  OAI222X4 U1709 ( .A0(n1064), .A1(n517), .B0(n1060), .B1(n1283), .C0(n1075), 
        .C1(n1347), .Y(block_next[71]) );
  CLKINVX1 U1710 ( .A(mem_rdata[71]), .Y(n1347) );
  OAI222X4 U1711 ( .A0(n1063), .A1(n518), .B0(n1060), .B1(n1282), .C0(n1074), 
        .C1(n1346), .Y(block_next[72]) );
  CLKINVX1 U1712 ( .A(mem_rdata[72]), .Y(n1346) );
  OAI222X4 U1713 ( .A0(n1063), .A1(n519), .B0(n1281), .B1(n1060), .C0(n1074), 
        .C1(n1345), .Y(block_next[73]) );
  CLKINVX1 U1714 ( .A(mem_rdata[73]), .Y(n1345) );
  OAI222X4 U1715 ( .A0(n1063), .A1(n520), .B0(n1060), .B1(n1280), .C0(n1074), 
        .C1(n1344), .Y(block_next[74]) );
  CLKINVX1 U1716 ( .A(mem_rdata[74]), .Y(n1344) );
  OAI222X4 U1717 ( .A0(n1063), .A1(n521), .B0(n1060), .B1(n1279), .C0(n1074), 
        .C1(n1343), .Y(block_next[75]) );
  CLKINVX1 U1718 ( .A(mem_rdata[75]), .Y(n1343) );
  OAI222X4 U1719 ( .A0(n1063), .A1(n522), .B0(n1060), .B1(n1278), .C0(n1074), 
        .C1(n1342), .Y(block_next[76]) );
  CLKINVX1 U1720 ( .A(mem_rdata[76]), .Y(n1342) );
  OAI222X4 U1721 ( .A0(n1063), .A1(n523), .B0(n1061), .B1(n1277), .C0(n1074), 
        .C1(n1341), .Y(block_next[77]) );
  CLKINVX1 U1722 ( .A(mem_rdata[77]), .Y(n1341) );
  OAI222X4 U1723 ( .A0(n1063), .A1(n524), .B0(n1061), .B1(n1276), .C0(n1074), 
        .C1(n1340), .Y(block_next[78]) );
  CLKINVX1 U1724 ( .A(mem_rdata[78]), .Y(n1340) );
  OAI222X4 U1725 ( .A0(n1063), .A1(n525), .B0(n1061), .B1(n1275), .C0(n1074), 
        .C1(n1339), .Y(block_next[79]) );
  CLKINVX1 U1726 ( .A(mem_rdata[79]), .Y(n1339) );
  OAI222X4 U1727 ( .A0(n1063), .A1(n526), .B0(n1061), .B1(n1274), .C0(n1074), 
        .C1(n1338), .Y(block_next[80]) );
  CLKINVX1 U1728 ( .A(mem_rdata[80]), .Y(n1338) );
  OAI222X4 U1729 ( .A0(n1063), .A1(n527), .B0(n1061), .B1(n1273), .C0(n1074), 
        .C1(n1337), .Y(block_next[81]) );
  CLKINVX1 U1730 ( .A(mem_rdata[81]), .Y(n1337) );
  OAI222X4 U1731 ( .A0(n1063), .A1(n528), .B0(n1061), .B1(n1272), .C0(n1074), 
        .C1(n1336), .Y(block_next[82]) );
  CLKINVX1 U1732 ( .A(mem_rdata[82]), .Y(n1336) );
  OAI222X4 U1733 ( .A0(n1063), .A1(n529), .B0(n1061), .B1(n1271), .C0(n1074), 
        .C1(n1335), .Y(block_next[83]) );
  CLKINVX1 U1734 ( .A(mem_rdata[83]), .Y(n1335) );
  OAI222X4 U1735 ( .A0(n1062), .A1(n530), .B0(n1061), .B1(n1270), .C0(n1074), 
        .C1(n1334), .Y(block_next[84]) );
  CLKINVX1 U1736 ( .A(mem_rdata[84]), .Y(n1334) );
  OAI222X4 U1737 ( .A0(n1062), .A1(n531), .B0(n1061), .B1(n1269), .C0(n1074), 
        .C1(n1333), .Y(block_next[85]) );
  CLKINVX1 U1738 ( .A(mem_rdata[85]), .Y(n1333) );
  OAI222X4 U1739 ( .A0(n1062), .A1(n532), .B0(n1061), .B1(n1268), .C0(n1074), 
        .C1(n1332), .Y(block_next[86]) );
  CLKINVX1 U1740 ( .A(mem_rdata[86]), .Y(n1332) );
  OAI222X4 U1741 ( .A0(n1062), .A1(n533), .B0(n1061), .B1(n1267), .C0(n1073), 
        .C1(n1331), .Y(block_next[87]) );
  CLKINVX1 U1742 ( .A(mem_rdata[87]), .Y(n1331) );
  OAI222X4 U1743 ( .A0(n1062), .A1(n534), .B0(n1061), .B1(n1266), .C0(n1073), 
        .C1(n1330), .Y(block_next[88]) );
  CLKINVX1 U1744 ( .A(mem_rdata[88]), .Y(n1330) );
  OAI222X4 U1745 ( .A0(n1062), .A1(n535), .B0(n1061), .B1(n1265), .C0(n1073), 
        .C1(n1329), .Y(block_next[89]) );
  CLKINVX1 U1746 ( .A(mem_rdata[89]), .Y(n1329) );
  OAI222X4 U1747 ( .A0(n1062), .A1(n536), .B0(n1060), .B1(n1264), .C0(n1073), 
        .C1(n1328), .Y(block_next[90]) );
  CLKINVX1 U1748 ( .A(mem_rdata[90]), .Y(n1328) );
  OAI222X4 U1749 ( .A0(n1062), .A1(n537), .B0(n1061), .B1(n1263), .C0(n1073), 
        .C1(n1327), .Y(block_next[91]) );
  CLKINVX1 U1750 ( .A(mem_rdata[91]), .Y(n1327) );
  OAI222X4 U1751 ( .A0(n1062), .A1(n538), .B0(n1060), .B1(n1262), .C0(n1073), 
        .C1(n1326), .Y(block_next[92]) );
  CLKINVX1 U1752 ( .A(mem_rdata[92]), .Y(n1326) );
  OAI222X4 U1753 ( .A0(n1062), .A1(n539), .B0(n1061), .B1(n1261), .C0(n1073), 
        .C1(n1325), .Y(block_next[93]) );
  CLKINVX1 U1754 ( .A(mem_rdata[93]), .Y(n1325) );
  OAI222X4 U1755 ( .A0(n1062), .A1(n540), .B0(n1060), .B1(n1260), .C0(n1073), 
        .C1(n1324), .Y(block_next[94]) );
  CLKINVX1 U1756 ( .A(mem_rdata[94]), .Y(n1324) );
  OAI222X4 U1757 ( .A0(n1062), .A1(n541), .B0(n1060), .B1(n1259), .C0(n1073), 
        .C1(n1323), .Y(block_next[95]) );
  CLKINVX1 U1758 ( .A(mem_rdata[95]), .Y(n1323) );
  OAI222X4 U1759 ( .A0(n1067), .A1(n1217), .B0(n1066), .B1(n1290), .C0(n1073), 
        .C1(n1322), .Y(block_next[96]) );
  CLKINVX1 U1760 ( .A(mem_rdata[96]), .Y(n1322) );
  OAI222X4 U1761 ( .A0(n1067), .A1(n1218), .B0(n1065), .B1(n1289), .C0(n1073), 
        .C1(n1321), .Y(block_next[97]) );
  CLKINVX1 U1762 ( .A(mem_rdata[97]), .Y(n1321) );
  OAI222X4 U1763 ( .A0(n1067), .A1(n1219), .B0(n1066), .B1(n1288), .C0(n1073), 
        .C1(n1320), .Y(block_next[98]) );
  CLKINVX1 U1764 ( .A(mem_rdata[98]), .Y(n1320) );
  OAI222X4 U1765 ( .A0(n1067), .A1(n1220), .B0(n1065), .B1(n1287), .C0(n1073), 
        .C1(n1319), .Y(block_next[99]) );
  CLKINVX1 U1766 ( .A(mem_rdata[99]), .Y(n1319) );
  OAI222X4 U1767 ( .A0(n266), .A1(n1221), .B0(n1065), .B1(n1286), .C0(n1080), 
        .C1(n1318), .Y(block_next[100]) );
  CLKINVX1 U1768 ( .A(mem_rdata[100]), .Y(n1318) );
  OAI222X4 U1769 ( .A0(n266), .A1(n1222), .B0(n1065), .B1(n1285), .C0(n1080), 
        .C1(n1317), .Y(block_next[101]) );
  CLKINVX1 U1770 ( .A(mem_rdata[101]), .Y(n1317) );
  OAI222X4 U1771 ( .A0(n266), .A1(n1223), .B0(n1065), .B1(n1284), .C0(n1080), 
        .C1(n1316), .Y(block_next[102]) );
  CLKINVX1 U1772 ( .A(mem_rdata[102]), .Y(n1316) );
  OAI222X4 U1773 ( .A0(n266), .A1(n1224), .B0(n1065), .B1(n1283), .C0(n1080), 
        .C1(n1315), .Y(block_next[103]) );
  CLKINVX1 U1774 ( .A(mem_rdata[103]), .Y(n1315) );
  OAI222X4 U1775 ( .A0(n266), .A1(n1225), .B0(n1065), .B1(n1282), .C0(n1080), 
        .C1(n1314), .Y(block_next[104]) );
  CLKINVX1 U1776 ( .A(mem_rdata[104]), .Y(n1314) );
  OAI222X4 U1777 ( .A0(n266), .A1(n1226), .B0(n1281), .B1(n1065), .C0(n1080), 
        .C1(n1313), .Y(block_next[105]) );
  CLKINVX1 U1778 ( .A(mem_rdata[105]), .Y(n1313) );
  OAI222X4 U1779 ( .A0(n266), .A1(n1227), .B0(n1065), .B1(n1280), .C0(n1080), 
        .C1(n1312), .Y(block_next[106]) );
  CLKINVX1 U1780 ( .A(mem_rdata[106]), .Y(n1312) );
  OAI222X4 U1781 ( .A0(n266), .A1(n1228), .B0(n1066), .B1(n1279), .C0(n1080), 
        .C1(n1311), .Y(block_next[107]) );
  CLKINVX1 U1782 ( .A(mem_rdata[107]), .Y(n1311) );
  OAI222X4 U1783 ( .A0(n1068), .A1(n1229), .B0(n1065), .B1(n1278), .C0(n1080), 
        .C1(n1310), .Y(block_next[108]) );
  CLKINVX1 U1784 ( .A(mem_rdata[108]), .Y(n1310) );
  OAI222X4 U1785 ( .A0(n1068), .A1(n1230), .B0(n1065), .B1(n1277), .C0(n1080), 
        .C1(n1309), .Y(block_next[109]) );
  CLKINVX1 U1786 ( .A(mem_rdata[109]), .Y(n1309) );
  OAI222X4 U1787 ( .A0(n1068), .A1(n1231), .B0(n1065), .B1(n1276), .C0(n1080), 
        .C1(n1308), .Y(block_next[110]) );
  CLKINVX1 U1788 ( .A(mem_rdata[110]), .Y(n1308) );
  OAI222X4 U1789 ( .A0(n1068), .A1(n1232), .B0(n1065), .B1(n1275), .C0(n1080), 
        .C1(n1307), .Y(block_next[111]) );
  CLKINVX1 U1790 ( .A(mem_rdata[111]), .Y(n1307) );
  OAI222X4 U1791 ( .A0(n1068), .A1(n1233), .B0(n1065), .B1(n1274), .C0(n1080), 
        .C1(n1306), .Y(block_next[112]) );
  CLKINVX1 U1792 ( .A(mem_rdata[112]), .Y(n1306) );
  OAI222X4 U1793 ( .A0(n1068), .A1(n1234), .B0(n1066), .B1(n1273), .C0(n1080), 
        .C1(n1305), .Y(block_next[113]) );
  CLKINVX1 U1794 ( .A(mem_rdata[113]), .Y(n1305) );
  OAI222X4 U1795 ( .A0(n1068), .A1(n1235), .B0(n1066), .B1(n1272), .C0(n1080), 
        .C1(n1304), .Y(block_next[114]) );
  CLKINVX1 U1796 ( .A(mem_rdata[114]), .Y(n1304) );
  OAI222X4 U1797 ( .A0(n1068), .A1(n1236), .B0(n1066), .B1(n1271), .C0(n1079), 
        .C1(n1303), .Y(block_next[115]) );
  CLKINVX1 U1798 ( .A(mem_rdata[115]), .Y(n1303) );
  OAI222X4 U1799 ( .A0(n1068), .A1(n1237), .B0(n1066), .B1(n1270), .C0(n1079), 
        .C1(n1302), .Y(block_next[116]) );
  CLKINVX1 U1800 ( .A(mem_rdata[116]), .Y(n1302) );
  OAI222X4 U1801 ( .A0(n1068), .A1(n1238), .B0(n1066), .B1(n1269), .C0(n1079), 
        .C1(n1301), .Y(block_next[117]) );
  CLKINVX1 U1802 ( .A(mem_rdata[117]), .Y(n1301) );
  OAI222X4 U1803 ( .A0(n1068), .A1(n1239), .B0(n1066), .B1(n1268), .C0(n1079), 
        .C1(n1300), .Y(block_next[118]) );
  CLKINVX1 U1804 ( .A(mem_rdata[118]), .Y(n1300) );
  OAI222X4 U1805 ( .A0(n1068), .A1(n1240), .B0(n1066), .B1(n1267), .C0(n1079), 
        .C1(n1299), .Y(block_next[119]) );
  CLKINVX1 U1806 ( .A(mem_rdata[119]), .Y(n1299) );
  OAI222X4 U1807 ( .A0(n1067), .A1(n1241), .B0(n1066), .B1(n1266), .C0(n1079), 
        .C1(n1298), .Y(block_next[120]) );
  CLKINVX1 U1808 ( .A(mem_rdata[120]), .Y(n1298) );
  OAI222X4 U1809 ( .A0(n1067), .A1(n1242), .B0(n1066), .B1(n1265), .C0(n1079), 
        .C1(n1297), .Y(block_next[121]) );
  CLKINVX1 U1810 ( .A(mem_rdata[121]), .Y(n1297) );
  OAI222X4 U1811 ( .A0(n1067), .A1(n1243), .B0(n1066), .B1(n1264), .C0(n1079), 
        .C1(n1296), .Y(block_next[122]) );
  CLKINVX1 U1812 ( .A(mem_rdata[122]), .Y(n1296) );
  OAI222X4 U1813 ( .A0(n1067), .A1(n1244), .B0(n1066), .B1(n1263), .C0(n1079), 
        .C1(n1295), .Y(block_next[123]) );
  CLKINVX1 U1814 ( .A(mem_rdata[123]), .Y(n1295) );
  OAI222X4 U1815 ( .A0(n1067), .A1(n1245), .B0(n1066), .B1(n1262), .C0(n1079), 
        .C1(n1294), .Y(block_next[124]) );
  CLKINVX1 U1816 ( .A(mem_rdata[124]), .Y(n1294) );
  OAI222X4 U1817 ( .A0(n1067), .A1(n1246), .B0(n1065), .B1(n1261), .C0(n1079), 
        .C1(n1293), .Y(block_next[125]) );
  CLKINVX1 U1818 ( .A(mem_rdata[125]), .Y(n1293) );
  OAI222X4 U1819 ( .A0(n1067), .A1(n1247), .B0(n1066), .B1(n1260), .C0(n1079), 
        .C1(n1292), .Y(block_next[126]) );
  CLKINVX1 U1820 ( .A(mem_rdata[126]), .Y(n1292) );
  OAI222X4 U1821 ( .A0(n1067), .A1(n1248), .B0(n1065), .B1(n1259), .C0(n1079), 
        .C1(n1291), .Y(block_next[127]) );
  CLKINVX1 U1822 ( .A(mem_rdata[127]), .Y(n1291) );
  OAI222X1 U1823 ( .A0(n613), .A1(valid), .B0(n1174), .B1(n145), .C0(n261), 
        .C1(n256), .Y(n431) );
  MXI2X1 U1824 ( .A(n968), .B(n969), .S0(n1044), .Y(tag[0]) );
  MXI4X1 U1825 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(
        \blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n999), .S1(n1028), .Y(
        n968) );
  MXI2X1 U1826 ( .A(n966), .B(n967), .S0(n1044), .Y(tag[1]) );
  MXI4X1 U1827 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(
        \blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n999), .S1(n1028), .Y(
        n966) );
  MXI4X1 U1828 ( .A(\blocktag[4][1] ), .B(\blocktag[5][1] ), .C(
        \blocktag[6][1] ), .D(\blocktag[7][1] ), .S0(n999), .S1(n1028), .Y(
        n967) );
  MXI2X1 U1829 ( .A(n962), .B(n963), .S0(n1044), .Y(tag[3]) );
  MXI4X1 U1830 ( .A(\blocktag[0][3] ), .B(\blocktag[1][3] ), .C(
        \blocktag[2][3] ), .D(\blocktag[3][3] ), .S0(n999), .S1(n1028), .Y(
        n962) );
  MXI4X1 U1831 ( .A(\blocktag[4][3] ), .B(\blocktag[5][3] ), .C(
        \blocktag[6][3] ), .D(\blocktag[7][3] ), .S0(n677), .S1(n1028), .Y(
        n963) );
  MXI2X1 U1832 ( .A(n928), .B(n929), .S0(n1043), .Y(tag[20]) );
  MXI4X1 U1833 ( .A(\blocktag[0][20] ), .B(\blocktag[1][20] ), .C(
        \blocktag[2][20] ), .D(\blocktag[3][20] ), .S0(n996), .S1(n1031), .Y(
        n928) );
  MXI4X1 U1834 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n677), .S1(n1030), .Y(
        n929) );
  MXI2X1 U1835 ( .A(n960), .B(n961), .S0(n1044), .Y(tag[4]) );
  MXI4X1 U1836 ( .A(\blocktag[0][4] ), .B(\blocktag[1][4] ), .C(
        \blocktag[2][4] ), .D(\blocktag[3][4] ), .S0(n999), .S1(n1028), .Y(
        n960) );
  MXI4X1 U1837 ( .A(\blocktag[4][4] ), .B(\blocktag[5][4] ), .C(
        \blocktag[6][4] ), .D(\blocktag[7][4] ), .S0(n999), .S1(n1028), .Y(
        n961) );
  MXI2X1 U1838 ( .A(n942), .B(n943), .S0(n1043), .Y(tag[13]) );
  MXI4X1 U1839 ( .A(\blocktag[0][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[3][13] ), .S0(n997), .S1(n1031), .Y(
        n942) );
  MXI4X1 U1840 ( .A(\blocktag[4][13] ), .B(\blocktag[5][13] ), .C(
        \blocktag[6][13] ), .D(\blocktag[7][13] ), .S0(n997), .S1(n1030), .Y(
        n943) );
  MXI2X1 U1841 ( .A(n940), .B(n941), .S0(n1043), .Y(tag[14]) );
  MXI4X1 U1842 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n997), .S1(n1169), .Y(
        n940) );
  MXI4X1 U1843 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n997), .S1(n1169), .Y(
        n941) );
  MXI2X1 U1844 ( .A(n938), .B(n939), .S0(n1043), .Y(tag[15]) );
  MXI4X1 U1845 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n997), .S1(n1002), .Y(
        n938) );
  MXI4X1 U1846 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n997), .S1(n1002), .Y(
        n939) );
  MXI2X1 U1847 ( .A(n950), .B(n951), .S0(n1044), .Y(tag[9]) );
  MXI4X1 U1848 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(
        \blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n998), .S1(n1002), .Y(
        n950) );
  MXI4X1 U1849 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(
        \blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n998), .S1(n1002), .Y(
        n951) );
  MXI2X1 U1850 ( .A(n948), .B(n949), .S0(n1044), .Y(tag[10]) );
  MXI4X1 U1851 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n998), .S1(n1002), .Y(
        n948) );
  MXI4X1 U1852 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n998), .S1(n1031), .Y(
        n949) );
  MXI2X1 U1853 ( .A(n926), .B(n927), .S0(n1043), .Y(tag[21]) );
  MXI2X1 U1854 ( .A(n946), .B(n947), .S0(n1044), .Y(tag[11]) );
  MXI4X1 U1855 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n998), .S1(n1030), .Y(
        n946) );
  MXI4X1 U1856 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n998), .S1(n1031), .Y(
        n947) );
  XNOR2X1 U1857 ( .A(proc_addr[5]), .B(tag[0]), .Y(n445) );
  NOR4X1 U1858 ( .A(n438), .B(n439), .C(n440), .D(n441), .Y(n437) );
  XNOR2X1 U1859 ( .A(n551), .B(proc_addr[28]), .Y(n439) );
  XNOR2X1 U1860 ( .A(n552), .B(proc_addr[17]), .Y(n440) );
  XNOR2X1 U1861 ( .A(n553), .B(proc_addr[27]), .Y(n441) );
  MXI4X1 U1862 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(
        \blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n999), .S1(n1028), .Y(
        n964) );
  MXI4X1 U1863 ( .A(\blocktag[4][2] ), .B(\blocktag[5][2] ), .C(
        \blocktag[6][2] ), .D(\blocktag[7][2] ), .S0(n999), .S1(n1028), .Y(
        n965) );
  MXI4X1 U1864 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(
        \blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n999), .S1(n1028), .Y(
        n958) );
  MXI4X1 U1865 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(
        \blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n999), .S1(n1028), .Y(
        n959) );
  MXI4X1 U1866 ( .A(\blocktag[0][6] ), .B(\blocktag[1][6] ), .C(
        \blocktag[2][6] ), .D(\blocktag[3][6] ), .S0(n999), .S1(n1030), .Y(
        n956) );
  MXI4X1 U1867 ( .A(\blocktag[4][6] ), .B(\blocktag[5][6] ), .C(
        \blocktag[6][6] ), .D(\blocktag[7][6] ), .S0(n998), .S1(n1002), .Y(
        n957) );
  MXI4X1 U1868 ( .A(\blocktag[0][7] ), .B(\blocktag[1][7] ), .C(
        \blocktag[2][7] ), .D(\blocktag[3][7] ), .S0(n998), .S1(n1030), .Y(
        n954) );
  MXI4X1 U1869 ( .A(\blocktag[4][7] ), .B(\blocktag[5][7] ), .C(
        \blocktag[6][7] ), .D(\blocktag[7][7] ), .S0(n998), .S1(n1002), .Y(
        n955) );
  MXI4X1 U1870 ( .A(\blocktag[0][12] ), .B(\blocktag[1][12] ), .C(
        \blocktag[2][12] ), .D(\blocktag[3][12] ), .S0(n998), .S1(n1002), .Y(
        n944) );
  MXI4X1 U1871 ( .A(\blocktag[4][12] ), .B(\blocktag[5][12] ), .C(
        \blocktag[6][12] ), .D(\blocktag[7][12] ), .S0(n998), .S1(n1030), .Y(
        n945) );
  MXI4X1 U1872 ( .A(\blocktag[0][16] ), .B(\blocktag[1][16] ), .C(
        \blocktag[2][16] ), .D(\blocktag[3][16] ), .S0(n997), .S1(n1031), .Y(
        n936) );
  MXI4X1 U1873 ( .A(\blocktag[4][16] ), .B(\blocktag[5][16] ), .C(
        \blocktag[6][16] ), .D(\blocktag[7][16] ), .S0(n997), .S1(n1002), .Y(
        n937) );
  MXI4X1 U1874 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n997), .S1(n1031), .Y(
        n934) );
  MXI4X1 U1875 ( .A(\blocktag[4][17] ), .B(\blocktag[5][17] ), .C(
        \blocktag[6][17] ), .D(\blocktag[7][17] ), .S0(n997), .S1(n1031), .Y(
        n935) );
  MXI4X1 U1876 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n997), .S1(n1002), .Y(
        n932) );
  MXI4X1 U1877 ( .A(\blocktag[4][18] ), .B(\blocktag[5][18] ), .C(
        \blocktag[6][18] ), .D(\blocktag[7][18] ), .S0(n997), .S1(n1031), .Y(
        n933) );
  MXI4X1 U1878 ( .A(\blocktag[0][19] ), .B(\blocktag[1][19] ), .C(
        \blocktag[2][19] ), .D(\blocktag[3][19] ), .S0(n997), .S1(n1030), .Y(
        n930) );
  MXI4X1 U1879 ( .A(\blocktag[4][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[7][22] ), .S0(n996), .S1(n1030), .Y(
        n925) );
  MXI4X1 U1880 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n996), .S1(n1027), .Y(
        n921) );
  NAND4X1 U1881 ( .A(n442), .B(n443), .C(n444), .D(n445), .Y(n438) );
  XNOR2X1 U1882 ( .A(proc_addr[25]), .B(tag[20]), .Y(n442) );
  XNOR2X1 U1883 ( .A(proc_addr[8]), .B(tag[3]), .Y(n443) );
  XNOR2X1 U1884 ( .A(proc_addr[6]), .B(tag[1]), .Y(n444) );
  NOR2BX2 U1885 ( .AN(n163), .B(n164), .Y(n147) );
  MXI2X1 U1886 ( .A(n918), .B(n919), .S0(n1042), .Y(dirty) );
  OAI21XL U1887 ( .A0(n256), .A1(dirty), .B0(valid), .Y(n433) );
  OAI22XL U1888 ( .A0(n471), .A1(n1255), .B0(n147), .B1(n148), .Y(n487) );
  OAI22XL U1889 ( .A0(n472), .A1(n1256), .B0(n147), .B1(n150), .Y(n488) );
  OAI22XL U1890 ( .A0(n473), .A1(n1253), .B0(n147), .B1(n152), .Y(n489) );
  OAI22XL U1891 ( .A0(n474), .A1(n1254), .B0(n147), .B1(n154), .Y(n490) );
  OAI22XL U1892 ( .A0(n475), .A1(n1251), .B0(n147), .B1(n156), .Y(n491) );
  OAI22XL U1893 ( .A0(n476), .A1(n1252), .B0(n147), .B1(n158), .Y(n492) );
  OAI22XL U1894 ( .A0(n477), .A1(n1249), .B0(n147), .B1(n160), .Y(n493) );
  OAI22XL U1895 ( .A0(n478), .A1(n1250), .B0(n147), .B1(n162), .Y(n494) );
  AND2X2 U1896 ( .A(n255), .B(n613), .Y(n261) );
  AOI21X2 U1897 ( .A0(n1175), .A1(n613), .B0(valid), .Y(n166) );
  MXI2X1 U1898 ( .A(n742), .B(n743), .S0(n1037), .Y(blockdata[96]) );
  MXI4X1 U1899 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n982), .S1(n1011), .Y(n742) );
  MXI4X1 U1900 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n981), .S1(n1011), .Y(n743) );
  MXI2X1 U1901 ( .A(n740), .B(n741), .S0(n1037), .Y(blockdata[97]) );
  MXI4X1 U1902 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n981), .S1(n1011), .Y(n740) );
  MXI4X1 U1903 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n981), .S1(n1011), .Y(n741) );
  MXI2X1 U1904 ( .A(n738), .B(n739), .S0(n1037), .Y(blockdata[98]) );
  MXI4X1 U1905 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n981), .S1(n1011), .Y(n738) );
  MXI4X1 U1906 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n981), .S1(n1011), .Y(n739) );
  MXI2X1 U1907 ( .A(n736), .B(n737), .S0(n1037), .Y(blockdata[99]) );
  MXI4X1 U1908 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n981), .S1(n1010), .Y(n736) );
  MXI4X1 U1909 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n981), .S1(n1010), .Y(n737) );
  MXI2X1 U1910 ( .A(n734), .B(n735), .S0(n1037), .Y(blockdata[100]) );
  MXI4X1 U1911 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n981), .S1(n1010), .Y(n734) );
  MXI4X1 U1912 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n981), .S1(n1010), .Y(n735) );
  MXI2X1 U1913 ( .A(n732), .B(n733), .S0(n1037), .Y(blockdata[101]) );
  MXI4X1 U1914 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n981), .S1(n1010), .Y(n732) );
  MXI4X1 U1915 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n981), .S1(n1010), .Y(n733) );
  MXI2X1 U1916 ( .A(n730), .B(n731), .S0(n1037), .Y(blockdata[102]) );
  MXI4X1 U1917 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n981), .S1(n1010), .Y(n730) );
  MXI4X1 U1918 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n981), .S1(n1010), .Y(n731) );
  MXI2X1 U1919 ( .A(n728), .B(n729), .S0(n1037), .Y(blockdata[103]) );
  MXI4X1 U1920 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n980), .S1(n1010), .Y(n728) );
  MXI4X1 U1921 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n980), .S1(n1010), .Y(n729) );
  MXI2X1 U1922 ( .A(n726), .B(n727), .S0(n1037), .Y(blockdata[104]) );
  MXI4X1 U1923 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n980), .S1(n1010), .Y(n726) );
  MXI4X1 U1924 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n980), .S1(n1010), .Y(n727) );
  MXI2X1 U1925 ( .A(n724), .B(n725), .S0(n1036), .Y(blockdata[105]) );
  MXI4X1 U1926 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n980), .S1(n1009), .Y(n724) );
  MXI4X1 U1927 ( .A(\block[4][105] ), .B(\block[5][105] ), .C(\block[6][105] ), 
        .D(\block[7][105] ), .S0(n980), .S1(n1009), .Y(n725) );
  MXI2X1 U1928 ( .A(n722), .B(n723), .S0(n1036), .Y(blockdata[106]) );
  MXI4X1 U1929 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n980), .S1(n1009), .Y(n722) );
  MXI4X1 U1930 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n980), .S1(n1009), .Y(n723) );
  MXI2X1 U1931 ( .A(n720), .B(n721), .S0(n1036), .Y(blockdata[107]) );
  MXI4X1 U1932 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n980), .S1(n1009), .Y(n720) );
  MXI4X1 U1933 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n980), .S1(n1009), .Y(n721) );
  MXI2X1 U1934 ( .A(n718), .B(n719), .S0(n1036), .Y(blockdata[108]) );
  MXI4X1 U1935 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n980), .S1(n1009), .Y(n718) );
  MXI4X1 U1936 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n980), .S1(n1009), .Y(n719) );
  MXI2X1 U1937 ( .A(n716), .B(n717), .S0(n1036), .Y(blockdata[109]) );
  MXI4X1 U1938 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n980), .S1(n1009), .Y(n716) );
  MXI4X1 U1939 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n979), .S1(n1009), .Y(n717) );
  MXI2X1 U1940 ( .A(n714), .B(n715), .S0(n1036), .Y(blockdata[110]) );
  MXI4X1 U1941 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n979), .S1(n1009), .Y(n714) );
  MXI4X1 U1942 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n979), .S1(n1009), .Y(n715) );
  MXI2X1 U1943 ( .A(n712), .B(n713), .S0(n1036), .Y(blockdata[111]) );
  MXI4X1 U1944 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n979), .S1(n1008), .Y(n712) );
  MXI4X1 U1945 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n979), .S1(n1008), .Y(n713) );
  MXI2X1 U1946 ( .A(n710), .B(n711), .S0(n1036), .Y(blockdata[112]) );
  MXI4X1 U1947 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n979), .S1(n1008), .Y(n710) );
  MXI4X1 U1948 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n979), .S1(n1008), .Y(n711) );
  MXI2X1 U1949 ( .A(n708), .B(n709), .S0(n1036), .Y(blockdata[113]) );
  MXI4X1 U1950 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n979), .S1(n1008), .Y(n708) );
  MXI4X1 U1951 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n979), .S1(n1008), .Y(n709) );
  MXI2X1 U1952 ( .A(n706), .B(n707), .S0(n1036), .Y(blockdata[114]) );
  MXI4X1 U1953 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n979), .S1(n1008), .Y(n706) );
  MXI4X1 U1954 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n979), .S1(n1008), .Y(n707) );
  MXI2X1 U1955 ( .A(n704), .B(n705), .S0(n1036), .Y(blockdata[115]) );
  MXI4X1 U1956 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n979), .S1(n1008), .Y(n704) );
  MXI4X1 U1957 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n979), .S1(n1008), .Y(n705) );
  MXI2X1 U1958 ( .A(n702), .B(n703), .S0(n1036), .Y(blockdata[116]) );
  MXI4X1 U1959 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n978), .S1(n1008), .Y(n702) );
  MXI4X1 U1960 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n978), .S1(n1008), .Y(n703) );
  MXI2X1 U1961 ( .A(n700), .B(n701), .S0(n1035), .Y(blockdata[117]) );
  MXI4X1 U1962 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n978), .S1(n1007), .Y(n700) );
  MXI4X1 U1963 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n978), .S1(n1007), .Y(n701) );
  MXI2X1 U1964 ( .A(n698), .B(n699), .S0(n1035), .Y(blockdata[118]) );
  MXI4X1 U1965 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n978), .S1(n1007), .Y(n698) );
  MXI4X1 U1966 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n978), .S1(n1007), .Y(n699) );
  MXI2X1 U1967 ( .A(n696), .B(n697), .S0(n1035), .Y(blockdata[119]) );
  MXI4X1 U1968 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n978), .S1(n1007), .Y(n696) );
  MXI4X1 U1969 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n978), .S1(n1007), .Y(n697) );
  MXI2X1 U1970 ( .A(n694), .B(n695), .S0(n1035), .Y(blockdata[120]) );
  MXI4X1 U1971 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n978), .S1(n1007), .Y(n694) );
  MXI4X1 U1972 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n978), .S1(n1007), .Y(n695) );
  MXI2X1 U1973 ( .A(n692), .B(n693), .S0(n1035), .Y(blockdata[121]) );
  MXI4X1 U1974 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n978), .S1(n1007), .Y(n692) );
  MXI4X1 U1975 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n978), .S1(n1007), .Y(n693) );
  MXI2X1 U1976 ( .A(n690), .B(n691), .S0(n1035), .Y(blockdata[122]) );
  MXI4X1 U1977 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n994), .S1(n1007), .Y(n691) );
  MXI4X1 U1978 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n978), .S1(n1007), .Y(n690) );
  MXI2X1 U1979 ( .A(n688), .B(n689), .S0(n1035), .Y(blockdata[123]) );
  MXI4X1 U1980 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n985), .S1(n1015), .Y(n688) );
  MXI4X1 U1981 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n991), .S1(n1022), .Y(n689) );
  MXI2X1 U1982 ( .A(n686), .B(n687), .S0(n1035), .Y(blockdata[124]) );
  MXI4X1 U1983 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n989), .S1(n1014), .Y(n686) );
  MXI4X1 U1984 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n990), .S1(n1021), .Y(n687) );
  MXI2X1 U1985 ( .A(n684), .B(n685), .S0(n1035), .Y(blockdata[125]) );
  MXI4X1 U1986 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n988), .S1(n1013), .Y(n684) );
  MXI4X1 U1987 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n992), .S1(n1020), .Y(n685) );
  MXI2X1 U1988 ( .A(n682), .B(n683), .S0(n1035), .Y(blockdata[126]) );
  MXI4X1 U1989 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n985), .S1(n1012), .Y(n682) );
  MXI4X1 U1990 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n993), .S1(n1017), .Y(n683) );
  MXI2X1 U1991 ( .A(n680), .B(n681), .S0(n1035), .Y(blockdata[127]) );
  MXI4X1 U1992 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n989), .S1(n1016), .Y(n680) );
  MXI4X1 U1993 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n986), .S1(n1019), .Y(n681) );
  NOR2X1 U1994 ( .A(n615), .B(n150), .Y(N1769) );
  NOR2X1 U1995 ( .A(n615), .B(n148), .Y(N1768) );
  NOR2X1 U1996 ( .A(n615), .B(n152), .Y(N1771) );
  NOR2X1 U1997 ( .A(n615), .B(n154), .Y(N1772) );
  NOR2X1 U1998 ( .A(n615), .B(n156), .Y(N1773) );
  NOR2X1 U1999 ( .A(n615), .B(n158), .Y(N1774) );
  NOR2X1 U2000 ( .A(n615), .B(n160), .Y(N1776) );
  NOR2X1 U2001 ( .A(n615), .B(n162), .Y(N1777) );
  OAI22XL U2002 ( .A0(n479), .A1(n1255), .B0(n166), .B1(n148), .Y(n495) );
  OAI22XL U2003 ( .A0(n480), .A1(n1256), .B0(n166), .B1(n150), .Y(n496) );
  OAI22XL U2004 ( .A0(n481), .A1(n1253), .B0(n166), .B1(n152), .Y(n497) );
  OAI22XL U2005 ( .A0(n482), .A1(n1254), .B0(n166), .B1(n154), .Y(n498) );
  OAI22XL U2006 ( .A0(n483), .A1(n1251), .B0(n166), .B1(n156), .Y(n499) );
  OAI22XL U2007 ( .A0(n484), .A1(n1252), .B0(n166), .B1(n158), .Y(n500) );
  OAI22XL U2008 ( .A0(n485), .A1(n1249), .B0(n166), .B1(n160), .Y(n501) );
  OAI22XL U2009 ( .A0(n486), .A1(n1250), .B0(n166), .B1(n162), .Y(n503) );
  CLKINVX1 U2010 ( .A(proc_wdata[4]), .Y(n1286) );
  CLKINVX1 U2011 ( .A(proc_wdata[5]), .Y(n1285) );
  CLKINVX1 U2012 ( .A(proc_wdata[6]), .Y(n1284) );
  CLKINVX1 U2013 ( .A(proc_wdata[7]), .Y(n1283) );
  CLKINVX1 U2014 ( .A(proc_wdata[8]), .Y(n1282) );
  CLKINVX1 U2015 ( .A(proc_wdata[10]), .Y(n1280) );
  CLKINVX1 U2016 ( .A(proc_wdata[11]), .Y(n1279) );
  CLKINVX1 U2017 ( .A(proc_wdata[12]), .Y(n1278) );
  CLKINVX1 U2018 ( .A(proc_wdata[13]), .Y(n1277) );
  CLKINVX1 U2019 ( .A(proc_wdata[14]), .Y(n1276) );
  CLKINVX1 U2020 ( .A(proc_wdata[15]), .Y(n1275) );
  CLKINVX1 U2021 ( .A(proc_wdata[16]), .Y(n1274) );
  CLKINVX1 U2022 ( .A(proc_wdata[17]), .Y(n1273) );
  CLKINVX1 U2023 ( .A(proc_wdata[18]), .Y(n1272) );
  CLKINVX1 U2024 ( .A(proc_wdata[19]), .Y(n1271) );
  CLKINVX1 U2025 ( .A(proc_wdata[20]), .Y(n1270) );
  CLKINVX1 U2026 ( .A(proc_wdata[21]), .Y(n1269) );
  CLKINVX1 U2027 ( .A(proc_wdata[22]), .Y(n1268) );
  CLKINVX1 U2028 ( .A(proc_wdata[23]), .Y(n1267) );
  CLKINVX1 U2029 ( .A(proc_wdata[24]), .Y(n1266) );
  CLKINVX1 U2030 ( .A(proc_wdata[25]), .Y(n1265) );
  CLKINVX1 U2031 ( .A(proc_wdata[26]), .Y(n1264) );
  CLKINVX1 U2032 ( .A(proc_wdata[27]), .Y(n1263) );
  CLKINVX1 U2033 ( .A(proc_wdata[28]), .Y(n1262) );
  CLKINVX1 U2034 ( .A(proc_wdata[29]), .Y(n1261) );
  CLKINVX1 U2035 ( .A(proc_wdata[30]), .Y(n1260) );
  CLKINVX1 U2036 ( .A(proc_wdata[31]), .Y(n1259) );
  CLKINVX1 U2037 ( .A(proc_wdata[0]), .Y(n1290) );
  CLKINVX1 U2038 ( .A(proc_wdata[1]), .Y(n1289) );
  CLKINVX1 U2039 ( .A(proc_wdata[2]), .Y(n1288) );
  CLKINVX1 U2040 ( .A(proc_wdata[3]), .Y(n1287) );
  CLKINVX1 U2041 ( .A(proc_wdata[9]), .Y(n1281) );
  MXI4X1 U2042 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n986), .S1(n1016), .Y(n806) );
  MXI4X1 U2043 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n986), .S1(n1016), .Y(n807) );
  MXI4X1 U2044 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n986), .S1(n1016), .Y(n804) );
  MXI4X1 U2045 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n986), .S1(n1016), .Y(n805) );
  MXI4X1 U2046 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n986), .S1(n1016), .Y(n802) );
  MXI4X1 U2047 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n986), .S1(n1016), .Y(n803) );
  MXI4X1 U2048 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n986), .S1(n1016), .Y(n800) );
  MXI4X1 U2049 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n986), .S1(n1016), .Y(n801) );
  MXI4X1 U2050 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n986), .S1(n1016), .Y(n798) );
  MXI4X1 U2051 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n986), .S1(n1016), .Y(n799) );
  MXI4X1 U2052 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n986), .S1(n1015), .Y(n796) );
  MXI4X1 U2053 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n986), .S1(n1015), .Y(n797) );
  MXI4X1 U2054 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n986), .S1(n1015), .Y(n794) );
  MXI4X1 U2055 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n985), .S1(n1015), .Y(n795) );
  MXI4X1 U2056 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n985), .S1(n1015), .Y(n792) );
  MXI4X1 U2057 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n985), .S1(n1015), .Y(n793) );
  MXI4X1 U2058 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n985), .S1(n1015), .Y(n790) );
  MXI4X1 U2059 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n985), .S1(n1015), .Y(n791) );
  MXI4X1 U2060 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n985), .S1(n1015), .Y(n788) );
  MXI4X1 U2061 ( .A(\block[4][73] ), .B(\block[5][73] ), .C(\block[6][73] ), 
        .D(\block[7][73] ), .S0(n985), .S1(n1015), .Y(n789) );
  MXI4X1 U2062 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n985), .S1(n1015), .Y(n786) );
  MXI4X1 U2063 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n985), .S1(n1015), .Y(n787) );
  MXI4X1 U2064 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n985), .S1(n1014), .Y(n784) );
  MXI4X1 U2065 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n985), .S1(n1014), .Y(n785) );
  MXI4X1 U2066 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n985), .S1(n1014), .Y(n782) );
  MXI4X1 U2067 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n985), .S1(n1014), .Y(n783) );
  MXI4X1 U2068 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n984), .S1(n1014), .Y(n780) );
  MXI4X1 U2069 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n984), .S1(n1014), .Y(n781) );
  MXI4X1 U2070 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n984), .S1(n1014), .Y(n778) );
  MXI4X1 U2071 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n984), .S1(n1014), .Y(n779) );
  MXI4X1 U2072 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n984), .S1(n1014), .Y(n776) );
  MXI4X1 U2073 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n984), .S1(n1014), .Y(n777) );
  MXI4X1 U2074 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n984), .S1(n1014), .Y(n774) );
  MXI4X1 U2075 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n984), .S1(n1014), .Y(n775) );
  MXI4X1 U2076 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n984), .S1(n1013), .Y(n772) );
  MXI4X1 U2077 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n984), .S1(n1013), .Y(n773) );
  MXI4X1 U2078 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n984), .S1(n1013), .Y(n770) );
  MXI4X1 U2079 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n984), .S1(n1013), .Y(n771) );
  MXI4X1 U2080 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n984), .S1(n1013), .Y(n768) );
  MXI4X1 U2081 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n983), .S1(n1013), .Y(n769) );
  MXI4X1 U2082 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n983), .S1(n1013), .Y(n766) );
  MXI4X1 U2083 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n983), .S1(n1013), .Y(n767) );
  MXI4X1 U2084 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n983), .S1(n1013), .Y(n764) );
  MXI4X1 U2085 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n983), .S1(n1013), .Y(n765) );
  MXI4X1 U2086 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n983), .S1(n1013), .Y(n762) );
  MXI4X1 U2087 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n983), .S1(n1013), .Y(n763) );
  MXI4X1 U2088 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n983), .S1(n1012), .Y(n760) );
  MXI4X1 U2089 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n983), .S1(n1012), .Y(n761) );
  MXI4X1 U2090 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n983), .S1(n1012), .Y(n758) );
  MXI4X1 U2091 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n983), .S1(n1012), .Y(n759) );
  MXI4X1 U2092 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n983), .S1(n1012), .Y(n756) );
  MXI4X1 U2093 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n983), .S1(n1012), .Y(n757) );
  MXI4X1 U2094 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n982), .S1(n1012), .Y(n754) );
  MXI4X1 U2095 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n982), .S1(n1012), .Y(n755) );
  MXI4X1 U2096 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n982), .S1(n1012), .Y(n752) );
  MXI4X1 U2097 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n982), .S1(n1012), .Y(n753) );
  MXI4X1 U2098 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n982), .S1(n1012), .Y(n750) );
  MXI4X1 U2099 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n982), .S1(n1012), .Y(n751) );
  MXI4X1 U2100 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n982), .S1(n1011), .Y(n748) );
  MXI4X1 U2101 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n982), .S1(n1011), .Y(n749) );
  MXI4X1 U2102 ( .A(\block[0][94] ), .B(\block[1][94] ), .C(\block[2][94] ), 
        .D(\block[3][94] ), .S0(n982), .S1(n1011), .Y(n746) );
  MXI4X1 U2103 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), 
        .D(\block[7][94] ), .S0(n982), .S1(n1011), .Y(n747) );
  MXI4X1 U2104 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n982), .S1(n1011), .Y(n744) );
  MXI4X1 U2105 ( .A(\block[4][95] ), .B(\block[5][95] ), .C(\block[6][95] ), 
        .D(\block[7][95] ), .S0(n982), .S1(n1011), .Y(n745) );
  MXI4X1 U2106 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n990), .S1(n1022), .Y(n870) );
  MXI4X1 U2107 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n990), .S1(n1022), .Y(n871) );
  MXI4X1 U2108 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n990), .S1(n1021), .Y(n868) );
  MXI4X1 U2109 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n990), .S1(n1021), .Y(n869) );
  MXI4X1 U2110 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n990), .S1(n1021), .Y(n866) );
  MXI4X1 U2111 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n990), .S1(n1021), .Y(n867) );
  MXI4X1 U2112 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n990), .S1(n1021), .Y(n864) );
  MXI4X1 U2113 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n990), .S1(n1021), .Y(n865) );
  MXI4X1 U2114 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n990), .S1(n1021), .Y(n862) );
  MXI4X1 U2115 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n990), .S1(n1021), .Y(n863) );
  MXI4X1 U2116 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n990), .S1(n1021), .Y(n860) );
  MXI4X1 U2117 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n990), .S1(n1021), .Y(n861) );
  MXI4X1 U2118 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n989), .S1(n1021), .Y(n858) );
  MXI4X1 U2119 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n989), .S1(n1021), .Y(n859) );
  MXI4X1 U2120 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n989), .S1(n1020), .Y(n856) );
  MXI4X1 U2121 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n989), .S1(n1020), .Y(n857) );
  MXI4X1 U2122 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n989), .S1(n1020), .Y(n854) );
  MXI4X1 U2123 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n989), .S1(n1020), .Y(n855) );
  MXI4X1 U2124 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n989), .S1(n1020), .Y(n852) );
  MXI4X1 U2125 ( .A(\block[4][41] ), .B(\block[5][41] ), .C(\block[6][41] ), 
        .D(\block[7][41] ), .S0(n989), .S1(n1020), .Y(n853) );
  MXI4X1 U2126 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n989), .S1(n1020), .Y(n850) );
  MXI4X1 U2127 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n989), .S1(n1020), .Y(n851) );
  MXI4X1 U2128 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n989), .S1(n1020), .Y(n848) );
  MXI4X1 U2129 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n989), .S1(n1020), .Y(n849) );
  MXI4X1 U2130 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n989), .S1(n1020), .Y(n846) );
  MXI4X1 U2131 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n988), .S1(n1020), .Y(n847) );
  MXI4X1 U2132 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n988), .S1(n1019), .Y(n844) );
  MXI4X1 U2133 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n988), .S1(n1019), .Y(n845) );
  MXI4X1 U2134 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n988), .S1(n1019), .Y(n842) );
  MXI4X1 U2135 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n988), .S1(n1019), .Y(n843) );
  MXI4X1 U2136 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n988), .S1(n1019), .Y(n840) );
  MXI4X1 U2137 ( .A(\block[4][47] ), .B(\block[5][47] ), .C(\block[6][47] ), 
        .D(\block[7][47] ), .S0(n988), .S1(n1019), .Y(n841) );
  MXI4X1 U2138 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n988), .S1(n1019), .Y(n838) );
  MXI4X1 U2139 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n988), .S1(n1019), .Y(n839) );
  MXI4X1 U2140 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n988), .S1(n1019), .Y(n836) );
  MXI4X1 U2141 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n988), .S1(n1019), .Y(n837) );
  MXI4X1 U2142 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n988), .S1(n1019), .Y(n834) );
  MXI4X1 U2143 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n988), .S1(n1019), .Y(n835) );
  MXI4X1 U2144 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n987), .S1(n1018), .Y(n832) );
  MXI4X1 U2145 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n987), .S1(n1018), .Y(n833) );
  MXI4X1 U2146 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n987), .S1(n1018), .Y(n830) );
  MXI4X1 U2147 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n987), .S1(n1018), .Y(n831) );
  MXI4X1 U2148 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n987), .S1(n1018), .Y(n828) );
  MXI4X1 U2149 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n987), .S1(n1018), .Y(n829) );
  MXI4X1 U2150 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n987), .S1(n1018), .Y(n826) );
  MXI4X1 U2151 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n987), .S1(n1018), .Y(n827) );
  MXI4X1 U2152 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n987), .S1(n1018), .Y(n824) );
  MXI4X1 U2153 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n987), .S1(n1018), .Y(n825) );
  MXI4X1 U2154 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n987), .S1(n1018), .Y(n822) );
  MXI4X1 U2155 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n987), .S1(n1018), .Y(n823) );
  MXI4X1 U2156 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n987), .S1(n1017), .Y(n820) );
  MXI4X1 U2157 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n993), .S1(n1017), .Y(n821) );
  MXI4X1 U2158 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n993), .S1(n1017), .Y(n818) );
  MXI4X1 U2159 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n992), .S1(n1017), .Y(n819) );
  MXI4X1 U2160 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n988), .S1(n1017), .Y(n816) );
  MXI4X1 U2161 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n988), .S1(n1017), .Y(n817) );
  MXI4X1 U2162 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n992), .S1(n1017), .Y(n814) );
  MXI4X1 U2163 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n991), .S1(n1017), .Y(n815) );
  MXI4X1 U2164 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n990), .S1(n1017), .Y(n812) );
  MXI4X1 U2165 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n985), .S1(n1017), .Y(n813) );
  MXI4X1 U2166 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n986), .S1(n1017), .Y(n810) );
  MXI4X1 U2167 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n986), .S1(n1017), .Y(n811) );
  MXI4X1 U2168 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n991), .S1(n1016), .Y(n808) );
  MXI4X1 U2169 ( .A(\block[4][63] ), .B(\block[5][63] ), .C(\block[6][63] ), 
        .D(\block[7][63] ), .S0(n990), .S1(n1016), .Y(n809) );
  MXI4X1 U2170 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n994), .S1(n1025), .Y(n916) );
  MXI4X1 U2171 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n994), .S1(n1025), .Y(n917) );
  MXI4X1 U2172 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n994), .S1(n1025), .Y(n914) );
  MXI4X1 U2173 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n994), .S1(n1025), .Y(n915) );
  MXI4X1 U2174 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n994), .S1(n1025), .Y(n912) );
  MXI4X1 U2175 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n994), .S1(n1025), .Y(n913) );
  MXI4X1 U2176 ( .A(\block[0][12] ), .B(\block[1][12] ), .C(\block[2][12] ), 
        .D(\block[3][12] ), .S0(n993), .S1(n1025), .Y(n910) );
  MXI4X1 U2177 ( .A(\block[4][12] ), .B(\block[5][12] ), .C(\block[6][12] ), 
        .D(\block[7][12] ), .S0(n993), .S1(n1025), .Y(n911) );
  MXI4X1 U2178 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n993), .S1(n1025), .Y(n908) );
  MXI4X1 U2179 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n993), .S1(n1025), .Y(n909) );
  MXI4X1 U2180 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n993), .S1(n1025), .Y(n906) );
  MXI4X1 U2181 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n993), .S1(n1025), .Y(n907) );
  MXI4X1 U2182 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n993), .S1(n1024), .Y(n904) );
  MXI4X1 U2183 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n993), .S1(n1024), .Y(n905) );
  MXI4X1 U2184 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n993), .S1(n1024), .Y(n902) );
  MXI4X1 U2185 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n993), .S1(n1024), .Y(n903) );
  MXI4X1 U2186 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n993), .S1(n1024), .Y(n900) );
  MXI4X1 U2187 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n993), .S1(n1024), .Y(n901) );
  MXI4X1 U2188 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n993), .S1(n1024), .Y(n898) );
  MXI4X1 U2189 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n992), .S1(n1024), .Y(n899) );
  MXI4X1 U2190 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n992), .S1(n1024), .Y(n896) );
  MXI4X1 U2191 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n992), .S1(n1024), .Y(n897) );
  MXI4X1 U2192 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n992), .S1(n1024), .Y(n894) );
  MXI4X1 U2193 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n992), .S1(n1024), .Y(n895) );
  MXI4X1 U2194 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n992), .S1(n1023), .Y(n892) );
  MXI4X1 U2195 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n992), .S1(n1023), .Y(n893) );
  MXI4X1 U2196 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n992), .S1(n1023), .Y(n890) );
  MXI4X1 U2197 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n992), .S1(n1023), .Y(n891) );
  MXI4X1 U2198 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n992), .S1(n1023), .Y(n888) );
  MXI4X1 U2199 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n992), .S1(n1023), .Y(n889) );
  MXI4X1 U2200 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n992), .S1(n1023), .Y(n886) );
  MXI4X1 U2201 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n992), .S1(n1023), .Y(n887) );
  MXI4X1 U2202 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n991), .S1(n1023), .Y(n884) );
  MXI4X1 U2203 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n991), .S1(n1023), .Y(n885) );
  MXI4X1 U2204 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n991), .S1(n1023), .Y(n882) );
  MXI4X1 U2205 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n991), .S1(n1023), .Y(n883) );
  MXI4X1 U2206 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n991), .S1(n1022), .Y(n880) );
  MXI4X1 U2207 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n991), .S1(n1022), .Y(n881) );
  MXI4X1 U2208 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n991), .S1(n1022), .Y(n878) );
  MXI4X1 U2209 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n991), .S1(n1022), .Y(n879) );
  MXI4X1 U2210 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n991), .S1(n1022), .Y(n876) );
  MXI4X1 U2211 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n991), .S1(n1022), .Y(n877) );
  MXI4X1 U2212 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n991), .S1(n1022), .Y(n874) );
  MXI4X1 U2213 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n991), .S1(n1022), .Y(n875) );
  MXI4X1 U2214 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n991), .S1(n1022), .Y(n872) );
  MXI4X1 U2215 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n990), .S1(n1022), .Y(n873) );
  CLKINVX1 U2216 ( .A(proc_read), .Y(n1174) );
  CLKINVX1 U2217 ( .A(proc_addr[5]), .Y(n1203) );
  CLKINVX1 U2218 ( .A(proc_addr[6]), .Y(n1202) );
  CLKINVX1 U2219 ( .A(proc_addr[7]), .Y(n1201) );
  CLKINVX1 U2220 ( .A(proc_addr[8]), .Y(n1200) );
  CLKINVX1 U2221 ( .A(proc_addr[9]), .Y(n1199) );
  CLKINVX1 U2222 ( .A(proc_addr[10]), .Y(n1198) );
  CLKINVX1 U2223 ( .A(proc_addr[11]), .Y(n1197) );
  CLKINVX1 U2224 ( .A(proc_addr[12]), .Y(n1196) );
  CLKINVX1 U2225 ( .A(proc_addr[13]), .Y(n1195) );
  CLKINVX1 U2226 ( .A(proc_addr[14]), .Y(n1194) );
  CLKINVX1 U2227 ( .A(proc_addr[15]), .Y(n1193) );
  CLKINVX1 U2228 ( .A(proc_addr[16]), .Y(n1192) );
  CLKINVX1 U2229 ( .A(proc_addr[17]), .Y(n1191) );
  CLKINVX1 U2230 ( .A(proc_addr[18]), .Y(n1190) );
  CLKINVX1 U2231 ( .A(proc_addr[19]), .Y(n1189) );
  CLKINVX1 U2232 ( .A(proc_addr[20]), .Y(n1188) );
  CLKINVX1 U2233 ( .A(proc_addr[21]), .Y(n1187) );
  CLKINVX1 U2234 ( .A(proc_addr[22]), .Y(n1186) );
  CLKINVX1 U2235 ( .A(proc_addr[23]), .Y(n1185) );
  CLKINVX1 U2236 ( .A(proc_addr[24]), .Y(n1184) );
  CLKINVX1 U2237 ( .A(proc_addr[25]), .Y(n1183) );
  CLKINVX1 U2238 ( .A(proc_addr[26]), .Y(n1182) );
  CLKINVX1 U2239 ( .A(proc_addr[27]), .Y(n1181) );
  CLKINVX1 U2240 ( .A(proc_addr[28]), .Y(n1180) );
  CLKINVX1 U2241 ( .A(proc_addr[29]), .Y(n1178) );
  INVX3 U2242 ( .A(n615), .Y(n1173) );
endmodule

