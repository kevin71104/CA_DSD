
module IF_DEC_regFile ( clk, rst_n, flush, stallcache, stall_lw_use, 
        instruction_next, PCplus4, branchOffset, opcode, Rs, Rt, Rd, shamt, 
        funct, immediate, instruction_regI, PCplus4_regI );
  input [31:0] instruction_next;
  input [31:0] PCplus4;
  output [15:0] branchOffset;
  output [5:0] opcode;
  output [4:0] Rs;
  output [4:0] Rt;
  output [4:0] Rd;
  output [4:0] shamt;
  output [5:0] funct;
  output [15:0] immediate;
  output [31:0] instruction_regI;
  output [31:0] PCplus4_regI;
  input clk, rst_n, flush, stallcache, stall_lw_use;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n1, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145;

  DFFRX4 \instruction_regI_reg[29]  ( .D(n32), .CK(clk), .RN(n137), .Q(
        opcode[3]) );
  DFFRX4 \instruction_regI_reg[28]  ( .D(n31), .CK(clk), .RN(n137), .Q(
        opcode[2]) );
  DFFRX4 \instruction_regI_reg[27]  ( .D(n30), .CK(clk), .RN(n137), .Q(
        opcode[1]) );
  DFFRX4 \instruction_regI_reg[25]  ( .D(n28), .CK(clk), .RN(n137), .Q(Rs[4])
         );
  DFFRX4 \instruction_regI_reg[22]  ( .D(n25), .CK(clk), .RN(n136), .Q(Rs[1])
         );
  DFFRX1 \PCplus4_regI_reg[31]  ( .D(n66), .CK(clk), .RN(n140), .Q(
        PCplus4_regI[31]) );
  DFFRX1 \PCplus4_regI_reg[30]  ( .D(n65), .CK(clk), .RN(n140), .Q(
        PCplus4_regI[30]) );
  DFFRX1 \PCplus4_regI_reg[29]  ( .D(n64), .CK(clk), .RN(n140), .Q(
        PCplus4_regI[29]) );
  DFFRX1 \PCplus4_regI_reg[28]  ( .D(n63), .CK(clk), .RN(n140), .Q(
        PCplus4_regI[28]) );
  DFFRX1 \PCplus4_regI_reg[27]  ( .D(n62), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[27]) );
  DFFRX1 \PCplus4_regI_reg[26]  ( .D(n61), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[26]) );
  DFFRX1 \PCplus4_regI_reg[25]  ( .D(n60), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[25]) );
  DFFRX1 \PCplus4_regI_reg[24]  ( .D(n59), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[24]) );
  DFFRX1 \PCplus4_regI_reg[23]  ( .D(n58), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[23]) );
  DFFRX1 \PCplus4_regI_reg[22]  ( .D(n57), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[22]) );
  DFFRX1 \PCplus4_regI_reg[21]  ( .D(n56), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[21]) );
  DFFRX1 \PCplus4_regI_reg[20]  ( .D(n55), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[20]) );
  DFFRX1 \PCplus4_regI_reg[19]  ( .D(n54), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[19]) );
  DFFRX1 \PCplus4_regI_reg[18]  ( .D(n53), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[18]) );
  DFFRX1 \PCplus4_regI_reg[17]  ( .D(n52), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[17]) );
  DFFRX1 \PCplus4_regI_reg[16]  ( .D(n51), .CK(clk), .RN(n139), .Q(
        PCplus4_regI[16]) );
  DFFRX1 \PCplus4_regI_reg[15]  ( .D(n50), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[15]) );
  DFFRX1 \PCplus4_regI_reg[14]  ( .D(n49), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[14]) );
  DFFRX1 \PCplus4_regI_reg[13]  ( .D(n48), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[13]) );
  DFFRX1 \PCplus4_regI_reg[12]  ( .D(n47), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[12]) );
  DFFRX1 \PCplus4_regI_reg[11]  ( .D(n46), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[11]) );
  DFFRX1 \PCplus4_regI_reg[10]  ( .D(n45), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[10]) );
  DFFRX1 \PCplus4_regI_reg[9]  ( .D(n44), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[9]) );
  DFFRX1 \PCplus4_regI_reg[8]  ( .D(n43), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[8]) );
  DFFRX1 \PCplus4_regI_reg[7]  ( .D(n42), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[7]) );
  DFFRX1 \PCplus4_regI_reg[6]  ( .D(n41), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[6]) );
  DFFRX1 \PCplus4_regI_reg[5]  ( .D(n40), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[5]) );
  DFFRX1 \PCplus4_regI_reg[4]  ( .D(n39), .CK(clk), .RN(n138), .Q(
        PCplus4_regI[4]) );
  DFFRX1 \PCplus4_regI_reg[3]  ( .D(n38), .CK(clk), .RN(n137), .Q(
        PCplus4_regI[3]) );
  DFFRX1 \PCplus4_regI_reg[2]  ( .D(n37), .CK(clk), .RN(n137), .Q(
        PCplus4_regI[2]) );
  DFFRX1 \PCplus4_regI_reg[1]  ( .D(n36), .CK(clk), .RN(n137), .Q(
        PCplus4_regI[1]) );
  DFFRX1 \PCplus4_regI_reg[0]  ( .D(n35), .CK(clk), .RN(n137), .Q(
        PCplus4_regI[0]) );
  DFFRX1 \instruction_regI_reg[30]  ( .D(n33), .CK(clk), .RN(n137), .Q(
        opcode[4]) );
  DFFRX2 \instruction_regI_reg[5]  ( .D(n8), .CK(clk), .RN(n135), .Q(funct[5])
         );
  DFFRX2 \instruction_regI_reg[2]  ( .D(n5), .CK(clk), .RN(n135), .Q(funct[2])
         );
  DFFRX2 \instruction_regI_reg[4]  ( .D(n7), .CK(clk), .RN(n135), .Q(funct[4])
         );
  DFFRX2 \instruction_regI_reg[0]  ( .D(n3), .CK(clk), .RN(n135), .Q(funct[0])
         );
  DFFRX2 \instruction_regI_reg[3]  ( .D(n6), .CK(clk), .RN(n135), .Q(funct[3])
         );
  DFFRX2 \instruction_regI_reg[26]  ( .D(n29), .CK(clk), .RN(n137), .Q(
        opcode[0]) );
  DFFRX2 \instruction_regI_reg[1]  ( .D(n4), .CK(clk), .RN(n135), .Q(funct[1])
         );
  DFFRX1 \instruction_regI_reg[24]  ( .D(n27), .CK(clk), .RN(n137), .Q(Rs[3])
         );
  DFFRX1 \instruction_regI_reg[23]  ( .D(n26), .CK(clk), .RN(n136), .Q(Rs[2])
         );
  DFFRX1 \instruction_regI_reg[19]  ( .D(n22), .CK(clk), .RN(n136), .Q(Rt[3])
         );
  DFFRX1 \instruction_regI_reg[18]  ( .D(n21), .CK(clk), .RN(n136), .Q(Rt[2])
         );
  DFFRX1 \instruction_regI_reg[9]  ( .D(n12), .CK(clk), .RN(n135), .Q(shamt[3]) );
  DFFRX1 \instruction_regI_reg[8]  ( .D(n11), .CK(clk), .RN(n135), .Q(shamt[2]) );
  DFFRX1 \instruction_regI_reg[7]  ( .D(n10), .CK(clk), .RN(n135), .Q(shamt[1]) );
  DFFRX1 \instruction_regI_reg[6]  ( .D(n9), .CK(clk), .RN(n135), .Q(shamt[0])
         );
  DFFRX1 \instruction_regI_reg[14]  ( .D(n17), .CK(clk), .RN(n136), .Q(Rd[3])
         );
  DFFRX1 \instruction_regI_reg[13]  ( .D(n16), .CK(clk), .RN(n136), .Q(Rd[2])
         );
  DFFRX1 \instruction_regI_reg[12]  ( .D(n15), .CK(clk), .RN(n136), .Q(Rd[1])
         );
  DFFRX1 \instruction_regI_reg[11]  ( .D(n14), .CK(clk), .RN(n135), .Q(Rd[0])
         );
  DFFRX1 \instruction_regI_reg[15]  ( .D(n18), .CK(clk), .RN(n136), .Q(Rd[4])
         );
  DFFRX1 \instruction_regI_reg[10]  ( .D(n13), .CK(clk), .RN(n135), .Q(
        shamt[4]) );
  DFFRX2 \instruction_regI_reg[31]  ( .D(n34), .CK(clk), .RN(n137), .Q(
        opcode[5]) );
  DFFRX2 \instruction_regI_reg[20]  ( .D(n23), .CK(clk), .RN(n136), .Q(Rt[4])
         );
  DFFRX2 \instruction_regI_reg[21]  ( .D(n24), .CK(clk), .RN(n136), .Q(Rs[0])
         );
  DFFRX2 \instruction_regI_reg[16]  ( .D(n19), .CK(clk), .RN(n136), .Q(Rt[0])
         );
  DFFRX2 \instruction_regI_reg[17]  ( .D(n20), .CK(clk), .RN(n136), .Q(Rt[1])
         );
  AO22X1 U2 ( .A0(instruction_next[28]), .A1(n131), .B0(opcode[2]), .B1(n144), 
        .Y(n31) );
  CLKINVX8 U3 ( .A(n142), .Y(n145) );
  AO22X2 U4 ( .A0(PCplus4[0]), .A1(n130), .B0(PCplus4_regI[0]), .B1(n144), .Y(
        n35) );
  AO22X2 U5 ( .A0(PCplus4[1]), .A1(n130), .B0(PCplus4_regI[1]), .B1(n144), .Y(
        n36) );
  AO22X2 U6 ( .A0(PCplus4[3]), .A1(n130), .B0(PCplus4_regI[3]), .B1(n144), .Y(
        n38) );
  AO22X2 U7 ( .A0(PCplus4[4]), .A1(n130), .B0(PCplus4_regI[4]), .B1(n144), .Y(
        n39) );
  AO22X2 U8 ( .A0(PCplus4[7]), .A1(n130), .B0(PCplus4_regI[7]), .B1(n144), .Y(
        n42) );
  AO22X2 U9 ( .A0(PCplus4[8]), .A1(n130), .B0(PCplus4_regI[8]), .B1(n144), .Y(
        n43) );
  AO22X2 U10 ( .A0(PCplus4[9]), .A1(n130), .B0(PCplus4_regI[9]), .B1(n144), 
        .Y(n44) );
  AO22X2 U11 ( .A0(PCplus4[10]), .A1(n130), .B0(PCplus4_regI[10]), .B1(n144), 
        .Y(n45) );
  AO22X2 U12 ( .A0(instruction_next[6]), .A1(n132), .B0(shamt[0]), .B1(n144), 
        .Y(n9) );
  AO22X2 U13 ( .A0(instruction_next[7]), .A1(n132), .B0(shamt[1]), .B1(n144), 
        .Y(n10) );
  AO22X2 U14 ( .A0(instruction_next[15]), .A1(n132), .B0(Rd[4]), .B1(n144), 
        .Y(n18) );
  AO22X2 U15 ( .A0(instruction_next[11]), .A1(n132), .B0(Rd[0]), .B1(n144), 
        .Y(n14) );
  AO22X2 U16 ( .A0(instruction_next[9]), .A1(n132), .B0(shamt[3]), .B1(n144), 
        .Y(n12) );
  AO22X1 U17 ( .A0(instruction_next[10]), .A1(n132), .B0(shamt[4]), .B1(n144), 
        .Y(n13) );
  AO22X2 U18 ( .A0(instruction_next[12]), .A1(n132), .B0(Rd[1]), .B1(n144), 
        .Y(n15) );
  AO22X2 U19 ( .A0(instruction_next[13]), .A1(n132), .B0(Rd[2]), .B1(n144), 
        .Y(n16) );
  BUFX20 U20 ( .A(n145), .Y(n132) );
  BUFX20 U21 ( .A(n145), .Y(n131) );
  INVX8 U22 ( .A(flush), .Y(n141) );
  NAND2X2 U23 ( .A(n1), .B(n141), .Y(n142) );
  BUFX20 U24 ( .A(n145), .Y(n130) );
  AO22XL U25 ( .A0(instruction_next[29]), .A1(n132), .B0(opcode[3]), .B1(n144), 
        .Y(n32) );
  OAI21XL U26 ( .A0(stall_lw_use), .A1(stallcache), .B0(n141), .Y(n1) );
  OAI21X4 U27 ( .A0(stall_lw_use), .A1(stallcache), .B0(n141), .Y(n143) );
  INVX20 U28 ( .A(n143), .Y(n144) );
  CLKBUFX2 U29 ( .A(shamt[4]), .Y(instruction_regI[10]) );
  CLKBUFX3 U30 ( .A(Rd[0]), .Y(instruction_regI[11]) );
  CLKBUFX3 U31 ( .A(Rd[1]), .Y(instruction_regI[12]) );
  CLKBUFX3 U32 ( .A(Rd[2]), .Y(instruction_regI[13]) );
  CLKBUFX3 U33 ( .A(Rd[3]), .Y(instruction_regI[14]) );
  CLKBUFX3 U34 ( .A(Rd[4]), .Y(instruction_regI[15]) );
  CLKBUFX3 U35 ( .A(shamt[0]), .Y(instruction_regI[6]) );
  CLKBUFX3 U36 ( .A(shamt[1]), .Y(instruction_regI[7]) );
  CLKBUFX3 U37 ( .A(shamt[2]), .Y(instruction_regI[8]) );
  CLKBUFX3 U38 ( .A(shamt[3]), .Y(instruction_regI[9]) );
  CLKBUFX2 U39 ( .A(opcode[4]), .Y(instruction_regI[30]) );
  CLKBUFX2 U40 ( .A(funct[3]), .Y(instruction_regI[3]) );
  CLKBUFX2 U41 ( .A(opcode[0]), .Y(instruction_regI[26]) );
  CLKBUFX2 U42 ( .A(Rt[2]), .Y(instruction_regI[18]) );
  CLKBUFX2 U43 ( .A(Rt[3]), .Y(instruction_regI[19]) );
  CLKBUFX2 U44 ( .A(Rs[2]), .Y(instruction_regI[23]) );
  CLKBUFX2 U45 ( .A(Rs[3]), .Y(instruction_regI[24]) );
  CLKBUFX2 U46 ( .A(funct[1]), .Y(instruction_regI[1]) );
  CLKBUFX2 U47 ( .A(funct[4]), .Y(instruction_regI[4]) );
  CLKBUFX2 U48 ( .A(funct[2]), .Y(instruction_regI[2]) );
  CLKBUFX2 U49 ( .A(funct[5]), .Y(instruction_regI[5]) );
  CLKBUFX2 U50 ( .A(opcode[5]), .Y(instruction_regI[31]) );
  CLKBUFX2 U51 ( .A(funct[0]), .Y(instruction_regI[0]) );
  CLKBUFX2 U52 ( .A(opcode[3]), .Y(instruction_regI[29]) );
  CLKBUFX2 U53 ( .A(opcode[2]), .Y(instruction_regI[28]) );
  CLKBUFX2 U54 ( .A(Rt[1]), .Y(instruction_regI[17]) );
  CLKBUFX2 U55 ( .A(Rt[0]), .Y(instruction_regI[16]) );
  CLKBUFX2 U56 ( .A(Rt[4]), .Y(instruction_regI[20]) );
  CLKBUFX2 U57 ( .A(Rs[0]), .Y(instruction_regI[21]) );
  CLKBUFX2 U58 ( .A(opcode[1]), .Y(instruction_regI[27]) );
  CLKBUFX2 U59 ( .A(Rs[1]), .Y(instruction_regI[22]) );
  CLKBUFX2 U60 ( .A(Rs[4]), .Y(instruction_regI[25]) );
  BUFX12 U61 ( .A(n145), .Y(n133) );
  AO22XL U62 ( .A0(instruction_next[22]), .A1(n133), .B0(Rs[1]), .B1(n144), 
        .Y(n25) );
  AO22XL U63 ( .A0(instruction_next[25]), .A1(n133), .B0(Rs[4]), .B1(n144), 
        .Y(n28) );
  AO22XL U64 ( .A0(instruction_next[27]), .A1(n133), .B0(opcode[1]), .B1(n144), 
        .Y(n30) );
  CLKBUFX2 U65 ( .A(rst_n), .Y(n134) );
  AO22XL U66 ( .A0(PCplus4[18]), .A1(n130), .B0(PCplus4_regI[18]), .B1(n144), 
        .Y(n53) );
  CLKBUFX2 U67 ( .A(funct[0]), .Y(immediate[0]) );
  CLKBUFX2 U68 ( .A(funct[0]), .Y(branchOffset[0]) );
  CLKBUFX3 U69 ( .A(n134), .Y(n135) );
  CLKBUFX3 U70 ( .A(n140), .Y(n136) );
  CLKBUFX3 U71 ( .A(n134), .Y(n137) );
  CLKBUFX3 U72 ( .A(n134), .Y(n138) );
  CLKBUFX3 U73 ( .A(n134), .Y(n139) );
  CLKBUFX3 U74 ( .A(n134), .Y(n140) );
  AO22XL U75 ( .A0(instruction_next[1]), .A1(n131), .B0(funct[1]), .B1(n144), 
        .Y(n4) );
  AO22XL U76 ( .A0(instruction_next[2]), .A1(n131), .B0(funct[2]), .B1(n144), 
        .Y(n5) );
  AO22XL U77 ( .A0(instruction_next[5]), .A1(n132), .B0(funct[5]), .B1(n144), 
        .Y(n8) );
  AO22XL U78 ( .A0(instruction_next[3]), .A1(n131), .B0(funct[3]), .B1(n144), 
        .Y(n6) );
  AO22XL U79 ( .A0(instruction_next[4]), .A1(n132), .B0(funct[4]), .B1(n144), 
        .Y(n7) );
  AO22XL U80 ( .A0(instruction_next[0]), .A1(n131), .B0(funct[0]), .B1(n144), 
        .Y(n3) );
  AO22XL U81 ( .A0(instruction_next[14]), .A1(n132), .B0(Rd[3]), .B1(n144), 
        .Y(n17) );
  AO22XL U82 ( .A0(instruction_next[8]), .A1(n132), .B0(shamt[2]), .B1(n144), 
        .Y(n11) );
  AO22XL U83 ( .A0(instruction_next[26]), .A1(n133), .B0(opcode[0]), .B1(n144), 
        .Y(n29) );
  AO22XL U84 ( .A0(instruction_next[16]), .A1(n133), .B0(Rt[0]), .B1(n144), 
        .Y(n19) );
  AO22XL U85 ( .A0(instruction_next[17]), .A1(n133), .B0(Rt[1]), .B1(n144), 
        .Y(n20) );
  AO22XL U86 ( .A0(instruction_next[18]), .A1(n133), .B0(Rt[2]), .B1(n144), 
        .Y(n21) );
  AO22XL U87 ( .A0(instruction_next[19]), .A1(n133), .B0(Rt[3]), .B1(n144), 
        .Y(n22) );
  AO22XL U88 ( .A0(instruction_next[20]), .A1(n133), .B0(Rt[4]), .B1(n144), 
        .Y(n23) );
  AO22XL U89 ( .A0(instruction_next[21]), .A1(n133), .B0(Rs[0]), .B1(n144), 
        .Y(n24) );
  AO22XL U90 ( .A0(instruction_next[23]), .A1(n133), .B0(Rs[2]), .B1(n144), 
        .Y(n26) );
  AO22XL U91 ( .A0(instruction_next[24]), .A1(n133), .B0(Rs[3]), .B1(n144), 
        .Y(n27) );
  AO22XL U92 ( .A0(PCplus4[2]), .A1(n130), .B0(PCplus4_regI[2]), .B1(n144), 
        .Y(n37) );
  AO22XL U93 ( .A0(PCplus4[5]), .A1(n130), .B0(PCplus4_regI[5]), .B1(n144), 
        .Y(n40) );
  AO22XL U94 ( .A0(PCplus4[6]), .A1(n130), .B0(PCplus4_regI[6]), .B1(n144), 
        .Y(n41) );
  AO22XL U95 ( .A0(PCplus4[11]), .A1(n130), .B0(PCplus4_regI[11]), .B1(n144), 
        .Y(n46) );
  AO22XL U96 ( .A0(PCplus4[12]), .A1(n132), .B0(PCplus4_regI[12]), .B1(n144), 
        .Y(n47) );
  AO22XL U97 ( .A0(PCplus4[13]), .A1(n131), .B0(PCplus4_regI[13]), .B1(n144), 
        .Y(n48) );
  AO22XL U98 ( .A0(PCplus4[14]), .A1(n130), .B0(PCplus4_regI[14]), .B1(n144), 
        .Y(n49) );
  AO22XL U99 ( .A0(PCplus4[15]), .A1(n132), .B0(PCplus4_regI[15]), .B1(n144), 
        .Y(n50) );
  AO22XL U100 ( .A0(PCplus4[16]), .A1(n131), .B0(PCplus4_regI[16]), .B1(n144), 
        .Y(n51) );
  AO22XL U101 ( .A0(PCplus4[17]), .A1(n130), .B0(PCplus4_regI[17]), .B1(n144), 
        .Y(n52) );
  AO22XL U102 ( .A0(PCplus4[19]), .A1(n132), .B0(PCplus4_regI[19]), .B1(n144), 
        .Y(n54) );
  AO22XL U103 ( .A0(PCplus4[20]), .A1(n131), .B0(PCplus4_regI[20]), .B1(n144), 
        .Y(n55) );
  AO22XL U104 ( .A0(PCplus4[21]), .A1(n130), .B0(PCplus4_regI[21]), .B1(n144), 
        .Y(n56) );
  AO22XL U105 ( .A0(PCplus4[22]), .A1(n132), .B0(PCplus4_regI[22]), .B1(n144), 
        .Y(n57) );
  AO22XL U106 ( .A0(PCplus4[23]), .A1(n131), .B0(PCplus4_regI[23]), .B1(n144), 
        .Y(n58) );
  AO22XL U107 ( .A0(PCplus4[24]), .A1(n131), .B0(PCplus4_regI[24]), .B1(n144), 
        .Y(n59) );
  AO22XL U108 ( .A0(PCplus4[25]), .A1(n131), .B0(PCplus4_regI[25]), .B1(n144), 
        .Y(n60) );
  AO22XL U109 ( .A0(PCplus4[26]), .A1(n131), .B0(PCplus4_regI[26]), .B1(n144), 
        .Y(n61) );
  AO22XL U110 ( .A0(PCplus4[27]), .A1(n131), .B0(PCplus4_regI[27]), .B1(n144), 
        .Y(n62) );
  AO22XL U111 ( .A0(PCplus4[28]), .A1(n131), .B0(PCplus4_regI[28]), .B1(n144), 
        .Y(n63) );
  AO22XL U112 ( .A0(PCplus4[29]), .A1(n131), .B0(PCplus4_regI[29]), .B1(n144), 
        .Y(n64) );
  AO22XL U113 ( .A0(PCplus4[30]), .A1(n131), .B0(PCplus4_regI[30]), .B1(n144), 
        .Y(n65) );
  AO22XL U114 ( .A0(PCplus4[31]), .A1(n131), .B0(PCplus4_regI[31]), .B1(n144), 
        .Y(n66) );
  CLKBUFX3 U115 ( .A(funct[1]), .Y(immediate[1]) );
  CLKBUFX3 U116 ( .A(funct[1]), .Y(branchOffset[1]) );
  CLKBUFX3 U117 ( .A(Rd[4]), .Y(immediate[15]) );
  CLKBUFX3 U118 ( .A(Rd[4]), .Y(branchOffset[15]) );
  CLKBUFX3 U119 ( .A(Rd[3]), .Y(immediate[14]) );
  CLKBUFX3 U120 ( .A(Rd[3]), .Y(branchOffset[14]) );
  CLKBUFX3 U121 ( .A(Rd[2]), .Y(immediate[13]) );
  CLKBUFX3 U122 ( .A(Rd[2]), .Y(branchOffset[13]) );
  CLKBUFX3 U123 ( .A(Rd[1]), .Y(immediate[12]) );
  CLKBUFX3 U124 ( .A(Rd[1]), .Y(branchOffset[12]) );
  CLKBUFX3 U125 ( .A(Rd[0]), .Y(immediate[11]) );
  CLKBUFX3 U126 ( .A(Rd[0]), .Y(branchOffset[11]) );
  CLKBUFX3 U127 ( .A(shamt[4]), .Y(immediate[10]) );
  CLKBUFX3 U128 ( .A(shamt[4]), .Y(branchOffset[10]) );
  CLKBUFX3 U129 ( .A(shamt[3]), .Y(immediate[9]) );
  CLKBUFX3 U130 ( .A(shamt[3]), .Y(branchOffset[9]) );
  CLKBUFX3 U131 ( .A(shamt[2]), .Y(immediate[8]) );
  CLKBUFX3 U132 ( .A(shamt[2]), .Y(branchOffset[8]) );
  CLKBUFX3 U133 ( .A(shamt[1]), .Y(immediate[7]) );
  CLKBUFX3 U134 ( .A(shamt[1]), .Y(branchOffset[7]) );
  CLKBUFX3 U135 ( .A(shamt[0]), .Y(immediate[6]) );
  CLKBUFX3 U136 ( .A(shamt[0]), .Y(branchOffset[6]) );
  CLKBUFX3 U137 ( .A(funct[5]), .Y(immediate[5]) );
  CLKBUFX3 U138 ( .A(funct[5]), .Y(branchOffset[5]) );
  CLKBUFX3 U139 ( .A(funct[4]), .Y(immediate[4]) );
  CLKBUFX3 U140 ( .A(funct[4]), .Y(branchOffset[4]) );
  CLKBUFX3 U141 ( .A(funct[3]), .Y(immediate[3]) );
  CLKBUFX3 U142 ( .A(funct[3]), .Y(branchOffset[3]) );
  CLKBUFX3 U143 ( .A(funct[2]), .Y(immediate[2]) );
  CLKBUFX3 U144 ( .A(funct[2]), .Y(branchOffset[2]) );
  AO22XL U145 ( .A0(instruction_next[30]), .A1(n130), .B0(opcode[4]), .B1(n144), .Y(n33) );
  AO22XL U146 ( .A0(instruction_next[31]), .A1(n131), .B0(opcode[5]), .B1(n144), .Y(n34) );
endmodule


module DEC_EX_regFile ( clk, rst_n, stallcache, MemtoReg, ALUOp, JumpReg, 
        MemRead, MemWrite, ALUsrc, RegWrite, Branch, PCplus4_regI, funct, 
        branchOffset_D, A, B, ExtOut, Rs, Rt, wsel, MemtoReg_regD, ALUOp_regD, 
        MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, funct_regD, 
        A_regD, B_regD, ExtOut_regD, Rs_regD, Rt_regD, wsel_regD, JumpReg_regD, 
        Branch_regD, PCplus4_regD, branchOffset_regD );
  input [1:0] MemtoReg;
  input [5:0] ALUOp;
  input [31:0] PCplus4_regI;
  input [5:0] funct;
  input [15:0] branchOffset_D;
  input [31:0] A;
  input [31:0] B;
  input [31:0] ExtOut;
  input [4:0] Rs;
  input [4:0] Rt;
  input [4:0] wsel;
  output [1:0] MemtoReg_regD;
  output [5:0] ALUOp_regD;
  output [5:0] funct_regD;
  output [31:0] A_regD;
  output [31:0] B_regD;
  output [31:0] ExtOut_regD;
  output [4:0] Rs_regD;
  output [4:0] Rt_regD;
  output [4:0] wsel_regD;
  output [31:0] PCplus4_regD;
  output [15:0] branchOffset_regD;
  input clk, rst_n, stallcache, JumpReg, MemRead, MemWrite, ALUsrc, RegWrite,
         Branch;
  output MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, JumpReg_regD,
         Branch_regD;
  wire   n2, n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n113, n114, n115, n116, n117, n118, n119, n122,
         n123, n124, n127, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n13, n111, n112, n120, n121, n125,
         n126, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440;

  DFFRX1 \MemtoReg_regD_reg[1]  ( .D(n300), .CK(clk), .RN(n146), .Q(
        MemtoReg_regD[1]) );
  DFFRX1 \MemtoReg_regD_reg[0]  ( .D(n299), .CK(clk), .RN(n146), .Q(
        MemtoReg_regD[0]) );
  DFFRX1 RegWrite_regD_reg ( .D(n290), .CK(clk), .RN(n145), .Q(RegWrite_regD)
         );
  DFFRX1 \wsel_regD_reg[4]  ( .D(n182), .CK(clk), .RN(n136), .Q(wsel_regD[4])
         );
  DFFRX1 \wsel_regD_reg[3]  ( .D(n181), .CK(clk), .RN(n136), .Q(wsel_regD[3])
         );
  DFFRX1 \wsel_regD_reg[2]  ( .D(n180), .CK(clk), .RN(n136), .Q(wsel_regD[2])
         );
  DFFRX1 \wsel_regD_reg[1]  ( .D(n179), .CK(clk), .RN(n136), .Q(wsel_regD[1])
         );
  DFFRX1 \wsel_regD_reg[0]  ( .D(n178), .CK(clk), .RN(n136), .Q(wsel_regD[0])
         );
  DFFRX1 \PCplus4_regD_reg[31]  ( .D(n354), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[31]) );
  DFFRX1 \funct_regD_reg[4]  ( .D(n305), .CK(clk), .RN(n146), .Q(funct_regD[4]) );
  DFFRX1 \branchOffset_regD_reg[11]  ( .D(n318), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[11]) );
  DFFRX1 \branchOffset_regD_reg[15]  ( .D(n322), .CK(clk), .RN(n148), .Q(
        branchOffset_regD[15]) );
  DFFRX1 \branchOffset_regD_reg[14]  ( .D(n321), .CK(clk), .RN(n148), .Q(
        branchOffset_regD[14]) );
  DFFRX1 \branchOffset_regD_reg[13]  ( .D(n320), .CK(clk), .RN(n148), .Q(
        branchOffset_regD[13]) );
  DFFRX1 \branchOffset_regD_reg[12]  ( .D(n319), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[12]) );
  DFFRX1 \branchOffset_regD_reg[10]  ( .D(n317), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[10]) );
  DFFRX1 \branchOffset_regD_reg[9]  ( .D(n316), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[9]) );
  DFFRX1 \branchOffset_regD_reg[8]  ( .D(n315), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[8]) );
  DFFRX1 \branchOffset_regD_reg[7]  ( .D(n314), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[7]) );
  DFFRX1 \branchOffset_regD_reg[5]  ( .D(n312), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[5]) );
  DFFRX1 \branchOffset_regD_reg[4]  ( .D(n311), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[4]) );
  DFFRX1 \branchOffset_regD_reg[3]  ( .D(n310), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[3]) );
  DFFRX1 \branchOffset_regD_reg[2]  ( .D(n309), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[2]) );
  DFFRX1 \branchOffset_regD_reg[1]  ( .D(n308), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[1]) );
  DFFRX1 \branchOffset_regD_reg[0]  ( .D(n307), .CK(clk), .RN(n146), .Q(
        branchOffset_regD[0]) );
  DFFRX1 \ExtOut_regD_reg[31]  ( .D(n224), .CK(clk), .RN(n140), .Q(
        ExtOut_regD[31]), .QN(n45) );
  DFFRX1 \ExtOut_regD_reg[29]  ( .D(n222), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[29]), .QN(n43) );
  DFFRX1 \ExtOut_regD_reg[30]  ( .D(n223), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[30]), .QN(n44) );
  DFFRX1 \ExtOut_regD_reg[7]  ( .D(n200), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[7]), .QN(n21) );
  DFFRX1 \ExtOut_regD_reg[24]  ( .D(n217), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[24]), .QN(n38) );
  DFFRX1 \ExtOut_regD_reg[10]  ( .D(n203), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[10]), .QN(n24) );
  DFFRX1 \ExtOut_regD_reg[14]  ( .D(n207), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[14]), .QN(n28) );
  DFFRX1 \ExtOut_regD_reg[18]  ( .D(n211), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[18]), .QN(n32) );
  DFFRX1 \ExtOut_regD_reg[20]  ( .D(n213), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[20]), .QN(n34) );
  DFFRX1 \ExtOut_regD_reg[21]  ( .D(n214), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[21]), .QN(n35) );
  DFFRX1 \ExtOut_regD_reg[16]  ( .D(n209), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[16]), .QN(n30) );
  DFFRX1 \ExtOut_regD_reg[11]  ( .D(n204), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[11]), .QN(n25) );
  DFFRX1 \ExtOut_regD_reg[22]  ( .D(n215), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[22]), .QN(n36) );
  DFFRX1 \ExtOut_regD_reg[8]  ( .D(n201), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[8]), .QN(n22) );
  DFFRX1 \ExtOut_regD_reg[25]  ( .D(n218), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[25]), .QN(n39) );
  DFFRX1 \ExtOut_regD_reg[17]  ( .D(n210), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[17]), .QN(n31) );
  DFFRX1 \ExtOut_regD_reg[13]  ( .D(n206), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[13]), .QN(n27) );
  DFFRX1 \ExtOut_regD_reg[9]  ( .D(n202), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[9]), .QN(n23) );
  DFFRX1 \ExtOut_regD_reg[23]  ( .D(n216), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[23]), .QN(n37) );
  DFFRX1 \ExtOut_regD_reg[27]  ( .D(n220), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[27]), .QN(n41) );
  DFFRX1 \ExtOut_regD_reg[19]  ( .D(n212), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[19]), .QN(n33) );
  DFFRX1 \ExtOut_regD_reg[6]  ( .D(n199), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[6]), .QN(n20) );
  DFFRX1 \ExtOut_regD_reg[1]  ( .D(n194), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[1]), .QN(n15) );
  DFFRX1 \ExtOut_regD_reg[2]  ( .D(n195), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[2]), .QN(n16) );
  DFFRX1 \ExtOut_regD_reg[26]  ( .D(n219), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[26]), .QN(n40) );
  DFFRX1 \ExtOut_regD_reg[12]  ( .D(n205), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[12]), .QN(n26) );
  DFFRX1 \ExtOut_regD_reg[4]  ( .D(n197), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[4]), .QN(n18) );
  DFFRX1 \ExtOut_regD_reg[15]  ( .D(n208), .CK(clk), .RN(n138), .Q(
        ExtOut_regD[15]), .QN(n29) );
  DFFRX1 \ExtOut_regD_reg[5]  ( .D(n198), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[5]), .QN(n19) );
  DFFRX1 \ExtOut_regD_reg[0]  ( .D(n193), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[0]), .QN(n14) );
  DFFRX1 \ExtOut_regD_reg[3]  ( .D(n196), .CK(clk), .RN(n137), .Q(
        ExtOut_regD[3]), .QN(n17) );
  DFFRX1 \ExtOut_regD_reg[28]  ( .D(n221), .CK(clk), .RN(n139), .Q(
        ExtOut_regD[28]), .QN(n42) );
  DFFRX1 \branchOffset_regD_reg[6]  ( .D(n313), .CK(clk), .RN(n147), .Q(
        branchOffset_regD[6]) );
  DFFRX1 \ALUOp_regD_reg[5]  ( .D(n298), .CK(clk), .RN(n146), .Q(ALUOp_regD[5]), .QN(n119) );
  DFFRX1 \PCplus4_regD_reg[16]  ( .D(n339), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[16]) );
  DFFRX1 \PCplus4_regD_reg[15]  ( .D(n338), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[15]) );
  DFFRX1 \PCplus4_regD_reg[14]  ( .D(n337), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[14]) );
  DFFRX1 \PCplus4_regD_reg[11]  ( .D(n334), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[11]) );
  DFFRX1 \PCplus4_regD_reg[1]  ( .D(n324), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[1]) );
  DFFRX1 \PCplus4_regD_reg[0]  ( .D(n323), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[0]) );
  DFFRX1 \PCplus4_regD_reg[27]  ( .D(n350), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[27]) );
  DFFRX1 \PCplus4_regD_reg[26]  ( .D(n349), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[26]) );
  DFFRX1 \PCplus4_regD_reg[25]  ( .D(n348), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[25]) );
  DFFRX1 \PCplus4_regD_reg[23]  ( .D(n346), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[23]) );
  DFFRX1 \PCplus4_regD_reg[22]  ( .D(n345), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[22]) );
  DFFRX1 \PCplus4_regD_reg[21]  ( .D(n344), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[21]) );
  DFFRX1 \PCplus4_regD_reg[20]  ( .D(n343), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[20]) );
  DFFRX1 \PCplus4_regD_reg[19]  ( .D(n342), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[19]) );
  DFFRX1 \PCplus4_regD_reg[18]  ( .D(n341), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[18]) );
  DFFRX1 \PCplus4_regD_reg[13]  ( .D(n336), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[13]) );
  DFFRX1 \PCplus4_regD_reg[12]  ( .D(n335), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[12]) );
  DFFRX1 \PCplus4_regD_reg[9]  ( .D(n332), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[9]) );
  DFFRX1 \PCplus4_regD_reg[7]  ( .D(n330), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[7]) );
  DFFRX1 \PCplus4_regD_reg[6]  ( .D(n329), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[6]) );
  DFFRX1 \PCplus4_regD_reg[5]  ( .D(n328), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[5]) );
  DFFRX1 \PCplus4_regD_reg[4]  ( .D(n327), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[4]) );
  DFFRX1 \PCplus4_regD_reg[3]  ( .D(n326), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[3]) );
  DFFRX1 \PCplus4_regD_reg[8]  ( .D(n331), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[8]) );
  DFFRX1 \funct_regD_reg[2]  ( .D(n303), .CK(clk), .RN(n146), .Q(funct_regD[2]), .QN(n124) );
  DFFRX1 \PCplus4_regD_reg[10]  ( .D(n333), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[10]) );
  DFFRX1 \PCplus4_regD_reg[24]  ( .D(n347), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[24]) );
  DFFRX1 \PCplus4_regD_reg[17]  ( .D(n340), .CK(clk), .RN(n149), .Q(
        PCplus4_regD[17]) );
  DFFRX1 \PCplus4_regD_reg[2]  ( .D(n325), .CK(clk), .RN(n148), .Q(
        PCplus4_regD[2]) );
  DFFRX1 \PCplus4_regD_reg[30]  ( .D(n353), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[30]) );
  DFFRX1 \PCplus4_regD_reg[29]  ( .D(n352), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[29]) );
  DFFRX1 \PCplus4_regD_reg[28]  ( .D(n351), .CK(clk), .RN(n150), .Q(
        PCplus4_regD[28]) );
  DFFRX1 \ALUOp_regD_reg[4]  ( .D(n297), .CK(clk), .RN(n146), .Q(ALUOp_regD[4]), .QN(n118) );
  DFFRX1 \ALUOp_regD_reg[0]  ( .D(n293), .CK(clk), .RN(n145), .Q(ALUOp_regD[0]), .QN(n114) );
  DFFRX1 \ALUOp_regD_reg[3]  ( .D(n296), .CK(clk), .RN(n146), .Q(ALUOp_regD[3]), .QN(n117) );
  DFFRX1 \ALUOp_regD_reg[2]  ( .D(n295), .CK(clk), .RN(n145), .Q(ALUOp_regD[2]), .QN(n116) );
  DFFRX1 \funct_regD_reg[5]  ( .D(n306), .CK(clk), .RN(n146), .Q(funct_regD[5]), .QN(n127) );
  DFFRX1 \funct_regD_reg[1]  ( .D(n302), .CK(clk), .RN(n146), .Q(funct_regD[1]), .QN(n123) );
  DFFRX1 \ALUOp_regD_reg[1]  ( .D(n294), .CK(clk), .RN(n145), .Q(ALUOp_regD[1]), .QN(n115) );
  DFFRX1 \B_regD_reg[16]  ( .D(n241), .CK(clk), .RN(n141), .Q(B_regD[16]), 
        .QN(n62) );
  DFFRX1 \B_regD_reg[20]  ( .D(n245), .CK(clk), .RN(n141), .Q(B_regD[20]), 
        .QN(n66) );
  DFFRX1 \B_regD_reg[13]  ( .D(n238), .CK(clk), .RN(n141), .Q(B_regD[13]), 
        .QN(n59) );
  DFFRX1 \B_regD_reg[17]  ( .D(n242), .CK(clk), .RN(n141), .Q(B_regD[17]), 
        .QN(n63) );
  DFFRX1 \B_regD_reg[9]  ( .D(n234), .CK(clk), .RN(n140), .Q(B_regD[9]), .QN(
        n55) );
  DFFRX1 \B_regD_reg[22]  ( .D(n247), .CK(clk), .RN(n141), .Q(B_regD[22]), 
        .QN(n68) );
  DFFRX1 \B_regD_reg[8]  ( .D(n233), .CK(clk), .RN(n140), .Q(B_regD[8]), .QN(
        n54) );
  DFFRX1 \B_regD_reg[14]  ( .D(n239), .CK(clk), .RN(n141), .Q(B_regD[14]), 
        .QN(n60) );
  DFFRX1 \B_regD_reg[21]  ( .D(n246), .CK(clk), .RN(n141), .Q(B_regD[21]), 
        .QN(n67) );
  DFFRX1 \B_regD_reg[12]  ( .D(n237), .CK(clk), .RN(n141), .Q(B_regD[12]), 
        .QN(n58) );
  DFFRX1 \B_regD_reg[10]  ( .D(n235), .CK(clk), .RN(n140), .Q(B_regD[10]), 
        .QN(n56) );
  DFFRX1 \B_regD_reg[23]  ( .D(n248), .CK(clk), .RN(n142), .Q(B_regD[23]), 
        .QN(n69) );
  DFFRX1 \B_regD_reg[11]  ( .D(n236), .CK(clk), .RN(n141), .Q(B_regD[11]), 
        .QN(n57) );
  DFFRX1 \B_regD_reg[15]  ( .D(n240), .CK(clk), .RN(n141), .Q(B_regD[15]), 
        .QN(n61) );
  DFFRX1 \A_regD_reg[16]  ( .D(n273), .CK(clk), .RN(n144), .Q(A_regD[16]), 
        .QN(n94) );
  DFFRX1 \A_regD_reg[20]  ( .D(n277), .CK(clk), .RN(n144), .Q(A_regD[20]), 
        .QN(n98) );
  DFFRX1 \A_regD_reg[13]  ( .D(n270), .CK(clk), .RN(n143), .Q(A_regD[13]), 
        .QN(n91) );
  DFFRX1 \A_regD_reg[12]  ( .D(n269), .CK(clk), .RN(n143), .Q(A_regD[12]), 
        .QN(n90) );
  DFFRX1 \A_regD_reg[15]  ( .D(n272), .CK(clk), .RN(n144), .Q(A_regD[15]), 
        .QN(n93) );
  DFFRX1 \A_regD_reg[17]  ( .D(n274), .CK(clk), .RN(n144), .Q(A_regD[17]), 
        .QN(n95) );
  DFFRX1 \A_regD_reg[8]  ( .D(n265), .CK(clk), .RN(n143), .Q(A_regD[8]), .QN(
        n86) );
  DFFRX1 \A_regD_reg[10]  ( .D(n267), .CK(clk), .RN(n143), .Q(A_regD[10]), 
        .QN(n88) );
  DFFRX1 \A_regD_reg[22]  ( .D(n279), .CK(clk), .RN(n144), .Q(A_regD[22]), 
        .QN(n100) );
  DFFRX1 \A_regD_reg[14]  ( .D(n271), .CK(clk), .RN(n143), .Q(A_regD[14]), 
        .QN(n92) );
  DFFRX1 \A_regD_reg[11]  ( .D(n268), .CK(clk), .RN(n143), .Q(A_regD[11]), 
        .QN(n89) );
  DFFRX1 \B_regD_reg[31]  ( .D(n256), .CK(clk), .RN(n142), .Q(B_regD[31]), 
        .QN(n77) );
  DFFRX1 \B_regD_reg[30]  ( .D(n255), .CK(clk), .RN(n142), .Q(B_regD[30]), 
        .QN(n76) );
  DFFRX1 \B_regD_reg[29]  ( .D(n254), .CK(clk), .RN(n142), .Q(B_regD[29]), 
        .QN(n75) );
  DFFRX1 \B_regD_reg[26]  ( .D(n251), .CK(clk), .RN(n142), .Q(B_regD[26]), 
        .QN(n72) );
  DFFRX1 \B_regD_reg[25]  ( .D(n250), .CK(clk), .RN(n142), .Q(B_regD[25]), 
        .QN(n71) );
  DFFRX1 \B_regD_reg[19]  ( .D(n244), .CK(clk), .RN(n141), .Q(B_regD[19]), 
        .QN(n65) );
  DFFRX1 \B_regD_reg[18]  ( .D(n243), .CK(clk), .RN(n141), .Q(B_regD[18]), 
        .QN(n64) );
  DFFRX1 \B_regD_reg[6]  ( .D(n231), .CK(clk), .RN(n140), .Q(B_regD[6]), .QN(
        n52) );
  DFFRX1 \A_regD_reg[23]  ( .D(n280), .CK(clk), .RN(n144), .Q(A_regD[23]), 
        .QN(n101) );
  DFFRX1 \A_regD_reg[21]  ( .D(n278), .CK(clk), .RN(n144), .Q(A_regD[21]), 
        .QN(n99) );
  DFFRX2 JumpReg_regD_reg ( .D(n177), .CK(clk), .RN(n136), .Q(JumpReg_regD), 
        .QN(n3) );
  DFFRX2 Branch_regD_reg ( .D(n176), .CK(clk), .RN(n136), .Q(Branch_regD), 
        .QN(n2) );
  DFFRX2 \funct_regD_reg[0]  ( .D(n301), .CK(clk), .RN(n146), .Q(funct_regD[0]), .QN(n122) );
  DFFRX1 MemRead_regD_reg ( .D(n292), .CK(clk), .RN(n145), .Q(MemRead_regD), 
        .QN(n113) );
  DFFRX1 \A_regD_reg[28]  ( .D(n285), .CK(clk), .RN(n145), .Q(A_regD[28]), 
        .QN(n106) );
  DFFRX1 \A_regD_reg[24]  ( .D(n281), .CK(clk), .RN(n144), .Q(A_regD[24]), 
        .QN(n102) );
  DFFRX1 \A_regD_reg[7]  ( .D(n264), .CK(clk), .RN(n143), .Q(A_regD[7]), .QN(
        n85) );
  DFFRX1 \A_regD_reg[2]  ( .D(n259), .CK(clk), .RN(n142), .Q(A_regD[2]), .QN(
        n80) );
  DFFRX1 \B_regD_reg[28]  ( .D(n253), .CK(clk), .RN(n142), .Q(B_regD[28]), 
        .QN(n74) );
  DFFRX1 \B_regD_reg[27]  ( .D(n252), .CK(clk), .RN(n142), .Q(B_regD[27]), 
        .QN(n73) );
  DFFRX1 \B_regD_reg[24]  ( .D(n249), .CK(clk), .RN(n142), .Q(B_regD[24]), 
        .QN(n70) );
  DFFRX1 \B_regD_reg[7]  ( .D(n232), .CK(clk), .RN(n140), .Q(B_regD[7]), .QN(
        n53) );
  DFFRX1 \B_regD_reg[5]  ( .D(n230), .CK(clk), .RN(n140), .Q(B_regD[5]), .QN(
        n51) );
  DFFRX1 \B_regD_reg[3]  ( .D(n228), .CK(clk), .RN(n140), .Q(B_regD[3]), .QN(
        n49) );
  DFFRX1 \B_regD_reg[2]  ( .D(n227), .CK(clk), .RN(n140), .Q(B_regD[2]), .QN(
        n48) );
  DFFRX1 \B_regD_reg[1]  ( .D(n226), .CK(clk), .RN(n140), .Q(B_regD[1]), .QN(
        n47) );
  DFFRX1 \B_regD_reg[0]  ( .D(n225), .CK(clk), .RN(n140), .Q(B_regD[0]), .QN(
        n46) );
  DFFRX1 \A_regD_reg[31]  ( .D(n288), .CK(clk), .RN(n145), .Q(A_regD[31]), 
        .QN(n109) );
  DFFRX1 \A_regD_reg[30]  ( .D(n287), .CK(clk), .RN(n145), .Q(A_regD[30]), 
        .QN(n108) );
  DFFRX1 \A_regD_reg[29]  ( .D(n286), .CK(clk), .RN(n145), .Q(A_regD[29]), 
        .QN(n107) );
  DFFRX1 \A_regD_reg[27]  ( .D(n284), .CK(clk), .RN(n145), .Q(A_regD[27]), 
        .QN(n105) );
  DFFRX1 \A_regD_reg[26]  ( .D(n283), .CK(clk), .RN(n144), .Q(A_regD[26]), 
        .QN(n104) );
  DFFRX1 \A_regD_reg[25]  ( .D(n282), .CK(clk), .RN(n144), .Q(A_regD[25]), 
        .QN(n103) );
  DFFRX1 \A_regD_reg[19]  ( .D(n276), .CK(clk), .RN(n144), .Q(A_regD[19]), 
        .QN(n97) );
  DFFRX1 \A_regD_reg[18]  ( .D(n275), .CK(clk), .RN(n144), .Q(A_regD[18]), 
        .QN(n96) );
  DFFRX1 \A_regD_reg[9]  ( .D(n266), .CK(clk), .RN(n143), .Q(A_regD[9]), .QN(
        n87) );
  DFFRX1 \A_regD_reg[6]  ( .D(n263), .CK(clk), .RN(n143), .Q(A_regD[6]), .QN(
        n84) );
  DFFRX1 \A_regD_reg[5]  ( .D(n262), .CK(clk), .RN(n143), .Q(A_regD[5]), .QN(
        n83) );
  DFFRX1 \A_regD_reg[4]  ( .D(n261), .CK(clk), .RN(n143), .Q(A_regD[4]), .QN(
        n82) );
  DFFRX1 \A_regD_reg[3]  ( .D(n260), .CK(clk), .RN(n143), .Q(A_regD[3]), .QN(
        n81) );
  DFFRX1 \A_regD_reg[1]  ( .D(n258), .CK(clk), .RN(n142), .Q(A_regD[1]), .QN(
        n79) );
  DFFRX1 \A_regD_reg[0]  ( .D(n257), .CK(clk), .RN(n142), .Q(A_regD[0]), .QN(
        n78) );
  DFFRX2 \B_regD_reg[4]  ( .D(n229), .CK(clk), .RN(n140), .Q(B_regD[4]), .QN(
        n50) );
  DFFRHQX8 \Rs_regD_reg[4]  ( .D(n192), .CK(clk), .RN(n137), .Q(Rs_regD[4]) );
  DFFRHQX8 \Rs_regD_reg[2]  ( .D(n190), .CK(clk), .RN(n137), .Q(Rs_regD[2]) );
  DFFRHQX8 \Rt_regD_reg[2]  ( .D(n185), .CK(clk), .RN(n136), .Q(Rt_regD[2]) );
  DFFRHQX8 \Rs_regD_reg[3]  ( .D(n191), .CK(clk), .RN(n137), .Q(Rs_regD[3]) );
  DFFRHQX8 \Rs_regD_reg[1]  ( .D(n189), .CK(clk), .RN(n137), .Q(Rs_regD[1]) );
  DFFRHQX8 \Rs_regD_reg[0]  ( .D(n188), .CK(clk), .RN(n137), .Q(Rs_regD[0]) );
  DFFRHQX8 \Rt_regD_reg[3]  ( .D(n186), .CK(clk), .RN(n136), .Q(Rt_regD[3]) );
  DFFRHQX8 \Rt_regD_reg[4]  ( .D(n187), .CK(clk), .RN(n136), .Q(Rt_regD[4]) );
  DFFRHQX8 \Rt_regD_reg[1]  ( .D(n184), .CK(clk), .RN(n136), .Q(Rt_regD[1]) );
  DFFRHQX8 \Rt_regD_reg[0]  ( .D(n183), .CK(clk), .RN(n136), .Q(Rt_regD[0]) );
  DFFRX1 MemWrite_regD_reg ( .D(n291), .CK(clk), .RN(rst_n), .Q(MemWrite_regD)
         );
  DFFRX1 \funct_regD_reg[3]  ( .D(n304), .CK(clk), .RN(rst_n), .Q(
        funct_regD[3]) );
  DFFRX4 ALUsrc_regD_reg ( .D(n289), .CK(clk), .RN(n145), .Q(ALUsrc_regD), 
        .QN(n110) );
  CLKMX2X2 U2 ( .A(Rs[4]), .B(Rs_regD[4]), .S0(n128), .Y(n192) );
  CLKMX2X2 U3 ( .A(A[0]), .B(n397), .S0(n125), .Y(n257) );
  CLKMX2X2 U4 ( .A(A[26]), .B(n423), .S0(n128), .Y(n283) );
  CLKMX2X2 U5 ( .A(B[15]), .B(n380), .S0(n121), .Y(n240) );
  CLKMX2X2 U6 ( .A(B[11]), .B(n376), .S0(n121), .Y(n236) );
  CLKMX2X2 U7 ( .A(B[10]), .B(n375), .S0(n121), .Y(n235) );
  MX2X1 U8 ( .A(B[12]), .B(n377), .S0(n121), .Y(n237) );
  CLKMX2X2 U9 ( .A(B[14]), .B(n379), .S0(n121), .Y(n239) );
  CLKMX2X2 U10 ( .A(B[13]), .B(n378), .S0(n121), .Y(n238) );
  BUFX8 U11 ( .A(n132), .Y(n131) );
  BUFX4 U12 ( .A(n13), .Y(n133) );
  BUFX8 U13 ( .A(n133), .Y(n132) );
  BUFX20 U14 ( .A(n130), .Y(n125) );
  CLKBUFX6 U15 ( .A(n134), .Y(n130) );
  CLKMX2X3 U16 ( .A(B[30]), .B(n395), .S0(n125), .Y(n255) );
  CLKMX2X2 U17 ( .A(ExtOut[9]), .B(n163), .S0(n111), .Y(n202) );
  CLKMX2X2 U18 ( .A(funct[3]), .B(funct_regD[3]), .S0(n128), .Y(n304) );
  CLKMX2X2 U19 ( .A(funct[1]), .B(n430), .S0(n111), .Y(n302) );
  CLKMX2X2 U20 ( .A(funct[2]), .B(n431), .S0(n128), .Y(n303) );
  CLKMX2X2 U21 ( .A(funct[4]), .B(funct_regD[4]), .S0(n111), .Y(n305) );
  CLKMX2X2 U22 ( .A(funct[5]), .B(n432), .S0(n128), .Y(n306) );
  CLKMX2X2 U23 ( .A(A[27]), .B(n424), .S0(n128), .Y(n284) );
  CLKMX2X2 U24 ( .A(A[28]), .B(n425), .S0(n128), .Y(n285) );
  CLKMX2X2 U25 ( .A(A[29]), .B(n426), .S0(n128), .Y(n286) );
  CLKMX2X2 U26 ( .A(A[30]), .B(n427), .S0(n128), .Y(n287) );
  CLKMX2X2 U27 ( .A(A[31]), .B(n428), .S0(n128), .Y(n288) );
  BUFX20 U28 ( .A(n132), .Y(n111) );
  CLKBUFX4 U29 ( .A(n13), .Y(n134) );
  BUFX20 U30 ( .A(n131), .Y(n112) );
  BUFX20 U31 ( .A(n131), .Y(n120) );
  BUFX20 U32 ( .A(n129), .Y(n128) );
  CLKBUFX4 U33 ( .A(n134), .Y(n129) );
  CLKBUFX4 U34 ( .A(n129), .Y(n126) );
  MX2X1 U35 ( .A(A[1]), .B(n398), .S0(n126), .Y(n258) );
  CLKMX2X2 U36 ( .A(A[2]), .B(n399), .S0(n126), .Y(n259) );
  CLKMX2X2 U37 ( .A(A[3]), .B(n400), .S0(n126), .Y(n260) );
  CLKMX2X2 U38 ( .A(A[4]), .B(n401), .S0(n126), .Y(n261) );
  CLKMX2X2 U39 ( .A(A[5]), .B(n402), .S0(n126), .Y(n262) );
  CLKMX2X2 U40 ( .A(A[6]), .B(n403), .S0(n126), .Y(n263) );
  CLKMX2X2 U41 ( .A(A[7]), .B(n404), .S0(n126), .Y(n264) );
  CLKMX2X2 U42 ( .A(A[8]), .B(n405), .S0(n126), .Y(n265) );
  CLKMX2X2 U43 ( .A(A[9]), .B(n406), .S0(n126), .Y(n266) );
  CLKBUFX4 U44 ( .A(n130), .Y(n121) );
  CLKMX2X2 U45 ( .A(B[9]), .B(n374), .S0(n121), .Y(n234) );
  CLKMX2X4 U46 ( .A(B[21]), .B(n386), .S0(n125), .Y(n246) );
  MX2X2 U47 ( .A(B[22]), .B(n387), .S0(n125), .Y(n247) );
  MX2X2 U48 ( .A(B[23]), .B(n388), .S0(n125), .Y(n248) );
  MX2X2 U49 ( .A(B[24]), .B(n389), .S0(n125), .Y(n249) );
  MX2X2 U50 ( .A(B[25]), .B(n390), .S0(n125), .Y(n250) );
  MX2X2 U51 ( .A(B[26]), .B(n391), .S0(n125), .Y(n251) );
  MX2X2 U52 ( .A(B[27]), .B(n392), .S0(n125), .Y(n252) );
  MX2X2 U53 ( .A(B[28]), .B(n393), .S0(n125), .Y(n253) );
  MX2X2 U54 ( .A(B[29]), .B(n394), .S0(n125), .Y(n254) );
  CLKMX2X2 U55 ( .A(ALUsrc), .B(n433), .S0(n128), .Y(n289) );
  CLKBUFX2 U56 ( .A(rst_n), .Y(n135) );
  MX2XL U57 ( .A(Branch), .B(n152), .S0(n132), .Y(n176) );
  MX2XL U58 ( .A(ExtOut[0]), .B(n154), .S0(n132), .Y(n193) );
  MX2XL U59 ( .A(ExtOut[13]), .B(n167), .S0(n112), .Y(n206) );
  MX2XL U60 ( .A(ExtOut[26]), .B(n359), .S0(n120), .Y(n219) );
  MX2XL U61 ( .A(B[7]), .B(n372), .S0(n121), .Y(n232) );
  MX2XL U62 ( .A(A[14]), .B(n411), .S0(n128), .Y(n271) );
  MX2XL U63 ( .A(branchOffset_D[0]), .B(branchOffset_regD[0]), .S0(n111), .Y(
        n307) );
  MX2XL U64 ( .A(branchOffset_D[13]), .B(branchOffset_regD[13]), .S0(n111), 
        .Y(n320) );
  MX2XL U65 ( .A(PCplus4_regI[10]), .B(PCplus4_regD[10]), .S0(n125), .Y(n333)
         );
  MX2XL U66 ( .A(MemtoReg[1]), .B(MemtoReg_regD[1]), .S0(n125), .Y(n300) );
  CLKBUFX3 U67 ( .A(n151), .Y(n137) );
  CLKBUFX3 U68 ( .A(n151), .Y(n138) );
  CLKBUFX3 U69 ( .A(n135), .Y(n139) );
  CLKBUFX3 U70 ( .A(n151), .Y(n140) );
  CLKBUFX3 U71 ( .A(n135), .Y(n141) );
  CLKBUFX3 U72 ( .A(n151), .Y(n142) );
  CLKBUFX3 U73 ( .A(n135), .Y(n143) );
  CLKBUFX3 U74 ( .A(n135), .Y(n144) );
  CLKBUFX3 U75 ( .A(n151), .Y(n145) );
  CLKBUFX3 U76 ( .A(n151), .Y(n146) );
  CLKBUFX3 U77 ( .A(n135), .Y(n147) );
  CLKBUFX3 U78 ( .A(n151), .Y(n148) );
  CLKBUFX3 U79 ( .A(n135), .Y(n149) );
  CLKBUFX3 U80 ( .A(n151), .Y(n150) );
  CLKBUFX3 U81 ( .A(n135), .Y(n136) );
  CLKBUFX3 U82 ( .A(n135), .Y(n151) );
  CLKINVX1 U83 ( .A(n123), .Y(n430) );
  MX2XL U84 ( .A(funct[0]), .B(n429), .S0(n128), .Y(n301) );
  CLKINVX1 U85 ( .A(n122), .Y(n429) );
  MX2XL U86 ( .A(MemtoReg[0]), .B(MemtoReg_regD[0]), .S0(n125), .Y(n299) );
  MX2XL U87 ( .A(MemWrite), .B(MemWrite_regD), .S0(n128), .Y(n291) );
  MX2XL U88 ( .A(MemRead), .B(n434), .S0(n128), .Y(n292) );
  CLKINVX1 U89 ( .A(n113), .Y(n434) );
  MX2XL U90 ( .A(ALUOp[0]), .B(n435), .S0(n125), .Y(n293) );
  CLKINVX1 U91 ( .A(n114), .Y(n435) );
  MX2XL U92 ( .A(ALUOp[1]), .B(n436), .S0(n125), .Y(n294) );
  CLKINVX1 U93 ( .A(n115), .Y(n436) );
  MX2XL U94 ( .A(ALUOp[2]), .B(n437), .S0(n128), .Y(n295) );
  CLKINVX1 U95 ( .A(n116), .Y(n437) );
  MX2XL U96 ( .A(ALUOp[3]), .B(n438), .S0(n125), .Y(n296) );
  CLKINVX1 U97 ( .A(n117), .Y(n438) );
  MX2XL U98 ( .A(ALUOp[4]), .B(n439), .S0(n128), .Y(n297) );
  CLKINVX1 U99 ( .A(n118), .Y(n439) );
  MX2XL U100 ( .A(ALUOp[5]), .B(n440), .S0(n131), .Y(n298) );
  CLKINVX1 U101 ( .A(n119), .Y(n440) );
  MX2XL U102 ( .A(Rs[0]), .B(Rs_regD[0]), .S0(n125), .Y(n188) );
  MX2XL U103 ( .A(Rs[1]), .B(Rs_regD[1]), .S0(n128), .Y(n189) );
  MX2XL U104 ( .A(Rs[2]), .B(Rs_regD[2]), .S0(n125), .Y(n190) );
  MX2XL U105 ( .A(Rs[3]), .B(Rs_regD[3]), .S0(n128), .Y(n191) );
  CLKINVX1 U106 ( .A(n2), .Y(n152) );
  MX2XL U107 ( .A(JumpReg), .B(n153), .S0(n125), .Y(n177) );
  CLKINVX1 U108 ( .A(n3), .Y(n153) );
  MX2XL U109 ( .A(wsel[0]), .B(wsel_regD[0]), .S0(n132), .Y(n178) );
  MX2XL U110 ( .A(wsel[1]), .B(wsel_regD[1]), .S0(n132), .Y(n179) );
  MX2XL U111 ( .A(wsel[2]), .B(wsel_regD[2]), .S0(n132), .Y(n180) );
  MX2XL U112 ( .A(wsel[3]), .B(wsel_regD[3]), .S0(n132), .Y(n181) );
  MX2XL U113 ( .A(wsel[4]), .B(wsel_regD[4]), .S0(n132), .Y(n182) );
  MX2XL U114 ( .A(Rt[0]), .B(Rt_regD[0]), .S0(n125), .Y(n183) );
  MX2XL U115 ( .A(Rt[1]), .B(Rt_regD[1]), .S0(n128), .Y(n184) );
  MX2XL U116 ( .A(Rt[2]), .B(Rt_regD[2]), .S0(n125), .Y(n185) );
  MX2XL U117 ( .A(Rt[3]), .B(Rt_regD[3]), .S0(n128), .Y(n186) );
  MX2XL U118 ( .A(Rt[4]), .B(Rt_regD[4]), .S0(n125), .Y(n187) );
  CLKINVX1 U119 ( .A(n14), .Y(n154) );
  MX2XL U120 ( .A(ExtOut[1]), .B(n155), .S0(n132), .Y(n194) );
  CLKINVX1 U121 ( .A(n15), .Y(n155) );
  MX2XL U122 ( .A(ExtOut[2]), .B(n156), .S0(n132), .Y(n195) );
  CLKINVX1 U123 ( .A(n16), .Y(n156) );
  MX2XL U124 ( .A(ExtOut[3]), .B(n157), .S0(n132), .Y(n196) );
  CLKINVX1 U125 ( .A(n17), .Y(n157) );
  MX2XL U126 ( .A(ExtOut[4]), .B(n158), .S0(n125), .Y(n197) );
  CLKINVX1 U127 ( .A(n18), .Y(n158) );
  MX2XL U128 ( .A(ExtOut[5]), .B(n159), .S0(n132), .Y(n198) );
  CLKINVX1 U129 ( .A(n19), .Y(n159) );
  MX2XL U130 ( .A(ExtOut[6]), .B(n160), .S0(n128), .Y(n199) );
  CLKINVX1 U131 ( .A(n20), .Y(n160) );
  MX2XL U132 ( .A(ExtOut[7]), .B(n161), .S0(n125), .Y(n200) );
  CLKINVX1 U133 ( .A(n21), .Y(n161) );
  MX2XL U134 ( .A(ExtOut[8]), .B(n162), .S0(n128), .Y(n201) );
  CLKINVX1 U135 ( .A(n22), .Y(n162) );
  CLKINVX1 U136 ( .A(n23), .Y(n163) );
  MX2XL U137 ( .A(ExtOut[10]), .B(n164), .S0(n125), .Y(n203) );
  CLKINVX1 U138 ( .A(n24), .Y(n164) );
  MX2XL U139 ( .A(ExtOut[11]), .B(n165), .S0(n128), .Y(n204) );
  CLKINVX1 U140 ( .A(n25), .Y(n165) );
  MX2XL U141 ( .A(ExtOut[12]), .B(n166), .S0(n132), .Y(n205) );
  CLKINVX1 U142 ( .A(n26), .Y(n166) );
  CLKINVX1 U143 ( .A(n27), .Y(n167) );
  MX2XL U144 ( .A(ExtOut[14]), .B(n168), .S0(n112), .Y(n207) );
  CLKINVX1 U145 ( .A(n28), .Y(n168) );
  MX2XL U146 ( .A(ExtOut[15]), .B(n169), .S0(n112), .Y(n208) );
  CLKINVX1 U147 ( .A(n29), .Y(n169) );
  MX2XL U148 ( .A(ExtOut[16]), .B(n170), .S0(n112), .Y(n209) );
  CLKINVX1 U149 ( .A(n30), .Y(n170) );
  MX2XL U150 ( .A(ExtOut[17]), .B(n171), .S0(n112), .Y(n210) );
  CLKINVX1 U151 ( .A(n31), .Y(n171) );
  MX2XL U152 ( .A(ExtOut[18]), .B(n172), .S0(n112), .Y(n211) );
  CLKINVX1 U153 ( .A(n32), .Y(n172) );
  MX2XL U154 ( .A(ExtOut[19]), .B(n173), .S0(n112), .Y(n212) );
  CLKINVX1 U155 ( .A(n33), .Y(n173) );
  MX2XL U156 ( .A(ExtOut[20]), .B(n174), .S0(n112), .Y(n213) );
  CLKINVX1 U157 ( .A(n34), .Y(n174) );
  MX2XL U158 ( .A(ExtOut[21]), .B(n175), .S0(n112), .Y(n214) );
  CLKINVX1 U159 ( .A(n35), .Y(n175) );
  MX2XL U160 ( .A(ExtOut[22]), .B(n355), .S0(n112), .Y(n215) );
  CLKINVX1 U161 ( .A(n36), .Y(n355) );
  MX2XL U162 ( .A(ExtOut[23]), .B(n356), .S0(n112), .Y(n216) );
  CLKINVX1 U163 ( .A(n37), .Y(n356) );
  MX2XL U164 ( .A(ExtOut[24]), .B(n357), .S0(n112), .Y(n217) );
  CLKINVX1 U165 ( .A(n38), .Y(n357) );
  MX2XL U166 ( .A(ExtOut[25]), .B(n358), .S0(n112), .Y(n218) );
  CLKINVX1 U167 ( .A(n39), .Y(n358) );
  CLKINVX1 U168 ( .A(n40), .Y(n359) );
  MX2XL U169 ( .A(ExtOut[27]), .B(n360), .S0(n120), .Y(n220) );
  CLKINVX1 U170 ( .A(n41), .Y(n360) );
  MX2XL U171 ( .A(ExtOut[28]), .B(n361), .S0(n120), .Y(n221) );
  CLKINVX1 U172 ( .A(n42), .Y(n361) );
  MX2XL U173 ( .A(ExtOut[29]), .B(n362), .S0(n120), .Y(n222) );
  CLKINVX1 U174 ( .A(n43), .Y(n362) );
  MX2XL U175 ( .A(ExtOut[30]), .B(n363), .S0(n120), .Y(n223) );
  CLKINVX1 U176 ( .A(n44), .Y(n363) );
  MX2XL U177 ( .A(ExtOut[31]), .B(n364), .S0(n120), .Y(n224) );
  CLKINVX1 U178 ( .A(n45), .Y(n364) );
  MX2XL U179 ( .A(B[0]), .B(n365), .S0(n120), .Y(n225) );
  CLKINVX1 U180 ( .A(n46), .Y(n365) );
  MX2XL U181 ( .A(B[1]), .B(n366), .S0(n120), .Y(n226) );
  CLKINVX1 U182 ( .A(n47), .Y(n366) );
  MX2XL U183 ( .A(B[2]), .B(n367), .S0(n120), .Y(n227) );
  CLKINVX1 U184 ( .A(n48), .Y(n367) );
  MX2XL U185 ( .A(B[3]), .B(n368), .S0(n120), .Y(n228) );
  CLKINVX1 U186 ( .A(n49), .Y(n368) );
  MX2XL U187 ( .A(B[4]), .B(n369), .S0(n120), .Y(n229) );
  CLKINVX1 U188 ( .A(n50), .Y(n369) );
  MX2XL U189 ( .A(B[5]), .B(n370), .S0(n120), .Y(n230) );
  CLKINVX1 U190 ( .A(n51), .Y(n370) );
  MX2XL U191 ( .A(B[6]), .B(n371), .S0(n120), .Y(n231) );
  CLKINVX1 U192 ( .A(n52), .Y(n371) );
  CLKINVX1 U193 ( .A(n53), .Y(n372) );
  MX2XL U194 ( .A(B[8]), .B(n373), .S0(n121), .Y(n233) );
  CLKINVX1 U195 ( .A(n54), .Y(n373) );
  CLKINVX1 U196 ( .A(n55), .Y(n374) );
  CLKINVX1 U197 ( .A(n56), .Y(n375) );
  CLKINVX1 U198 ( .A(n57), .Y(n376) );
  CLKINVX1 U199 ( .A(n58), .Y(n377) );
  CLKINVX1 U200 ( .A(n59), .Y(n378) );
  CLKINVX1 U201 ( .A(n60), .Y(n379) );
  CLKINVX1 U202 ( .A(n61), .Y(n380) );
  MX2XL U203 ( .A(B[16]), .B(n381), .S0(n121), .Y(n241) );
  CLKINVX1 U204 ( .A(n62), .Y(n381) );
  MX2XL U205 ( .A(B[17]), .B(n382), .S0(n121), .Y(n242) );
  CLKINVX1 U206 ( .A(n63), .Y(n382) );
  MX2XL U207 ( .A(B[18]), .B(n383), .S0(n121), .Y(n243) );
  CLKINVX1 U208 ( .A(n64), .Y(n383) );
  MX2XL U209 ( .A(B[19]), .B(n384), .S0(n121), .Y(n244) );
  CLKINVX1 U210 ( .A(n65), .Y(n384) );
  CLKMX2X2 U211 ( .A(B[20]), .B(n385), .S0(n125), .Y(n245) );
  CLKINVX1 U212 ( .A(n66), .Y(n385) );
  CLKINVX1 U213 ( .A(n67), .Y(n386) );
  CLKINVX1 U214 ( .A(n68), .Y(n387) );
  CLKINVX1 U215 ( .A(n69), .Y(n388) );
  CLKINVX1 U216 ( .A(n70), .Y(n389) );
  CLKINVX1 U217 ( .A(n71), .Y(n390) );
  CLKINVX1 U218 ( .A(n72), .Y(n391) );
  CLKINVX1 U219 ( .A(n73), .Y(n392) );
  CLKINVX1 U220 ( .A(n74), .Y(n393) );
  CLKINVX1 U221 ( .A(n75), .Y(n394) );
  CLKINVX1 U222 ( .A(n76), .Y(n395) );
  MX2XL U223 ( .A(B[31]), .B(n396), .S0(n125), .Y(n256) );
  CLKINVX1 U224 ( .A(n77), .Y(n396) );
  CLKINVX1 U225 ( .A(n78), .Y(n397) );
  CLKINVX1 U226 ( .A(n79), .Y(n398) );
  CLKINVX1 U227 ( .A(n80), .Y(n399) );
  CLKINVX1 U228 ( .A(n81), .Y(n400) );
  CLKINVX1 U229 ( .A(n82), .Y(n401) );
  CLKINVX1 U230 ( .A(n83), .Y(n402) );
  CLKINVX1 U231 ( .A(n84), .Y(n403) );
  CLKINVX1 U232 ( .A(n85), .Y(n404) );
  CLKINVX1 U233 ( .A(n86), .Y(n405) );
  CLKINVX1 U234 ( .A(n87), .Y(n406) );
  MX2XL U235 ( .A(A[10]), .B(n407), .S0(n126), .Y(n267) );
  CLKINVX1 U236 ( .A(n88), .Y(n407) );
  MX2XL U237 ( .A(A[11]), .B(n408), .S0(n126), .Y(n268) );
  CLKINVX1 U238 ( .A(n89), .Y(n408) );
  MX2XL U239 ( .A(A[12]), .B(n409), .S0(n126), .Y(n269) );
  CLKINVX1 U240 ( .A(n90), .Y(n409) );
  MX2XL U241 ( .A(A[13]), .B(n410), .S0(n126), .Y(n270) );
  CLKINVX1 U242 ( .A(n91), .Y(n410) );
  CLKINVX1 U243 ( .A(n92), .Y(n411) );
  MX2XL U244 ( .A(A[15]), .B(n412), .S0(n128), .Y(n272) );
  CLKINVX1 U245 ( .A(n93), .Y(n412) );
  MX2XL U246 ( .A(A[16]), .B(n413), .S0(n128), .Y(n273) );
  CLKINVX1 U247 ( .A(n94), .Y(n413) );
  MX2XL U248 ( .A(A[17]), .B(n414), .S0(n128), .Y(n274) );
  CLKINVX1 U249 ( .A(n95), .Y(n414) );
  MX2XL U250 ( .A(A[18]), .B(n415), .S0(n128), .Y(n275) );
  CLKINVX1 U251 ( .A(n96), .Y(n415) );
  MX2XL U252 ( .A(A[19]), .B(n416), .S0(n128), .Y(n276) );
  CLKINVX1 U253 ( .A(n97), .Y(n416) );
  MX2XL U254 ( .A(A[20]), .B(n417), .S0(n128), .Y(n277) );
  CLKINVX1 U255 ( .A(n98), .Y(n417) );
  MX2XL U256 ( .A(A[21]), .B(n418), .S0(n128), .Y(n278) );
  CLKINVX1 U257 ( .A(n99), .Y(n418) );
  MX2XL U258 ( .A(A[22]), .B(n419), .S0(n128), .Y(n279) );
  CLKINVX1 U259 ( .A(n100), .Y(n419) );
  MX2XL U260 ( .A(A[23]), .B(n420), .S0(n128), .Y(n280) );
  CLKINVX1 U261 ( .A(n101), .Y(n420) );
  MX2XL U262 ( .A(A[24]), .B(n421), .S0(n128), .Y(n281) );
  CLKINVX1 U263 ( .A(n102), .Y(n421) );
  MX2XL U264 ( .A(A[25]), .B(n422), .S0(n128), .Y(n282) );
  CLKINVX1 U265 ( .A(n103), .Y(n422) );
  CLKINVX1 U266 ( .A(n104), .Y(n423) );
  MX2XL U267 ( .A(branchOffset_D[1]), .B(branchOffset_regD[1]), .S0(n111), .Y(
        n308) );
  MX2XL U268 ( .A(branchOffset_D[2]), .B(branchOffset_regD[2]), .S0(n111), .Y(
        n309) );
  MX2XL U269 ( .A(branchOffset_D[3]), .B(branchOffset_regD[3]), .S0(n111), .Y(
        n310) );
  MX2XL U270 ( .A(branchOffset_D[4]), .B(branchOffset_regD[4]), .S0(n111), .Y(
        n311) );
  MX2XL U271 ( .A(branchOffset_D[5]), .B(branchOffset_regD[5]), .S0(n111), .Y(
        n312) );
  MX2XL U272 ( .A(branchOffset_D[6]), .B(branchOffset_regD[6]), .S0(n111), .Y(
        n313) );
  MX2XL U273 ( .A(branchOffset_D[7]), .B(branchOffset_regD[7]), .S0(n111), .Y(
        n314) );
  MX2XL U274 ( .A(branchOffset_D[8]), .B(branchOffset_regD[8]), .S0(n111), .Y(
        n315) );
  MX2XL U275 ( .A(branchOffset_D[9]), .B(branchOffset_regD[9]), .S0(n111), .Y(
        n316) );
  MX2XL U276 ( .A(branchOffset_D[10]), .B(branchOffset_regD[10]), .S0(n111), 
        .Y(n317) );
  MX2XL U277 ( .A(branchOffset_D[11]), .B(branchOffset_regD[11]), .S0(n111), 
        .Y(n318) );
  MX2XL U278 ( .A(branchOffset_D[12]), .B(branchOffset_regD[12]), .S0(n111), 
        .Y(n319) );
  MX2XL U279 ( .A(branchOffset_D[14]), .B(branchOffset_regD[14]), .S0(n111), 
        .Y(n321) );
  MX2XL U280 ( .A(branchOffset_D[15]), .B(branchOffset_regD[15]), .S0(n111), 
        .Y(n322) );
  MX2XL U281 ( .A(PCplus4_regI[0]), .B(PCplus4_regD[0]), .S0(n111), .Y(n323)
         );
  MX2XL U282 ( .A(PCplus4_regI[1]), .B(PCplus4_regD[1]), .S0(n111), .Y(n324)
         );
  MX2XL U283 ( .A(PCplus4_regI[2]), .B(PCplus4_regD[2]), .S0(n111), .Y(n325)
         );
  MX2XL U284 ( .A(PCplus4_regI[3]), .B(PCplus4_regD[3]), .S0(n111), .Y(n326)
         );
  MX2XL U285 ( .A(PCplus4_regI[4]), .B(PCplus4_regD[4]), .S0(n111), .Y(n327)
         );
  MX2XL U286 ( .A(PCplus4_regI[5]), .B(PCplus4_regD[5]), .S0(n111), .Y(n328)
         );
  MX2XL U287 ( .A(PCplus4_regI[6]), .B(PCplus4_regD[6]), .S0(n111), .Y(n329)
         );
  MX2XL U288 ( .A(PCplus4_regI[7]), .B(PCplus4_regD[7]), .S0(n111), .Y(n330)
         );
  MX2XL U289 ( .A(PCplus4_regI[8]), .B(PCplus4_regD[8]), .S0(n111), .Y(n331)
         );
  MX2XL U290 ( .A(PCplus4_regI[9]), .B(PCplus4_regD[9]), .S0(n128), .Y(n332)
         );
  MX2XL U291 ( .A(PCplus4_regI[11]), .B(PCplus4_regD[11]), .S0(n125), .Y(n334)
         );
  MX2XL U292 ( .A(PCplus4_regI[12]), .B(PCplus4_regD[12]), .S0(n125), .Y(n335)
         );
  MX2XL U293 ( .A(PCplus4_regI[13]), .B(PCplus4_regD[13]), .S0(n125), .Y(n336)
         );
  MX2XL U294 ( .A(PCplus4_regI[14]), .B(PCplus4_regD[14]), .S0(n125), .Y(n337)
         );
  MX2XL U295 ( .A(PCplus4_regI[15]), .B(PCplus4_regD[15]), .S0(n125), .Y(n338)
         );
  MX2XL U296 ( .A(PCplus4_regI[16]), .B(PCplus4_regD[16]), .S0(n125), .Y(n339)
         );
  MX2XL U297 ( .A(PCplus4_regI[17]), .B(PCplus4_regD[17]), .S0(n125), .Y(n340)
         );
  MX2XL U298 ( .A(PCplus4_regI[18]), .B(PCplus4_regD[18]), .S0(n125), .Y(n341)
         );
  MX2XL U299 ( .A(PCplus4_regI[19]), .B(PCplus4_regD[19]), .S0(n125), .Y(n342)
         );
  MX2XL U300 ( .A(PCplus4_regI[20]), .B(PCplus4_regD[20]), .S0(n125), .Y(n343)
         );
  MX2XL U301 ( .A(PCplus4_regI[21]), .B(PCplus4_regD[21]), .S0(n125), .Y(n344)
         );
  MX2XL U302 ( .A(PCplus4_regI[22]), .B(PCplus4_regD[22]), .S0(n128), .Y(n345)
         );
  MX2XL U303 ( .A(PCplus4_regI[23]), .B(PCplus4_regD[23]), .S0(n132), .Y(n346)
         );
  MX2XL U304 ( .A(PCplus4_regI[24]), .B(PCplus4_regD[24]), .S0(n132), .Y(n347)
         );
  MX2XL U305 ( .A(PCplus4_regI[25]), .B(PCplus4_regD[25]), .S0(n132), .Y(n348)
         );
  MX2XL U306 ( .A(PCplus4_regI[26]), .B(PCplus4_regD[26]), .S0(n132), .Y(n349)
         );
  MX2XL U307 ( .A(PCplus4_regI[27]), .B(PCplus4_regD[27]), .S0(n132), .Y(n350)
         );
  MX2XL U308 ( .A(PCplus4_regI[28]), .B(PCplus4_regD[28]), .S0(n132), .Y(n351)
         );
  MX2XL U309 ( .A(PCplus4_regI[29]), .B(PCplus4_regD[29]), .S0(n132), .Y(n352)
         );
  MX2XL U310 ( .A(PCplus4_regI[30]), .B(PCplus4_regD[30]), .S0(n132), .Y(n353)
         );
  MX2XL U311 ( .A(PCplus4_regI[31]), .B(PCplus4_regD[31]), .S0(n132), .Y(n354)
         );
  CLKINVX1 U312 ( .A(n124), .Y(n431) );
  CLKINVX1 U313 ( .A(n127), .Y(n432) );
  CLKINVX1 U314 ( .A(n105), .Y(n424) );
  CLKINVX1 U315 ( .A(n106), .Y(n425) );
  CLKINVX1 U316 ( .A(n107), .Y(n426) );
  CLKINVX1 U317 ( .A(n108), .Y(n427) );
  CLKINVX1 U318 ( .A(n109), .Y(n428) );
  CLKINVX1 U319 ( .A(n110), .Y(n433) );
  MX2XL U320 ( .A(RegWrite), .B(RegWrite_regD), .S0(n125), .Y(n290) );
  CLKBUFX2 U321 ( .A(stallcache), .Y(n13) );
endmodule


module EX_MEM_regFile ( clk, rst_n, stallcache, MemtoReg_regD, MemRead_regD, 
        MemWrite_regD, RegWrite_regD, B_regD, wsel_regD, ALUout, MemtoReg_regE, 
        MemRead_regE, MemWrite_regE, RegWrite_regE, B_regE, wsel_regE, 
        ALUout_regE );
  input [1:0] MemtoReg_regD;
  input [31:0] B_regD;
  input [4:0] wsel_regD;
  input [31:0] ALUout;
  output [1:0] MemtoReg_regE;
  output [31:0] B_regE;
  output [4:0] wsel_regE;
  output [31:0] ALUout_regE;
  input clk, rst_n, stallcache, MemRead_regD, MemWrite_regD, RegWrite_regD;
  output MemRead_regE, MemWrite_regE, RegWrite_regE;
  wire   n205, n206, n25, n30, n31, n32, n33, n35, n39, n41, n42, n45, n46,
         n48, n51, n54, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26,
         n27, n66, n68, n70, n146, n157, n160, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n182, n185, n187, n188, n191, n194, n195;

  DFFRX4 MemWrite_regE_reg ( .D(n104), .CK(clk), .RN(n175), .QN(n35) );
  DFFRX1 \ALUout_regE_reg[23]  ( .D(n136), .CK(clk), .RN(n178), .Q(
        ALUout_regE[23]) );
  DFFRX1 \ALUout_regE_reg[26]  ( .D(n139), .CK(clk), .RN(n178), .Q(
        ALUout_regE[26]) );
  DFFRX1 \MemtoReg_regE_reg[1]  ( .D(n107), .CK(clk), .RN(n176), .Q(
        MemtoReg_regE[1]) );
  DFFRX1 \MemtoReg_regE_reg[0]  ( .D(n106), .CK(clk), .RN(n175), .Q(
        MemtoReg_regE[0]) );
  DFFRHQX8 \ALUout_regE_reg[4]  ( .D(n117), .CK(clk), .RN(n176), .Q(
        ALUout_regE[4]) );
  DFFRX1 MemRead_regE_reg ( .D(n105), .CK(clk), .RN(n175), .Q(MemRead_regE) );
  DFFRX1 \ALUout_regE_reg[7]  ( .D(n120), .CK(clk), .RN(n177), .Q(
        ALUout_regE[7]), .QN(n46) );
  DFFRX4 \ALUout_regE_reg[28]  ( .D(n141), .CK(clk), .RN(n178), .Q(n205), .QN(
        n160) );
  DFFRX1 \ALUout_regE_reg[2]  ( .D(n115), .CK(clk), .RN(n176), .Q(n2), .QN(n41) );
  DFFRX2 \ALUout_regE_reg[24]  ( .D(n137), .CK(clk), .RN(n178), .Q(n206), .QN(
        n157) );
  DFFRX2 \ALUout_regE_reg[3]  ( .D(n116), .CK(clk), .RN(n176), .Q(
        ALUout_regE[3]), .QN(n42) );
  DFFRX4 \ALUout_regE_reg[6]  ( .D(n119), .CK(clk), .RN(n177), .QN(n45) );
  DFFRHQX8 \wsel_regE_reg[4]  ( .D(n112), .CK(clk), .RN(n176), .Q(wsel_regE[4]) );
  DFFRHQX8 \wsel_regE_reg[2]  ( .D(n110), .CK(clk), .RN(n176), .Q(wsel_regE[2]) );
  DFFRHQX8 \wsel_regE_reg[3]  ( .D(n111), .CK(clk), .RN(n176), .Q(wsel_regE[3]) );
  DFFRHQX8 \wsel_regE_reg[0]  ( .D(n108), .CK(clk), .RN(n176), .Q(wsel_regE[0]) );
  DFFRHQX8 \wsel_regE_reg[1]  ( .D(n109), .CK(clk), .RN(n176), .Q(wsel_regE[1]) );
  DFFRHQX8 RegWrite_regE_reg ( .D(n103), .CK(clk), .RN(n175), .Q(RegWrite_regE) );
  DFFRHQX8 \ALUout_regE_reg[10]  ( .D(n123), .CK(clk), .RN(rst_n), .Q(n188) );
  DFFSRX4 \ALUout_regE_reg[5]  ( .D(n118), .CK(clk), .SN(1'b1), .RN(rst_n), 
        .Q(ALUout_regE[5]) );
  DFFRX4 \ALUout_regE_reg[11]  ( .D(n124), .CK(clk), .RN(n177), .Q(
        ALUout_regE[11]) );
  DFFRX4 \ALUout_regE_reg[19]  ( .D(n132), .CK(clk), .RN(n178), .Q(
        ALUout_regE[19]) );
  DFFRX4 \ALUout_regE_reg[30]  ( .D(n143), .CK(clk), .RN(n179), .Q(
        ALUout_regE[30]) );
  DFFRX4 \ALUout_regE_reg[31]  ( .D(n144), .CK(clk), .RN(n179), .Q(
        ALUout_regE[31]) );
  DFFRX4 \ALUout_regE_reg[27]  ( .D(n140), .CK(clk), .RN(n178), .Q(
        ALUout_regE[27]) );
  DFFRX4 \ALUout_regE_reg[16]  ( .D(n129), .CK(clk), .RN(rst_n), .Q(
        ALUout_regE[16]) );
  DFFRX2 \ALUout_regE_reg[12]  ( .D(n125), .CK(clk), .RN(n177), .QN(n51) );
  DFFRX2 \ALUout_regE_reg[9]  ( .D(n122), .CK(clk), .RN(n177), .Q(
        ALUout_regE[9]), .QN(n48) );
  DFFRX2 \B_regE_reg[1]  ( .D(n72), .CK(clk), .RN(n173), .QN(n27) );
  DFFRX2 \B_regE_reg[0]  ( .D(n71), .CK(clk), .RN(n173), .QN(n26) );
  DFFRX2 \B_regE_reg[22]  ( .D(n93), .CK(clk), .RN(n174), .QN(n24) );
  DFFRX2 \B_regE_reg[20]  ( .D(n91), .CK(clk), .RN(n174), .QN(n23) );
  DFFRX2 \B_regE_reg[19]  ( .D(n90), .CK(clk), .RN(n174), .QN(n22) );
  DFFRX2 \B_regE_reg[24]  ( .D(n95), .CK(clk), .RN(n175), .QN(n21) );
  DFFRX2 \B_regE_reg[17]  ( .D(n88), .CK(clk), .RN(n174), .QN(n20) );
  DFFRX2 \B_regE_reg[18]  ( .D(n89), .CK(clk), .RN(n174), .QN(n19) );
  DFFRX2 \B_regE_reg[15]  ( .D(n86), .CK(clk), .RN(n174), .QN(n18) );
  DFFRX2 \B_regE_reg[16]  ( .D(n87), .CK(clk), .RN(n174), .QN(n17) );
  DFFRX2 \B_regE_reg[14]  ( .D(n85), .CK(clk), .RN(n174), .QN(n16) );
  DFFRX2 \B_regE_reg[25]  ( .D(n96), .CK(clk), .RN(n175), .QN(n15) );
  DFFRX2 \B_regE_reg[13]  ( .D(n84), .CK(clk), .RN(n174), .QN(n14) );
  DFFRX2 \B_regE_reg[10]  ( .D(n81), .CK(clk), .RN(n173), .QN(n13) );
  DFFRX2 \B_regE_reg[11]  ( .D(n82), .CK(clk), .RN(n173), .QN(n12) );
  DFFRX2 \B_regE_reg[12]  ( .D(n83), .CK(clk), .RN(n174), .QN(n11) );
  DFFRX2 \B_regE_reg[5]  ( .D(n76), .CK(clk), .RN(n173), .QN(n10) );
  DFFRX2 \B_regE_reg[3]  ( .D(n74), .CK(clk), .RN(n173), .QN(n9) );
  DFFRX2 \B_regE_reg[2]  ( .D(n73), .CK(clk), .RN(n173), .QN(n8) );
  DFFRX2 \B_regE_reg[7]  ( .D(n78), .CK(clk), .RN(n173), .QN(n7) );
  DFFRX2 \B_regE_reg[9]  ( .D(n80), .CK(clk), .RN(n173), .QN(n6) );
  DFFRX2 \B_regE_reg[8]  ( .D(n79), .CK(clk), .RN(n173), .QN(n5) );
  DFFRX2 \B_regE_reg[26]  ( .D(n97), .CK(clk), .RN(n175), .QN(n4) );
  DFFRX2 \B_regE_reg[27]  ( .D(n98), .CK(clk), .RN(n175), .QN(n3) );
  DFFRX2 \B_regE_reg[6]  ( .D(n77), .CK(clk), .RN(n173), .QN(n1) );
  DFFRX2 \B_regE_reg[31]  ( .D(n102), .CK(clk), .RN(n175), .QN(n33) );
  DFFRX2 \B_regE_reg[30]  ( .D(n101), .CK(clk), .RN(n175), .QN(n32) );
  DFFRX2 \B_regE_reg[29]  ( .D(n100), .CK(clk), .RN(n175), .QN(n31) );
  DFFRX2 \B_regE_reg[28]  ( .D(n99), .CK(clk), .RN(n175), .QN(n30) );
  DFFRX2 \B_regE_reg[23]  ( .D(n94), .CK(clk), .RN(n174), .QN(n25) );
  DFFSRHQX2 \B_regE_reg[4]  ( .D(n75), .CK(clk), .SN(1'b1), .RN(rst_n), .Q(
        n194) );
  DFFSRHQX2 \B_regE_reg[21]  ( .D(n92), .CK(clk), .SN(1'b1), .RN(rst_n), .Q(
        n195) );
  DFFRHQX4 \ALUout_regE_reg[13]  ( .D(n126), .CK(clk), .RN(rst_n), .Q(n191) );
  DFFRX4 \ALUout_regE_reg[29]  ( .D(n142), .CK(clk), .RN(n178), .Q(
        ALUout_regE[29]) );
  DFFRX4 \ALUout_regE_reg[8]  ( .D(n121), .CK(clk), .RN(n177), .Q(
        ALUout_regE[8]) );
  DFFRX4 \ALUout_regE_reg[25]  ( .D(n138), .CK(clk), .RN(n178), .Q(
        ALUout_regE[25]) );
  DFFRX4 \ALUout_regE_reg[18]  ( .D(n131), .CK(clk), .RN(n178), .Q(
        ALUout_regE[18]) );
  DFFRX4 \ALUout_regE_reg[20]  ( .D(n133), .CK(clk), .RN(n178), .Q(
        ALUout_regE[20]) );
  DFFRX4 \ALUout_regE_reg[14]  ( .D(n127), .CK(clk), .RN(n177), .Q(
        ALUout_regE[14]) );
  DFFRX4 \ALUout_regE_reg[17]  ( .D(n130), .CK(clk), .RN(n177), .Q(
        ALUout_regE[17]) );
  DFFRX4 \ALUout_regE_reg[15]  ( .D(n128), .CK(clk), .RN(n177), .QN(n54) );
  DFFRX4 \ALUout_regE_reg[0]  ( .D(n113), .CK(clk), .RN(n176), .QN(n39) );
  DFFRX4 \ALUout_regE_reg[21]  ( .D(n134), .CK(clk), .RN(n178), .Q(
        ALUout_regE[21]) );
  DFFRX4 \ALUout_regE_reg[22]  ( .D(n135), .CK(clk), .RN(n178), .Q(
        ALUout_regE[22]) );
  DFFRX4 \ALUout_regE_reg[1]  ( .D(n114), .CK(clk), .RN(n176), .Q(
        ALUout_regE[1]) );
  MX2X2 U2 ( .A(ALUout[28]), .B(n205), .S0(n166), .Y(n141) );
  MX2X2 U3 ( .A(ALUout[30]), .B(ALUout_regE[30]), .S0(n166), .Y(n143) );
  MX2X2 U4 ( .A(ALUout[17]), .B(ALUout_regE[17]), .S0(n165), .Y(n130) );
  MX2X2 U5 ( .A(ALUout[3]), .B(n182), .S0(n164), .Y(n116) );
  MX2X1 U6 ( .A(ALUout[22]), .B(ALUout_regE[22]), .S0(n165), .Y(n135) );
  INVX6 U7 ( .A(n39), .Y(ALUout_regE[0]) );
  CLKMX2X3 U8 ( .A(ALUout[19]), .B(ALUout_regE[19]), .S0(n165), .Y(n132) );
  INVX6 U9 ( .A(n45), .Y(ALUout_regE[6]) );
  MX2X1 U10 ( .A(ALUout[21]), .B(ALUout_regE[21]), .S0(n165), .Y(n134) );
  CLKINVX8 U11 ( .A(n54), .Y(ALUout_regE[15]) );
  MX2X1 U12 ( .A(ALUout[15]), .B(ALUout_regE[15]), .S0(n165), .Y(n128) );
  CLKMX2X2 U13 ( .A(ALUout[13]), .B(ALUout_regE[13]), .S0(n165), .Y(n126) );
  MX2X1 U14 ( .A(ALUout[14]), .B(ALUout_regE[14]), .S0(n165), .Y(n127) );
  MX2X1 U15 ( .A(ALUout[20]), .B(ALUout_regE[20]), .S0(n165), .Y(n133) );
  MX2X1 U16 ( .A(ALUout[18]), .B(ALUout_regE[18]), .S0(n165), .Y(n131) );
  MX2X2 U17 ( .A(ALUout[25]), .B(ALUout_regE[25]), .S0(n165), .Y(n138) );
  MX2X1 U18 ( .A(ALUout[8]), .B(ALUout_regE[8]), .S0(n164), .Y(n121) );
  MX2X1 U19 ( .A(ALUout[29]), .B(ALUout_regE[29]), .S0(n166), .Y(n142) );
  INVX16 U20 ( .A(n26), .Y(B_regE[0]) );
  INVX16 U21 ( .A(n27), .Y(B_regE[1]) );
  INVX16 U22 ( .A(n8), .Y(B_regE[2]) );
  INVX16 U23 ( .A(n9), .Y(B_regE[3]) );
  INVX16 U24 ( .A(n68), .Y(B_regE[4]) );
  CLKINVX1 U25 ( .A(n194), .Y(n68) );
  INVX16 U26 ( .A(n10), .Y(B_regE[5]) );
  INVX16 U27 ( .A(n1), .Y(B_regE[6]) );
  INVX16 U28 ( .A(n7), .Y(B_regE[7]) );
  INVX16 U29 ( .A(n5), .Y(B_regE[8]) );
  INVX16 U30 ( .A(n6), .Y(B_regE[9]) );
  INVX16 U31 ( .A(n13), .Y(B_regE[10]) );
  INVX16 U32 ( .A(n12), .Y(B_regE[11]) );
  INVX16 U33 ( .A(n11), .Y(B_regE[12]) );
  INVX16 U34 ( .A(n14), .Y(B_regE[13]) );
  INVX16 U35 ( .A(n16), .Y(B_regE[14]) );
  INVX16 U36 ( .A(n18), .Y(B_regE[15]) );
  INVX16 U37 ( .A(n17), .Y(B_regE[16]) );
  INVX16 U38 ( .A(n20), .Y(B_regE[17]) );
  INVX16 U39 ( .A(n19), .Y(B_regE[18]) );
  INVX16 U40 ( .A(n22), .Y(B_regE[19]) );
  INVX16 U41 ( .A(n23), .Y(B_regE[20]) );
  INVX16 U42 ( .A(n66), .Y(B_regE[21]) );
  CLKINVX1 U43 ( .A(n195), .Y(n66) );
  INVX16 U44 ( .A(n24), .Y(B_regE[22]) );
  INVX16 U45 ( .A(n25), .Y(B_regE[23]) );
  INVX16 U46 ( .A(n21), .Y(B_regE[24]) );
  INVX16 U47 ( .A(n15), .Y(B_regE[25]) );
  INVX16 U48 ( .A(n4), .Y(B_regE[26]) );
  INVX16 U49 ( .A(n3), .Y(B_regE[27]) );
  INVX16 U50 ( .A(n30), .Y(B_regE[28]) );
  INVX16 U51 ( .A(n31), .Y(B_regE[29]) );
  INVX16 U52 ( .A(n32), .Y(B_regE[30]) );
  INVX16 U53 ( .A(n33), .Y(B_regE[31]) );
  INVX16 U54 ( .A(n41), .Y(ALUout_regE[2]) );
  CLKMX2X4 U55 ( .A(ALUout[31]), .B(ALUout_regE[31]), .S0(n166), .Y(n144) );
  MX2X1 U56 ( .A(ALUout[5]), .B(ALUout_regE[5]), .S0(n164), .Y(n118) );
  CLKMX2X2 U57 ( .A(B_regD[27]), .B(B_regE[27]), .S0(n168), .Y(n98) );
  MX2X4 U58 ( .A(ALUout[10]), .B(ALUout_regE[10]), .S0(n164), .Y(n123) );
  INVX4 U59 ( .A(n51), .Y(ALUout_regE[12]) );
  CLKMX2X4 U60 ( .A(ALUout[9]), .B(n187), .S0(n164), .Y(n122) );
  MX2X2 U61 ( .A(ALUout[12]), .B(ALUout_regE[12]), .S0(n164), .Y(n125) );
  CLKMX2X2 U62 ( .A(B_regD[26]), .B(B_regE[26]), .S0(n168), .Y(n97) );
  MX2X1 U63 ( .A(ALUout[16]), .B(ALUout_regE[16]), .S0(n165), .Y(n129) );
  CLKMX2X3 U64 ( .A(ALUout[27]), .B(ALUout_regE[27]), .S0(n166), .Y(n140) );
  CLKMX2X4 U65 ( .A(ALUout[11]), .B(ALUout_regE[11]), .S0(n164), .Y(n124) );
  MX2X1 U66 ( .A(B_regD[29]), .B(B_regE[29]), .S0(n169), .Y(n100) );
  INVX12 U67 ( .A(n188), .Y(n70) );
  CLKINVX20 U68 ( .A(n70), .Y(ALUout_regE[10]) );
  INVX12 U69 ( .A(n191), .Y(n146) );
  CLKINVX20 U70 ( .A(n146), .Y(ALUout_regE[13]) );
  CLKMX2X2 U74 ( .A(B_regD[23]), .B(B_regE[23]), .S0(n168), .Y(n94) );
  MX2X1 U75 ( .A(B_regD[21]), .B(B_regE[21]), .S0(n168), .Y(n92) );
  MX2XL U76 ( .A(B_regD[30]), .B(B_regE[30]), .S0(n169), .Y(n101) );
  MX2XL U77 ( .A(wsel_regD[4]), .B(wsel_regE[4]), .S0(n166), .Y(n112) );
  MX2X1 U78 ( .A(wsel_regD[0]), .B(wsel_regE[0]), .S0(n166), .Y(n108) );
  CLKMX2X2 U79 ( .A(B_regD[4]), .B(B_regE[4]), .S0(n167), .Y(n75) );
  CLKMX2X2 U80 ( .A(ALUout[23]), .B(ALUout_regE[23]), .S0(n165), .Y(n136) );
  MX2X1 U81 ( .A(ALUout[4]), .B(ALUout_regE[4]), .S0(n164), .Y(n117) );
  MX2X2 U82 ( .A(ALUout[7]), .B(n185), .S0(n164), .Y(n120) );
  CLKMX2X2 U83 ( .A(ALUout[24]), .B(n206), .S0(n165), .Y(n137) );
  CLKMX2X2 U84 ( .A(ALUout[0]), .B(ALUout_regE[0]), .S0(n164), .Y(n113) );
  MX2X2 U85 ( .A(ALUout[6]), .B(ALUout_regE[6]), .S0(n164), .Y(n119) );
  CLKMX2X2 U86 ( .A(ALUout[1]), .B(ALUout_regE[1]), .S0(n164), .Y(n114) );
  CLKMX2X2 U87 ( .A(ALUout[2]), .B(n2), .S0(n164), .Y(n115) );
  MX2XL U88 ( .A(B_regD[8]), .B(B_regE[8]), .S0(n167), .Y(n79) );
  MX2XL U89 ( .A(B_regD[9]), .B(B_regE[9]), .S0(n167), .Y(n80) );
  MX2XL U90 ( .A(B_regD[6]), .B(B_regE[6]), .S0(n167), .Y(n77) );
  MX2XL U91 ( .A(B_regD[7]), .B(B_regE[7]), .S0(n167), .Y(n78) );
  MX2XL U92 ( .A(B_regD[2]), .B(B_regE[2]), .S0(n167), .Y(n73) );
  MX2XL U93 ( .A(B_regD[3]), .B(B_regE[3]), .S0(n167), .Y(n74) );
  MX2XL U94 ( .A(B_regD[5]), .B(B_regE[5]), .S0(n167), .Y(n76) );
  MX2XL U95 ( .A(B_regD[12]), .B(B_regE[12]), .S0(n167), .Y(n83) );
  MX2XL U96 ( .A(B_regD[11]), .B(B_regE[11]), .S0(n167), .Y(n82) );
  MX2XL U97 ( .A(B_regD[10]), .B(B_regE[10]), .S0(n167), .Y(n81) );
  MX2XL U98 ( .A(B_regD[13]), .B(B_regE[13]), .S0(n167), .Y(n84) );
  MX2XL U99 ( .A(B_regD[25]), .B(B_regE[25]), .S0(n168), .Y(n96) );
  MX2XL U100 ( .A(B_regD[14]), .B(B_regE[14]), .S0(n167), .Y(n85) );
  MX2XL U101 ( .A(B_regD[16]), .B(B_regE[16]), .S0(n168), .Y(n87) );
  MX2XL U102 ( .A(B_regD[15]), .B(B_regE[15]), .S0(n168), .Y(n86) );
  MX2XL U103 ( .A(B_regD[18]), .B(B_regE[18]), .S0(n168), .Y(n89) );
  MX2XL U104 ( .A(B_regD[17]), .B(B_regE[17]), .S0(n168), .Y(n88) );
  MX2XL U105 ( .A(B_regD[24]), .B(B_regE[24]), .S0(n168), .Y(n95) );
  MX2XL U106 ( .A(B_regD[19]), .B(B_regE[19]), .S0(n168), .Y(n90) );
  MX2XL U107 ( .A(B_regD[20]), .B(B_regE[20]), .S0(n168), .Y(n91) );
  MX2XL U108 ( .A(B_regD[22]), .B(B_regE[22]), .S0(n168), .Y(n93) );
  INVX20 U109 ( .A(n35), .Y(MemWrite_regE) );
  INVX20 U110 ( .A(n157), .Y(ALUout_regE[24]) );
  BUFX8 U111 ( .A(n163), .Y(n171) );
  CLKBUFX2 U112 ( .A(n163), .Y(n170) );
  MX2XL U113 ( .A(wsel_regD[3]), .B(wsel_regE[3]), .S0(n166), .Y(n111) );
  CLKMX2X2 U114 ( .A(ALUout[26]), .B(ALUout_regE[26]), .S0(n166), .Y(n139) );
  CLKBUFX2 U115 ( .A(rst_n), .Y(n172) );
  MX2XL U116 ( .A(B_regD[0]), .B(B_regE[0]), .S0(n166), .Y(n71) );
  MX2XL U117 ( .A(B_regD[1]), .B(B_regE[1]), .S0(n166), .Y(n72) );
  MX2XL U118 ( .A(B_regD[31]), .B(B_regE[31]), .S0(n169), .Y(n102) );
  MX2XL U119 ( .A(MemWrite_regD), .B(MemWrite_regE), .S0(n169), .Y(n104) );
  MX2XL U120 ( .A(wsel_regD[1]), .B(wsel_regE[1]), .S0(n166), .Y(n109) );
  INVX20 U121 ( .A(n160), .Y(ALUout_regE[28]) );
  CLKBUFX3 U122 ( .A(n170), .Y(n166) );
  CLKBUFX3 U123 ( .A(n171), .Y(n165) );
  CLKBUFX3 U124 ( .A(n171), .Y(n164) );
  CLKBUFX3 U125 ( .A(n170), .Y(n167) );
  CLKBUFX3 U126 ( .A(n171), .Y(n168) );
  CLKBUFX3 U127 ( .A(n171), .Y(n169) );
  CLKBUFX3 U128 ( .A(n172), .Y(n174) );
  CLKBUFX3 U129 ( .A(n172), .Y(n175) );
  CLKBUFX3 U130 ( .A(n172), .Y(n176) );
  CLKBUFX3 U131 ( .A(n179), .Y(n177) );
  CLKBUFX3 U132 ( .A(n172), .Y(n178) );
  CLKBUFX3 U133 ( .A(n172), .Y(n179) );
  CLKBUFX3 U134 ( .A(n179), .Y(n173) );
  MX2XL U135 ( .A(wsel_regD[2]), .B(wsel_regE[2]), .S0(n166), .Y(n110) );
  MX2XL U136 ( .A(B_regD[28]), .B(B_regE[28]), .S0(n169), .Y(n99) );
  MX2XL U137 ( .A(RegWrite_regD), .B(RegWrite_regE), .S0(n169), .Y(n103) );
  MX2XL U138 ( .A(MemRead_regD), .B(MemRead_regE), .S0(n169), .Y(n105) );
  MX2XL U139 ( .A(MemtoReg_regD[0]), .B(MemtoReg_regE[0]), .S0(n169), .Y(n106)
         );
  MX2XL U140 ( .A(MemtoReg_regD[1]), .B(MemtoReg_regE[1]), .S0(n169), .Y(n107)
         );
  CLKINVX1 U141 ( .A(n42), .Y(n182) );
  CLKINVX1 U142 ( .A(n46), .Y(n185) );
  CLKINVX1 U143 ( .A(n48), .Y(n187) );
  CLKBUFX2 U144 ( .A(stallcache), .Y(n163) );
endmodule


module MEM_WB_regFile ( clk, rst_n, stallcache, MemtoReg_regE, RegWrite_regE, 
        ALUout_regE, wsel_regE, dataOut, MemtoReg_regM, RegWrite_regM, 
        ALUout_regM, wsel_regM, dataOut_regM );
  input [1:0] MemtoReg_regE;
  input [31:0] ALUout_regE;
  input [4:0] wsel_regE;
  input [31:0] dataOut;
  output [1:0] MemtoReg_regM;
  output [31:0] ALUout_regM;
  output [4:0] wsel_regM;
  output [31:0] dataOut_regM;
  input clk, rst_n, stallcache, RegWrite_regE;
  output RegWrite_regM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224;

  DFFRX4 \dataOut_regM_reg[28]  ( .D(n137), .CK(clk), .RN(n158), .Q(
        dataOut_regM[28]), .QN(n65) );
  DFFRX4 \dataOut_regM_reg[7]  ( .D(n116), .CK(clk), .RN(n156), .Q(
        dataOut_regM[7]), .QN(n44) );
  DFFRX1 \dataOut_regM_reg[16]  ( .D(n125), .CK(clk), .RN(n157), .Q(
        dataOut_regM[16]), .QN(n53) );
  DFFRX1 \dataOut_regM_reg[20]  ( .D(n129), .CK(clk), .RN(n158), .Q(
        dataOut_regM[20]), .QN(n57) );
  DFFRX1 \dataOut_regM_reg[13]  ( .D(n122), .CK(clk), .RN(n157), .Q(
        dataOut_regM[13]), .QN(n50) );
  DFFRX1 \dataOut_regM_reg[12]  ( .D(n121), .CK(clk), .RN(n157), .Q(
        dataOut_regM[12]), .QN(n49) );
  DFFRX1 \dataOut_regM_reg[17]  ( .D(n126), .CK(clk), .RN(n157), .Q(
        dataOut_regM[17]), .QN(n54) );
  DFFRX1 \dataOut_regM_reg[8]  ( .D(n117), .CK(clk), .RN(n157), .Q(
        dataOut_regM[8]), .QN(n45) );
  DFFRX1 \dataOut_regM_reg[22]  ( .D(n131), .CK(clk), .RN(n158), .Q(
        dataOut_regM[22]), .QN(n59) );
  DFFRX1 \dataOut_regM_reg[15]  ( .D(n124), .CK(clk), .RN(n157), .Q(
        dataOut_regM[15]), .QN(n52) );
  DFFRX1 \dataOut_regM_reg[10]  ( .D(n119), .CK(clk), .RN(n157), .Q(
        dataOut_regM[10]), .QN(n47) );
  DFFRX1 \dataOut_regM_reg[14]  ( .D(n123), .CK(clk), .RN(n157), .Q(
        dataOut_regM[14]), .QN(n51) );
  DFFRX1 \dataOut_regM_reg[11]  ( .D(n120), .CK(clk), .RN(n157), .Q(
        dataOut_regM[11]), .QN(n48) );
  DFFRX1 \dataOut_regM_reg[21]  ( .D(n130), .CK(clk), .RN(n158), .Q(
        dataOut_regM[21]), .QN(n58) );
  DFFRX1 \dataOut_regM_reg[23]  ( .D(n132), .CK(clk), .RN(n158), .Q(
        dataOut_regM[23]), .QN(n60) );
  DFFRX1 \dataOut_regM_reg[9]  ( .D(n118), .CK(clk), .RN(n157), .Q(
        dataOut_regM[9]), .QN(n46) );
  DFFRX1 \dataOut_regM_reg[18]  ( .D(n127), .CK(clk), .RN(n157), .Q(
        dataOut_regM[18]), .QN(n55) );
  DFFRX1 \dataOut_regM_reg[19]  ( .D(n128), .CK(clk), .RN(n157), .Q(
        dataOut_regM[19]), .QN(n56) );
  DFFRX1 \dataOut_regM_reg[6]  ( .D(n115), .CK(clk), .RN(n156), .Q(
        dataOut_regM[6]), .QN(n43) );
  DFFRX1 \dataOut_regM_reg[5]  ( .D(n114), .CK(clk), .RN(n156), .Q(
        dataOut_regM[5]), .QN(n42) );
  DFFRX1 \dataOut_regM_reg[4]  ( .D(n113), .CK(clk), .RN(n156), .Q(
        dataOut_regM[4]), .QN(n41) );
  DFFRX1 \dataOut_regM_reg[0]  ( .D(n109), .CK(clk), .RN(n156), .Q(
        dataOut_regM[0]), .QN(n37) );
  DFFRX1 \dataOut_regM_reg[1]  ( .D(n110), .CK(clk), .RN(n156), .Q(
        dataOut_regM[1]), .QN(n38) );
  DFFRX1 \ALUout_regM_reg[16]  ( .D(n85), .CK(clk), .RN(n154), .Q(
        ALUout_regM[16]), .QN(n18) );
  DFFRX1 \ALUout_regM_reg[20]  ( .D(n89), .CK(clk), .RN(n154), .Q(
        ALUout_regM[20]), .QN(n22) );
  DFFRX1 \ALUout_regM_reg[13]  ( .D(n82), .CK(clk), .RN(n154), .Q(
        ALUout_regM[13]), .QN(n15) );
  DFFRX1 \ALUout_regM_reg[12]  ( .D(n81), .CK(clk), .RN(n154), .Q(
        ALUout_regM[12]), .QN(n14) );
  DFFRX1 \ALUout_regM_reg[17]  ( .D(n86), .CK(clk), .RN(n154), .Q(
        ALUout_regM[17]), .QN(n19) );
  DFFRX1 \ALUout_regM_reg[8]  ( .D(n77), .CK(clk), .RN(n153), .Q(
        ALUout_regM[8]), .QN(n10) );
  DFFRX1 \ALUout_regM_reg[22]  ( .D(n91), .CK(clk), .RN(n154), .Q(
        ALUout_regM[22]), .QN(n24) );
  DFFRX1 \ALUout_regM_reg[15]  ( .D(n84), .CK(clk), .RN(n154), .Q(
        ALUout_regM[15]), .QN(n17) );
  DFFRX1 \ALUout_regM_reg[10]  ( .D(n79), .CK(clk), .RN(n153), .Q(
        ALUout_regM[10]), .QN(n12) );
  DFFRX1 \ALUout_regM_reg[14]  ( .D(n83), .CK(clk), .RN(n154), .Q(
        ALUout_regM[14]), .QN(n16) );
  DFFRX1 \ALUout_regM_reg[11]  ( .D(n80), .CK(clk), .RN(n153), .Q(
        ALUout_regM[11]), .QN(n13) );
  DFFRX1 \ALUout_regM_reg[21]  ( .D(n90), .CK(clk), .RN(n154), .Q(
        ALUout_regM[21]), .QN(n23) );
  DFFRX1 \ALUout_regM_reg[23]  ( .D(n92), .CK(clk), .RN(n154), .Q(
        ALUout_regM[23]), .QN(n25) );
  DFFRX1 \ALUout_regM_reg[9]  ( .D(n78), .CK(clk), .RN(n153), .Q(
        ALUout_regM[9]), .QN(n11) );
  DFFRX1 \ALUout_regM_reg[18]  ( .D(n87), .CK(clk), .RN(n154), .Q(
        ALUout_regM[18]), .QN(n20) );
  DFFRX1 \ALUout_regM_reg[19]  ( .D(n88), .CK(clk), .RN(n154), .Q(
        ALUout_regM[19]), .QN(n21) );
  DFFRX1 \ALUout_regM_reg[6]  ( .D(n75), .CK(clk), .RN(n153), .Q(
        ALUout_regM[6]), .QN(n8) );
  DFFRX1 \ALUout_regM_reg[5]  ( .D(n74), .CK(clk), .RN(n153), .Q(
        ALUout_regM[5]), .QN(n7) );
  DFFRX1 \ALUout_regM_reg[26]  ( .D(n95), .CK(clk), .RN(n155), .Q(
        ALUout_regM[26]), .QN(n28) );
  DFFRX1 \ALUout_regM_reg[4]  ( .D(n73), .CK(clk), .RN(n153), .Q(
        ALUout_regM[4]), .QN(n6) );
  DFFRX1 \ALUout_regM_reg[25]  ( .D(n94), .CK(clk), .RN(n155), .Q(
        ALUout_regM[25]), .QN(n27) );
  DFFRX1 \dataOut_regM_reg[3]  ( .D(n112), .CK(clk), .RN(n156), .Q(
        dataOut_regM[3]), .QN(n40) );
  DFFRX1 \dataOut_regM_reg[2]  ( .D(n111), .CK(clk), .RN(n156), .Q(
        dataOut_regM[2]), .QN(n39) );
  DFFRX1 \ALUout_regM_reg[31]  ( .D(n100), .CK(clk), .RN(n155), .Q(
        ALUout_regM[31]), .QN(n33) );
  DFFRX1 \ALUout_regM_reg[30]  ( .D(n99), .CK(clk), .RN(n155), .Q(
        ALUout_regM[30]), .QN(n32) );
  DFFRX1 \ALUout_regM_reg[29]  ( .D(n98), .CK(clk), .RN(n155), .Q(
        ALUout_regM[29]), .QN(n31) );
  DFFRX1 \ALUout_regM_reg[3]  ( .D(n72), .CK(clk), .RN(n153), .Q(
        ALUout_regM[3]), .QN(n5) );
  DFFRX1 \ALUout_regM_reg[1]  ( .D(n70), .CK(clk), .RN(n153), .Q(
        ALUout_regM[1]), .QN(n3) );
  DFFRX1 \ALUout_regM_reg[0]  ( .D(n69), .CK(clk), .RN(n153), .Q(
        ALUout_regM[0]), .QN(n2) );
  DFFRX1 \dataOut_regM_reg[27]  ( .D(n136), .CK(clk), .RN(n158), .Q(
        dataOut_regM[27]), .QN(n64) );
  DFFRX1 \dataOut_regM_reg[24]  ( .D(n133), .CK(clk), .RN(n158), .Q(
        dataOut_regM[24]), .QN(n61) );
  DFFRX1 \ALUout_regM_reg[28]  ( .D(n97), .CK(clk), .RN(n155), .Q(
        ALUout_regM[28]), .QN(n30) );
  DFFRX1 \ALUout_regM_reg[27]  ( .D(n96), .CK(clk), .RN(n155), .Q(
        ALUout_regM[27]), .QN(n29) );
  DFFRX1 \ALUout_regM_reg[24]  ( .D(n93), .CK(clk), .RN(n155), .Q(
        ALUout_regM[24]), .QN(n26) );
  DFFRX1 \ALUout_regM_reg[7]  ( .D(n76), .CK(clk), .RN(n153), .Q(
        ALUout_regM[7]), .QN(n9) );
  DFFRX1 \ALUout_regM_reg[2]  ( .D(n71), .CK(clk), .RN(n153), .Q(
        ALUout_regM[2]), .QN(n4) );
  DFFRX4 \MemtoReg_regM_reg[0]  ( .D(n102), .CK(clk), .RN(n155), .Q(
        MemtoReg_regM[0]), .QN(n35) );
  DFFRX4 RegWrite_regM_reg ( .D(n101), .CK(clk), .RN(n155), .Q(RegWrite_regM), 
        .QN(n34) );
  DFFRHQX8 \wsel_regM_reg[0]  ( .D(n104), .CK(clk), .RN(n155), .Q(wsel_regM[0]) );
  DFFRHQX8 \wsel_regM_reg[3]  ( .D(n107), .CK(clk), .RN(n156), .Q(wsel_regM[3]) );
  DFFRHQX8 \wsel_regM_reg[4]  ( .D(n108), .CK(clk), .RN(n156), .Q(wsel_regM[4]) );
  DFFRHQX8 \wsel_regM_reg[1]  ( .D(n105), .CK(clk), .RN(n156), .Q(wsel_regM[1]) );
  DFFRHQX8 \wsel_regM_reg[2]  ( .D(n106), .CK(clk), .RN(n156), .Q(wsel_regM[2]) );
  DFFSRHQX4 \MemtoReg_regM_reg[1]  ( .D(n103), .CK(clk), .SN(1'b1), .RN(rst_n), 
        .Q(MemtoReg_regM[1]) );
  DFFRX2 \dataOut_regM_reg[25]  ( .D(n134), .CK(clk), .RN(n158), .Q(
        dataOut_regM[25]), .QN(n62) );
  DFFRX2 \dataOut_regM_reg[30]  ( .D(n139), .CK(clk), .RN(n158), .Q(
        dataOut_regM[30]), .QN(n67) );
  DFFRX2 \dataOut_regM_reg[31]  ( .D(n140), .CK(clk), .RN(n158), .Q(
        dataOut_regM[31]), .QN(n68) );
  DFFRX2 \dataOut_regM_reg[29]  ( .D(n138), .CK(clk), .RN(n158), .Q(
        dataOut_regM[29]), .QN(n66) );
  DFFRX2 \dataOut_regM_reg[26]  ( .D(n135), .CK(clk), .RN(n158), .Q(
        dataOut_regM[26]), .QN(n63) );
  MX2X1 U2 ( .A(dataOut[26]), .B(n185), .S0(n150), .Y(n135) );
  MX2X1 U3 ( .A(dataOut[25]), .B(n184), .S0(n147), .Y(n134) );
  CLKMX2X2 U4 ( .A(MemtoReg_regE[0]), .B(n224), .S0(n148), .Y(n102) );
  CLKMX2X2 U5 ( .A(dataOut[4]), .B(n163), .S0(n146), .Y(n113) );
  CLKBUFX3 U6 ( .A(n145), .Y(n150) );
  CLKBUFX3 U7 ( .A(n145), .Y(n149) );
  BUFX2 U8 ( .A(n145), .Y(n151) );
  CLKMX2X2 U9 ( .A(dataOut[24]), .B(n183), .S0(n147), .Y(n133) );
  MX2X2 U10 ( .A(dataOut[29]), .B(n188), .S0(stallcache), .Y(n138) );
  MX2X2 U11 ( .A(dataOut[31]), .B(n190), .S0(stallcache), .Y(n140) );
  MX2X2 U12 ( .A(dataOut[30]), .B(n189), .S0(stallcache), .Y(n139) );
  MX2XL U14 ( .A(wsel_regE[4]), .B(wsel_regM[4]), .S0(n150), .Y(n108) );
  MX2XL U15 ( .A(wsel_regE[0]), .B(wsel_regM[0]), .S0(n150), .Y(n104) );
  MX2XL U16 ( .A(wsel_regE[3]), .B(wsel_regM[3]), .S0(n150), .Y(n107) );
  CLKBUFX2 U17 ( .A(rst_n), .Y(n152) );
  MX2X1 U18 ( .A(dataOut[8]), .B(n167), .S0(n146), .Y(n117) );
  MX2X1 U19 ( .A(dataOut[9]), .B(n168), .S0(n146), .Y(n118) );
  MX2X1 U20 ( .A(dataOut[1]), .B(n160), .S0(n146), .Y(n110) );
  MX2X1 U21 ( .A(dataOut[2]), .B(n161), .S0(n146), .Y(n111) );
  MX2X1 U22 ( .A(dataOut[3]), .B(n162), .S0(n146), .Y(n112) );
  MX2X1 U23 ( .A(dataOut[5]), .B(n164), .S0(n146), .Y(n114) );
  MX2X1 U24 ( .A(dataOut[6]), .B(n165), .S0(n146), .Y(n115) );
  MX2X1 U25 ( .A(dataOut[10]), .B(n169), .S0(n146), .Y(n119) );
  MX2X1 U26 ( .A(dataOut[11]), .B(n170), .S0(n146), .Y(n120) );
  MX2X1 U27 ( .A(dataOut[12]), .B(n171), .S0(n146), .Y(n121) );
  MX2X1 U28 ( .A(dataOut[14]), .B(n173), .S0(n147), .Y(n123) );
  MX2X1 U29 ( .A(dataOut[15]), .B(n174), .S0(n147), .Y(n124) );
  MX2X1 U30 ( .A(dataOut[16]), .B(n175), .S0(n147), .Y(n125) );
  MX2X1 U31 ( .A(dataOut[17]), .B(n176), .S0(n147), .Y(n126) );
  MX2X1 U32 ( .A(dataOut[18]), .B(n177), .S0(n147), .Y(n127) );
  MX2X1 U33 ( .A(dataOut[19]), .B(n178), .S0(n147), .Y(n128) );
  MX2X1 U34 ( .A(dataOut[20]), .B(n179), .S0(n147), .Y(n129) );
  MX2X1 U35 ( .A(dataOut[21]), .B(n180), .S0(n147), .Y(n130) );
  MX2X1 U36 ( .A(dataOut[22]), .B(n181), .S0(n147), .Y(n131) );
  MX2X1 U37 ( .A(dataOut[23]), .B(n182), .S0(n147), .Y(n132) );
  MX2X1 U38 ( .A(dataOut[0]), .B(n159), .S0(n146), .Y(n109) );
  MX2X1 U39 ( .A(dataOut[13]), .B(n172), .S0(n147), .Y(n122) );
  MX2XL U40 ( .A(wsel_regE[1]), .B(wsel_regM[1]), .S0(n150), .Y(n105) );
  CLKBUFX3 U41 ( .A(n151), .Y(n146) );
  CLKBUFX3 U42 ( .A(n151), .Y(n147) );
  CLKBUFX3 U43 ( .A(n149), .Y(n148) );
  CLKBUFX3 U44 ( .A(n152), .Y(n153) );
  CLKBUFX3 U45 ( .A(n152), .Y(n154) );
  CLKBUFX3 U46 ( .A(n152), .Y(n155) );
  CLKBUFX3 U47 ( .A(n152), .Y(n156) );
  CLKBUFX3 U48 ( .A(n152), .Y(n157) );
  CLKBUFX3 U49 ( .A(n152), .Y(n158) );
  CLKINVX1 U50 ( .A(n37), .Y(n159) );
  CLKINVX1 U51 ( .A(n38), .Y(n160) );
  CLKINVX1 U52 ( .A(n39), .Y(n161) );
  CLKINVX1 U53 ( .A(n40), .Y(n162) );
  CLKINVX1 U54 ( .A(n41), .Y(n163) );
  CLKINVX1 U55 ( .A(n42), .Y(n164) );
  CLKINVX1 U56 ( .A(n43), .Y(n165) );
  CLKMX2X2 U57 ( .A(dataOut[7]), .B(n166), .S0(n146), .Y(n116) );
  INVX1 U58 ( .A(n44), .Y(n166) );
  CLKINVX1 U59 ( .A(n47), .Y(n169) );
  CLKINVX1 U60 ( .A(n48), .Y(n170) );
  CLKINVX1 U61 ( .A(n49), .Y(n171) );
  CLKINVX1 U62 ( .A(n50), .Y(n172) );
  CLKINVX1 U63 ( .A(n51), .Y(n173) );
  CLKINVX1 U64 ( .A(n52), .Y(n174) );
  CLKINVX1 U65 ( .A(n53), .Y(n175) );
  CLKINVX1 U66 ( .A(n54), .Y(n176) );
  CLKINVX1 U67 ( .A(n55), .Y(n177) );
  CLKINVX1 U68 ( .A(n56), .Y(n178) );
  CLKINVX1 U69 ( .A(n57), .Y(n179) );
  CLKINVX1 U70 ( .A(n58), .Y(n180) );
  CLKINVX1 U71 ( .A(n59), .Y(n181) );
  CLKINVX1 U72 ( .A(n60), .Y(n182) );
  CLKINVX1 U73 ( .A(n61), .Y(n183) );
  CLKINVX1 U74 ( .A(n62), .Y(n184) );
  CLKINVX1 U75 ( .A(n63), .Y(n185) );
  MX2XL U76 ( .A(dataOut[27]), .B(n186), .S0(n150), .Y(n136) );
  CLKINVX1 U77 ( .A(n64), .Y(n186) );
  CLKMX2X2 U78 ( .A(dataOut[28]), .B(n187), .S0(n150), .Y(n137) );
  INVX1 U79 ( .A(n65), .Y(n187) );
  CLKINVX1 U80 ( .A(n66), .Y(n188) );
  CLKINVX1 U81 ( .A(n67), .Y(n189) );
  CLKINVX1 U82 ( .A(n68), .Y(n190) );
  CLKINVX1 U83 ( .A(n45), .Y(n167) );
  CLKINVX1 U84 ( .A(n46), .Y(n168) );
  MX2XL U85 ( .A(ALUout_regE[28]), .B(n219), .S0(n148), .Y(n97) );
  CLKINVX1 U86 ( .A(n30), .Y(n219) );
  MX2XL U87 ( .A(ALUout_regE[24]), .B(n215), .S0(n148), .Y(n93) );
  CLKINVX1 U88 ( .A(n26), .Y(n215) );
  MX2XL U89 ( .A(ALUout_regE[21]), .B(n212), .S0(n149), .Y(n90) );
  CLKINVX1 U90 ( .A(n23), .Y(n212) );
  MX2XL U91 ( .A(ALUout_regE[13]), .B(n204), .S0(n148), .Y(n82) );
  CLKINVX1 U92 ( .A(n15), .Y(n204) );
  MX2XL U93 ( .A(ALUout_regE[16]), .B(n207), .S0(n149), .Y(n85) );
  CLKINVX1 U94 ( .A(n18), .Y(n207) );
  MX2XL U95 ( .A(ALUout_regE[11]), .B(n202), .S0(n148), .Y(n80) );
  CLKINVX1 U96 ( .A(n13), .Y(n202) );
  MX2XL U97 ( .A(ALUout_regE[10]), .B(n201), .S0(n148), .Y(n79) );
  CLKINVX1 U98 ( .A(n12), .Y(n201) );
  MX2XL U99 ( .A(ALUout_regE[2]), .B(n193), .S0(n148), .Y(n71) );
  CLKINVX1 U100 ( .A(n4), .Y(n193) );
  MX2XL U101 ( .A(ALUout_regE[25]), .B(n216), .S0(n151), .Y(n94) );
  CLKINVX1 U102 ( .A(n27), .Y(n216) );
  MX2XL U103 ( .A(ALUout_regE[9]), .B(n200), .S0(n151), .Y(n78) );
  CLKINVX1 U104 ( .A(n11), .Y(n200) );
  MX2XL U105 ( .A(ALUout_regE[22]), .B(n213), .S0(stallcache), .Y(n91) );
  CLKINVX1 U106 ( .A(n24), .Y(n213) );
  MX2XL U107 ( .A(ALUout_regE[27]), .B(n218), .S0(stallcache), .Y(n96) );
  CLKINVX1 U108 ( .A(n29), .Y(n218) );
  MX2XL U109 ( .A(ALUout_regE[7]), .B(n198), .S0(n148), .Y(n76) );
  CLKINVX1 U110 ( .A(n9), .Y(n198) );
  MX2XL U111 ( .A(ALUout_regE[17]), .B(n208), .S0(stallcache), .Y(n86) );
  CLKINVX1 U112 ( .A(n19), .Y(n208) );
  MX2XL U113 ( .A(ALUout_regE[12]), .B(n203), .S0(n150), .Y(n81) );
  CLKINVX1 U114 ( .A(n14), .Y(n203) );
  MX2XL U115 ( .A(ALUout_regE[20]), .B(n211), .S0(stallcache), .Y(n89) );
  CLKINVX1 U116 ( .A(n22), .Y(n211) );
  MX2XL U117 ( .A(ALUout_regE[23]), .B(n214), .S0(stallcache), .Y(n92) );
  CLKINVX1 U118 ( .A(n25), .Y(n214) );
  MX2XL U119 ( .A(ALUout_regE[18]), .B(n209), .S0(stallcache), .Y(n87) );
  CLKINVX1 U120 ( .A(n20), .Y(n209) );
  MX2XL U121 ( .A(ALUout_regE[31]), .B(n222), .S0(n148), .Y(n100) );
  CLKINVX1 U122 ( .A(n33), .Y(n222) );
  MX2XL U123 ( .A(ALUout_regE[14]), .B(n205), .S0(n150), .Y(n83) );
  CLKINVX1 U124 ( .A(n16), .Y(n205) );
  MX2XL U125 ( .A(ALUout_regE[30]), .B(n221), .S0(n148), .Y(n99) );
  CLKINVX1 U126 ( .A(n32), .Y(n221) );
  MX2XL U127 ( .A(ALUout_regE[8]), .B(n199), .S0(n151), .Y(n77) );
  CLKINVX1 U128 ( .A(n10), .Y(n199) );
  MX2XL U129 ( .A(ALUout_regE[3]), .B(n194), .S0(stallcache), .Y(n72) );
  CLKINVX1 U130 ( .A(n5), .Y(n194) );
  MX2XL U131 ( .A(ALUout_regE[29]), .B(n220), .S0(n148), .Y(n98) );
  CLKINVX1 U132 ( .A(n31), .Y(n220) );
  MX2XL U133 ( .A(ALUout_regE[19]), .B(n210), .S0(stallcache), .Y(n88) );
  CLKINVX1 U134 ( .A(n21), .Y(n210) );
  MX2XL U135 ( .A(ALUout_regE[26]), .B(n217), .S0(stallcache), .Y(n95) );
  CLKINVX1 U136 ( .A(n28), .Y(n217) );
  MX2XL U137 ( .A(ALUout_regE[15]), .B(n206), .S0(stallcache), .Y(n84) );
  CLKINVX1 U138 ( .A(n17), .Y(n206) );
  MX2XL U139 ( .A(RegWrite_regE), .B(n223), .S0(n148), .Y(n101) );
  CLKINVX1 U140 ( .A(n34), .Y(n223) );
  CLKINVX1 U141 ( .A(n35), .Y(n224) );
  MX2XL U142 ( .A(MemtoReg_regE[1]), .B(MemtoReg_regM[1]), .S0(n148), .Y(n103)
         );
  MX2XL U143 ( .A(ALUout_regE[4]), .B(n195), .S0(stallcache), .Y(n73) );
  CLKINVX1 U144 ( .A(n6), .Y(n195) );
  MX2XL U145 ( .A(ALUout_regE[5]), .B(n196), .S0(stallcache), .Y(n74) );
  CLKINVX1 U146 ( .A(n7), .Y(n196) );
  MX2XL U147 ( .A(ALUout_regE[6]), .B(n197), .S0(stallcache), .Y(n75) );
  CLKINVX1 U148 ( .A(n8), .Y(n197) );
  MX2XL U149 ( .A(ALUout_regE[0]), .B(n191), .S0(n150), .Y(n69) );
  CLKINVX1 U150 ( .A(n2), .Y(n191) );
  MX2XL U151 ( .A(ALUout_regE[1]), .B(n192), .S0(n150), .Y(n70) );
  CLKINVX1 U152 ( .A(n3), .Y(n192) );
  MX2XL U153 ( .A(wsel_regE[2]), .B(wsel_regM[2]), .S0(n150), .Y(n106) );
  CLKBUFX2 U154 ( .A(stallcache), .Y(n145) );
endmodule


module maincontrol ( opcode, funct, RegDst, MemtoReg, ALUOp, Branch, MemRead, 
        MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp );
  input [5:0] opcode;
  input [5:0] funct;
  output [1:0] RegDst;
  output [1:0] MemtoReg;
  output [5:0] ALUOp;
  output Branch, MemRead, MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n8, n9, n29, n30, n31, n32, n33, n34, n35;

  CLKBUFX2 U3 ( .A(opcode[1]), .Y(ALUOp[1]) );
  OAI221X1 U4 ( .A0(n27), .A1(n32), .B0(n23), .B1(n30), .C0(n28), .Y(n19) );
  CLKINVX8 U5 ( .A(opcode[0]), .Y(n33) );
  CLKINVX3 U6 ( .A(opcode[3]), .Y(n31) );
  AOI31X1 U7 ( .A0(n20), .A1(n32), .A2(opcode[0]), .B0(ALUOp[4]), .Y(n28) );
  CLKINVX6 U8 ( .A(opcode[1]), .Y(n32) );
  NOR2X6 U9 ( .A(n13), .B(ALUOp[4]), .Y(RegDst[1]) );
  CLKINVX8 U10 ( .A(opcode[5]), .Y(n30) );
  INVXL U11 ( .A(n21), .Y(n34) );
  NOR3XL U12 ( .A(n31), .B(ALUOp[4]), .C(n15), .Y(MemWrite) );
  NOR3X2 U13 ( .A(opcode[2]), .B(opcode[3]), .C(n11), .Y(n25) );
  NAND2X4 U14 ( .A(n8), .B(n29), .Y(RegDst[0]) );
  NOR3XL U15 ( .A(n15), .B(ALUOp[4]), .C(opcode[3]), .Y(MemRead) );
  CLKBUFX2 U16 ( .A(opcode[0]), .Y(ALUOp[0]) );
  CLKBUFX2 U17 ( .A(opcode[2]), .Y(ALUOp[2]) );
  CLKBUFX2 U18 ( .A(opcode[3]), .Y(ALUOp[3]) );
  NOR4BXL U19 ( .AN(opcode[2]), .B(ALUOp[4]), .C(opcode[3]), .D(n11), .Y(
        Branch) );
  NAND4X2 U20 ( .A(opcode[1]), .B(n23), .C(n31), .D(n30), .Y(n13) );
  OAI211XL U21 ( .A0(n35), .A1(n29), .B0(n17), .C0(n18), .Y(MemtoReg[0]) );
  NOR2XL U22 ( .A(n19), .B(n14), .Y(n18) );
  NAND3X2 U23 ( .A(n21), .B(n22), .C(funct[3]), .Y(n16) );
  BUFX8 U24 ( .A(opcode[4]), .Y(ALUOp[4]) );
  NAND3XL U25 ( .A(opcode[1]), .B(n23), .C(opcode[5]), .Y(n15) );
  NOR3XL U26 ( .A(ALUOp[4]), .B(funct[1]), .C(n34), .Y(n24) );
  CLKBUFX3 U27 ( .A(RegDst[0]), .Y(ExtOp) );
  OAI31XL U28 ( .A0(n29), .A1(ALUOp[4]), .A2(n16), .B0(n9), .Y(MemtoReg[1]) );
  CLKINVX1 U29 ( .A(RegDst[1]), .Y(n9) );
  CLKINVX1 U30 ( .A(n19), .Y(n8) );
  NAND3X1 U31 ( .A(n32), .B(n30), .C(n33), .Y(n11) );
  CLKINVX1 U32 ( .A(n25), .Y(n29) );
  CLKBUFX3 U33 ( .A(opcode[5]), .Y(ALUOp[5]) );
  AND3X2 U34 ( .A(funct[3]), .B(n24), .C(n25), .Y(JumpReg) );
  NAND3XL U35 ( .A(n26), .B(n13), .C(n8), .Y(ALUsrc) );
  OAI31XL U36 ( .A0(n34), .A1(funct[3]), .A2(n22), .B0(n25), .Y(n26) );
  NOR2BX1 U37 ( .AN(n10), .B(ALUOp[4]), .Y(RegWrite) );
  AOI32X1 U38 ( .A0(opcode[0]), .A1(n30), .A2(opcode[3]), .B0(opcode[2]), .B1(
        n31), .Y(n27) );
  OAI22XL U39 ( .A0(opcode[0]), .A1(n31), .B0(opcode[1]), .B1(n20), .Y(n14) );
  NOR3X1 U40 ( .A(funct[5]), .B(funct[4]), .C(funct[2]), .Y(n21) );
  OAI211XL U41 ( .A0(n11), .A1(opcode[2]), .B0(n12), .C0(n13), .Y(n10) );
  AOI2BB2XL U42 ( .B0(n30), .B1(n14), .A0N(opcode[3]), .A1N(n15), .Y(n12) );
  NOR2X1 U43 ( .A(n33), .B(opcode[2]), .Y(n23) );
  NOR2BX1 U44 ( .AN(funct[0]), .B(funct[1]), .Y(n22) );
  NAND2X1 U45 ( .A(opcode[3]), .B(opcode[2]), .Y(n20) );
  OAI21XL U46 ( .A0(opcode[2]), .A1(opcode[1]), .B0(n33), .Y(n17) );
  CLKINVX1 U47 ( .A(n16), .Y(n35) );
endmodule


module registerFile ( clk, rst_n, rsel1, rsel2, wsel, wen, wdata, rdata1, 
        rdata2 );
  input [4:0] rsel1;
  input [4:0] rsel2;
  input [4:0] wsel;
  input [31:0] wdata;
  output [31:0] rdata1;
  output [31:0] rdata2;
  input clk, rst_n, wen;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, \register[31][31] ,
         \register[31][30] , \register[31][29] , \register[31][28] ,
         \register[31][27] , \register[31][26] , \register[31][25] ,
         \register[31][24] , \register[31][23] , \register[31][22] ,
         \register[31][21] , \register[31][20] , \register[31][19] ,
         \register[31][18] , \register[31][17] , \register[31][16] ,
         \register[31][15] , \register[31][14] , \register[31][13] ,
         \register[31][12] , \register[31][11] , \register[31][10] ,
         \register[31][9] , \register[31][8] , \register[31][7] ,
         \register[31][6] , \register[31][5] , \register[31][4] ,
         \register[31][3] , \register[31][2] , \register[31][1] ,
         \register[31][0] , \register[30][31] , \register[30][30] ,
         \register[30][29] , \register[30][28] , \register[30][27] ,
         \register[30][26] , \register[30][25] , \register[30][24] ,
         \register[30][23] , \register[30][22] , \register[30][21] ,
         \register[30][20] , \register[30][19] , \register[30][18] ,
         \register[30][17] , \register[30][16] , \register[30][15] ,
         \register[30][14] , \register[30][13] , \register[30][12] ,
         \register[30][11] , \register[30][10] , \register[30][9] ,
         \register[30][8] , \register[30][7] , \register[30][6] ,
         \register[30][5] , \register[30][4] , \register[30][3] ,
         \register[30][2] , \register[30][1] , \register[30][0] ,
         \register[29][31] , \register[29][30] , \register[29][29] ,
         \register[29][28] , \register[29][27] , \register[29][26] ,
         \register[29][25] , \register[29][24] , \register[29][23] ,
         \register[29][22] , \register[29][21] , \register[29][20] ,
         \register[29][19] , \register[29][18] , \register[29][17] ,
         \register[29][16] , \register[29][15] , \register[29][14] ,
         \register[29][13] , \register[29][12] , \register[29][11] ,
         \register[29][10] , \register[29][9] , \register[29][8] ,
         \register[29][7] , \register[29][6] , \register[29][5] ,
         \register[29][4] , \register[29][3] , \register[29][2] ,
         \register[29][1] , \register[29][0] , \register[28][31] ,
         \register[28][30] , \register[28][29] , \register[28][28] ,
         \register[28][27] , \register[28][26] , \register[28][25] ,
         \register[28][24] , \register[28][23] , \register[28][22] ,
         \register[28][21] , \register[28][20] , \register[28][19] ,
         \register[28][18] , \register[28][17] , \register[28][16] ,
         \register[28][15] , \register[28][14] , \register[28][13] ,
         \register[28][12] , \register[28][11] , \register[28][10] ,
         \register[28][9] , \register[28][8] , \register[28][7] ,
         \register[28][6] , \register[28][5] , \register[28][4] ,
         \register[28][3] , \register[28][2] , \register[28][1] ,
         \register[28][0] , \register[27][31] , \register[27][30] ,
         \register[27][29] , \register[27][28] , \register[27][27] ,
         \register[27][26] , \register[27][25] , \register[27][24] ,
         \register[27][23] , \register[27][22] , \register[27][21] ,
         \register[27][20] , \register[27][19] , \register[27][18] ,
         \register[27][17] , \register[27][16] , \register[27][15] ,
         \register[27][14] , \register[27][13] , \register[27][12] ,
         \register[27][11] , \register[27][10] , \register[27][9] ,
         \register[27][8] , \register[27][7] , \register[27][6] ,
         \register[27][5] , \register[27][4] , \register[27][3] ,
         \register[27][2] , \register[27][1] , \register[27][0] ,
         \register[26][31] , \register[26][30] , \register[26][29] ,
         \register[26][28] , \register[26][27] , \register[26][26] ,
         \register[26][25] , \register[26][24] , \register[26][23] ,
         \register[26][22] , \register[26][21] , \register[26][20] ,
         \register[26][19] , \register[26][18] , \register[26][17] ,
         \register[26][16] , \register[26][15] , \register[26][14] ,
         \register[26][13] , \register[26][12] , \register[26][11] ,
         \register[26][10] , \register[26][9] , \register[26][8] ,
         \register[26][7] , \register[26][6] , \register[26][5] ,
         \register[26][4] , \register[26][3] , \register[26][2] ,
         \register[26][1] , \register[26][0] , \register[25][31] ,
         \register[25][30] , \register[25][29] , \register[25][28] ,
         \register[25][27] , \register[25][26] , \register[25][25] ,
         \register[25][24] , \register[25][23] , \register[25][22] ,
         \register[25][21] , \register[25][20] , \register[25][19] ,
         \register[25][18] , \register[25][17] , \register[25][16] ,
         \register[25][15] , \register[25][14] , \register[25][13] ,
         \register[25][12] , \register[25][11] , \register[25][10] ,
         \register[25][9] , \register[25][8] , \register[25][7] ,
         \register[25][6] , \register[25][5] , \register[25][4] ,
         \register[25][3] , \register[25][2] , \register[25][1] ,
         \register[25][0] , \register[24][31] , \register[24][30] ,
         \register[24][29] , \register[24][28] , \register[24][27] ,
         \register[24][26] , \register[24][25] , \register[24][24] ,
         \register[24][23] , \register[24][22] , \register[24][21] ,
         \register[24][20] , \register[24][19] , \register[24][18] ,
         \register[24][17] , \register[24][16] , \register[24][15] ,
         \register[24][14] , \register[24][13] , \register[24][12] ,
         \register[24][11] , \register[24][10] , \register[24][9] ,
         \register[24][8] , \register[24][7] , \register[24][6] ,
         \register[24][5] , \register[24][4] , \register[24][3] ,
         \register[24][2] , \register[24][1] , \register[24][0] ,
         \register[23][31] , \register[23][30] , \register[23][29] ,
         \register[23][28] , \register[23][27] , \register[23][26] ,
         \register[23][25] , \register[23][24] , \register[23][23] ,
         \register[23][22] , \register[23][21] , \register[23][20] ,
         \register[23][19] , \register[23][18] , \register[23][17] ,
         \register[23][16] , \register[23][15] , \register[23][14] ,
         \register[23][13] , \register[23][12] , \register[23][11] ,
         \register[23][10] , \register[23][9] , \register[23][8] ,
         \register[23][7] , \register[23][6] , \register[23][5] ,
         \register[23][4] , \register[23][3] , \register[23][2] ,
         \register[23][1] , \register[23][0] , \register[22][31] ,
         \register[22][30] , \register[22][29] , \register[22][28] ,
         \register[22][27] , \register[22][26] , \register[22][25] ,
         \register[22][24] , \register[22][23] , \register[22][22] ,
         \register[22][21] , \register[22][20] , \register[22][19] ,
         \register[22][18] , \register[22][17] , \register[22][16] ,
         \register[22][15] , \register[22][14] , \register[22][13] ,
         \register[22][12] , \register[22][11] , \register[22][10] ,
         \register[22][9] , \register[22][8] , \register[22][7] ,
         \register[22][6] , \register[22][5] , \register[22][4] ,
         \register[22][3] , \register[22][2] , \register[22][1] ,
         \register[22][0] , \register[21][31] , \register[21][30] ,
         \register[21][29] , \register[21][28] , \register[21][27] ,
         \register[21][26] , \register[21][25] , \register[21][24] ,
         \register[21][23] , \register[21][22] , \register[21][21] ,
         \register[21][20] , \register[21][19] , \register[21][18] ,
         \register[21][17] , \register[21][16] , \register[21][15] ,
         \register[21][14] , \register[21][13] , \register[21][12] ,
         \register[21][11] , \register[21][10] , \register[21][9] ,
         \register[21][8] , \register[21][7] , \register[21][6] ,
         \register[21][5] , \register[21][4] , \register[21][3] ,
         \register[21][2] , \register[21][1] , \register[21][0] ,
         \register[20][31] , \register[20][30] , \register[20][29] ,
         \register[20][28] , \register[20][27] , \register[20][26] ,
         \register[20][25] , \register[20][24] , \register[20][23] ,
         \register[20][22] , \register[20][21] , \register[20][20] ,
         \register[20][19] , \register[20][18] , \register[20][17] ,
         \register[20][16] , \register[20][15] , \register[20][14] ,
         \register[20][13] , \register[20][12] , \register[20][11] ,
         \register[20][10] , \register[20][9] , \register[20][8] ,
         \register[20][7] , \register[20][6] , \register[20][5] ,
         \register[20][4] , \register[20][3] , \register[20][2] ,
         \register[20][1] , \register[20][0] , \register[19][31] ,
         \register[19][30] , \register[19][29] , \register[19][28] ,
         \register[19][27] , \register[19][26] , \register[19][25] ,
         \register[19][24] , \register[19][23] , \register[19][22] ,
         \register[19][21] , \register[19][20] , \register[19][19] ,
         \register[19][18] , \register[19][17] , \register[19][16] ,
         \register[19][15] , \register[19][14] , \register[19][13] ,
         \register[19][12] , \register[19][11] , \register[19][10] ,
         \register[19][9] , \register[19][8] , \register[19][7] ,
         \register[19][6] , \register[19][5] , \register[19][4] ,
         \register[19][3] , \register[19][2] , \register[19][1] ,
         \register[19][0] , \register[18][31] , \register[18][30] ,
         \register[18][29] , \register[18][28] , \register[18][27] ,
         \register[18][26] , \register[18][25] , \register[18][24] ,
         \register[18][23] , \register[18][22] , \register[18][21] ,
         \register[18][20] , \register[18][19] , \register[18][18] ,
         \register[18][17] , \register[18][16] , \register[18][15] ,
         \register[18][14] , \register[18][13] , \register[18][12] ,
         \register[18][11] , \register[18][10] , \register[18][9] ,
         \register[18][8] , \register[18][7] , \register[18][6] ,
         \register[18][5] , \register[18][4] , \register[18][3] ,
         \register[18][2] , \register[18][1] , \register[18][0] ,
         \register[17][31] , \register[17][30] , \register[17][29] ,
         \register[17][28] , \register[17][27] , \register[17][26] ,
         \register[17][25] , \register[17][24] , \register[17][23] ,
         \register[17][22] , \register[17][21] , \register[17][20] ,
         \register[17][19] , \register[17][18] , \register[17][17] ,
         \register[17][16] , \register[17][15] , \register[17][14] ,
         \register[17][13] , \register[17][12] , \register[17][11] ,
         \register[17][10] , \register[17][9] , \register[17][8] ,
         \register[17][7] , \register[17][6] , \register[17][5] ,
         \register[17][4] , \register[17][3] , \register[17][2] ,
         \register[17][1] , \register[17][0] , \register[16][31] ,
         \register[16][30] , \register[16][29] , \register[16][28] ,
         \register[16][27] , \register[16][26] , \register[16][25] ,
         \register[16][24] , \register[16][23] , \register[16][22] ,
         \register[16][21] , \register[16][20] , \register[16][19] ,
         \register[16][18] , \register[16][17] , \register[16][16] ,
         \register[16][15] , \register[16][14] , \register[16][13] ,
         \register[16][12] , \register[16][11] , \register[16][10] ,
         \register[16][9] , \register[16][8] , \register[16][7] ,
         \register[16][6] , \register[16][5] , \register[16][4] ,
         \register[16][3] , \register[16][2] , \register[16][1] ,
         \register[16][0] , \register[15][31] , \register[15][30] ,
         \register[15][29] , \register[15][28] , \register[15][27] ,
         \register[15][26] , \register[15][25] , \register[15][24] ,
         \register[15][23] , \register[15][22] , \register[15][21] ,
         \register[15][20] , \register[15][19] , \register[15][18] ,
         \register[15][17] , \register[15][16] , \register[15][15] ,
         \register[15][14] , \register[15][13] , \register[15][12] ,
         \register[15][11] , \register[15][10] , \register[15][9] ,
         \register[15][8] , \register[15][7] , \register[15][6] ,
         \register[15][5] , \register[15][4] , \register[15][3] ,
         \register[15][2] , \register[15][1] , \register[15][0] ,
         \register[14][31] , \register[14][30] , \register[14][29] ,
         \register[14][28] , \register[14][27] , \register[14][26] ,
         \register[14][25] , \register[14][24] , \register[14][23] ,
         \register[14][22] , \register[14][21] , \register[14][20] ,
         \register[14][19] , \register[14][18] , \register[14][17] ,
         \register[14][16] , \register[14][15] , \register[14][14] ,
         \register[14][13] , \register[14][12] , \register[14][11] ,
         \register[14][10] , \register[14][9] , \register[14][8] ,
         \register[14][7] , \register[14][6] , \register[14][5] ,
         \register[14][4] , \register[14][3] , \register[14][2] ,
         \register[14][1] , \register[14][0] , \register[13][31] ,
         \register[13][30] , \register[13][29] , \register[13][28] ,
         \register[13][27] , \register[13][26] , \register[13][25] ,
         \register[13][24] , \register[13][23] , \register[13][22] ,
         \register[13][21] , \register[13][20] , \register[13][19] ,
         \register[13][18] , \register[13][17] , \register[13][16] ,
         \register[13][15] , \register[13][14] , \register[13][13] ,
         \register[13][12] , \register[13][11] , \register[13][10] ,
         \register[13][9] , \register[13][8] , \register[13][7] ,
         \register[13][6] , \register[13][5] , \register[13][4] ,
         \register[13][3] , \register[13][2] , \register[13][1] ,
         \register[13][0] , \register[12][31] , \register[12][30] ,
         \register[12][29] , \register[12][28] , \register[12][27] ,
         \register[12][26] , \register[12][25] , \register[12][24] ,
         \register[12][23] , \register[12][22] , \register[12][21] ,
         \register[12][20] , \register[12][19] , \register[12][18] ,
         \register[12][17] , \register[12][16] , \register[12][15] ,
         \register[12][14] , \register[12][13] , \register[12][12] ,
         \register[12][11] , \register[12][10] , \register[12][9] ,
         \register[12][8] , \register[12][7] , \register[12][6] ,
         \register[12][5] , \register[12][4] , \register[12][3] ,
         \register[12][2] , \register[12][1] , \register[12][0] ,
         \register[11][31] , \register[11][30] , \register[11][29] ,
         \register[11][28] , \register[11][27] , \register[11][26] ,
         \register[11][25] , \register[11][24] , \register[11][23] ,
         \register[11][22] , \register[11][21] , \register[11][20] ,
         \register[11][19] , \register[11][18] , \register[11][17] ,
         \register[11][16] , \register[11][15] , \register[11][14] ,
         \register[11][13] , \register[11][12] , \register[11][11] ,
         \register[11][10] , \register[11][9] , \register[11][8] ,
         \register[11][7] , \register[11][6] , \register[11][5] ,
         \register[11][4] , \register[11][3] , \register[11][2] ,
         \register[11][1] , \register[11][0] , \register[10][31] ,
         \register[10][30] , \register[10][29] , \register[10][28] ,
         \register[10][27] , \register[10][26] , \register[10][25] ,
         \register[10][24] , \register[10][23] , \register[10][22] ,
         \register[10][21] , \register[10][20] , \register[10][19] ,
         \register[10][18] , \register[10][17] , \register[10][16] ,
         \register[10][15] , \register[10][14] , \register[10][13] ,
         \register[10][12] , \register[10][11] , \register[10][10] ,
         \register[10][9] , \register[10][8] , \register[10][7] ,
         \register[10][6] , \register[10][5] , \register[10][4] ,
         \register[10][3] , \register[10][2] , \register[10][1] ,
         \register[10][0] , \register[9][31] , \register[9][30] ,
         \register[9][29] , \register[9][28] , \register[9][27] ,
         \register[9][26] , \register[9][25] , \register[9][24] ,
         \register[9][23] , \register[9][22] , \register[9][21] ,
         \register[9][20] , \register[9][19] , \register[9][18] ,
         \register[9][17] , \register[9][16] , \register[9][15] ,
         \register[9][14] , \register[9][13] , \register[9][12] ,
         \register[9][11] , \register[9][10] , \register[9][9] ,
         \register[9][8] , \register[9][7] , \register[9][6] ,
         \register[9][5] , \register[9][4] , \register[9][3] ,
         \register[9][2] , \register[9][1] , \register[9][0] ,
         \register[8][31] , \register[8][30] , \register[8][29] ,
         \register[8][28] , \register[8][27] , \register[8][26] ,
         \register[8][25] , \register[8][24] , \register[8][23] ,
         \register[8][22] , \register[8][21] , \register[8][20] ,
         \register[8][19] , \register[8][18] , \register[8][17] ,
         \register[8][16] , \register[8][15] , \register[8][14] ,
         \register[8][13] , \register[8][12] , \register[8][11] ,
         \register[8][10] , \register[8][9] , \register[8][8] ,
         \register[8][7] , \register[8][6] , \register[8][5] ,
         \register[8][4] , \register[8][3] , \register[8][2] ,
         \register[8][1] , \register[8][0] , \register[7][31] ,
         \register[7][30] , \register[7][29] , \register[7][28] ,
         \register[7][27] , \register[7][26] , \register[7][25] ,
         \register[7][24] , \register[7][23] , \register[7][22] ,
         \register[7][21] , \register[7][20] , \register[7][19] ,
         \register[7][18] , \register[7][17] , \register[7][16] ,
         \register[7][15] , \register[7][14] , \register[7][13] ,
         \register[7][12] , \register[7][11] , \register[7][10] ,
         \register[7][9] , \register[7][8] , \register[7][7] ,
         \register[7][6] , \register[7][5] , \register[7][4] ,
         \register[7][3] , \register[7][2] , \register[7][1] ,
         \register[7][0] , \register[6][31] , \register[6][30] ,
         \register[6][29] , \register[6][28] , \register[6][27] ,
         \register[6][26] , \register[6][25] , \register[6][24] ,
         \register[6][23] , \register[6][22] , \register[6][21] ,
         \register[6][20] , \register[6][19] , \register[6][18] ,
         \register[6][17] , \register[6][16] , \register[6][15] ,
         \register[6][14] , \register[6][13] , \register[6][12] ,
         \register[6][11] , \register[6][10] , \register[6][9] ,
         \register[6][8] , \register[6][7] , \register[6][6] ,
         \register[6][5] , \register[6][4] , \register[6][3] ,
         \register[6][2] , \register[6][1] , \register[6][0] ,
         \register[5][31] , \register[5][30] , \register[5][29] ,
         \register[5][28] , \register[5][27] , \register[5][26] ,
         \register[5][25] , \register[5][24] , \register[5][23] ,
         \register[5][22] , \register[5][21] , \register[5][20] ,
         \register[5][19] , \register[5][18] , \register[5][17] ,
         \register[5][16] , \register[5][15] , \register[5][14] ,
         \register[5][13] , \register[5][12] , \register[5][11] ,
         \register[5][10] , \register[5][9] , \register[5][8] ,
         \register[5][7] , \register[5][6] , \register[5][5] ,
         \register[5][4] , \register[5][3] , \register[5][2] ,
         \register[5][1] , \register[5][0] , \register[4][31] ,
         \register[4][30] , \register[4][29] , \register[4][28] ,
         \register[4][27] , \register[4][26] , \register[4][25] ,
         \register[4][24] , \register[4][23] , \register[4][22] ,
         \register[4][21] , \register[4][20] , \register[4][19] ,
         \register[4][18] , \register[4][17] , \register[4][16] ,
         \register[4][15] , \register[4][14] , \register[4][13] ,
         \register[4][12] , \register[4][11] , \register[4][10] ,
         \register[4][9] , \register[4][8] , \register[4][7] ,
         \register[4][6] , \register[4][5] , \register[4][4] ,
         \register[4][3] , \register[4][2] , \register[4][1] ,
         \register[4][0] , \register[3][31] , \register[3][30] ,
         \register[3][29] , \register[3][28] , \register[3][27] ,
         \register[3][26] , \register[3][25] , \register[3][24] ,
         \register[3][23] , \register[3][22] , \register[3][21] ,
         \register[3][20] , \register[3][19] , \register[3][18] ,
         \register[3][17] , \register[3][16] , \register[3][15] ,
         \register[3][14] , \register[3][13] , \register[3][12] ,
         \register[3][11] , \register[3][10] , \register[3][9] ,
         \register[3][8] , \register[3][7] , \register[3][6] ,
         \register[3][5] , \register[3][4] , \register[3][3] ,
         \register[3][2] , \register[3][1] , \register[3][0] ,
         \register[2][31] , \register[2][30] , \register[2][29] ,
         \register[2][28] , \register[2][27] , \register[2][26] ,
         \register[2][25] , \register[2][24] , \register[2][23] ,
         \register[2][22] , \register[2][21] , \register[2][20] ,
         \register[2][19] , \register[2][18] , \register[2][17] ,
         \register[2][16] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[1][31] ,
         \register[1][30] , \register[1][29] , \register[1][28] ,
         \register[1][27] , \register[1][26] , \register[1][25] ,
         \register[1][24] , \register[1][23] , \register[1][22] ,
         \register[1][21] , \register[1][20] , \register[1][19] ,
         \register[1][18] , \register[1][17] , \register[1][16] ,
         \register[1][15] , \register[1][14] , \register[1][13] ,
         \register[1][12] , \register[1][11] , \register[1][10] ,
         \register[1][9] , \register[1][8] , \register[1][7] ,
         \register[1][6] , \register[1][5] , \register[1][4] ,
         \register[1][3] , \register[1][2] , \register[1][1] ,
         \register[1][0] , N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n67, n68, n69, n70, n71, n72, n74, n76, n77, n78, n79,
         n80, n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n66, n73, n75, n82, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
  assign N12 = rsel1[0];
  assign N13 = rsel1[1];
  assign N14 = rsel1[2];
  assign N15 = rsel1[3];
  assign N16 = rsel1[4];
  assign N17 = rsel2[0];
  assign N18 = rsel2[1];
  assign N19 = rsel2[2];
  assign N20 = rsel2[3];
  assign N21 = rsel2[4];

  NOR3X4 U878 ( .A(n14), .B(wsel[3]), .C(n2621), .Y(n91) );
  DFFRX1 \register_reg[2][31]  ( .D(n171), .CK(clk), .RN(n2454), .Q(
        \register[2][31] ), .QN(n2585) );
  DFFRX1 \register_reg[2][30]  ( .D(n170), .CK(clk), .RN(n2454), .Q(
        \register[2][30] ), .QN(n2584) );
  DFFRX1 \register_reg[2][29]  ( .D(n169), .CK(clk), .RN(n2454), .Q(
        \register[2][29] ), .QN(n2583) );
  DFFRX1 \register_reg[2][28]  ( .D(n168), .CK(clk), .RN(n2454), .Q(
        \register[2][28] ), .QN(n2582) );
  DFFRX1 \register_reg[2][27]  ( .D(n167), .CK(clk), .RN(n2453), .Q(
        \register[2][27] ), .QN(n2581) );
  DFFRX1 \register_reg[2][26]  ( .D(n166), .CK(clk), .RN(n2453), .Q(
        \register[2][26] ), .QN(n2580) );
  DFFRX1 \register_reg[2][25]  ( .D(n165), .CK(clk), .RN(n2453), .Q(
        \register[2][25] ), .QN(n2579) );
  DFFRX1 \register_reg[2][24]  ( .D(n164), .CK(clk), .RN(n2453), .Q(
        \register[2][24] ), .QN(n2578) );
  DFFRX1 \register_reg[2][23]  ( .D(n163), .CK(clk), .RN(n2453), .Q(
        \register[2][23] ), .QN(n2577) );
  DFFRX1 \register_reg[2][22]  ( .D(n162), .CK(clk), .RN(n2453), .Q(
        \register[2][22] ), .QN(n2576) );
  DFFRX1 \register_reg[2][21]  ( .D(n161), .CK(clk), .RN(n2453), .Q(
        \register[2][21] ), .QN(n2575) );
  DFFRX1 \register_reg[2][20]  ( .D(n160), .CK(clk), .RN(n2453), .Q(
        \register[2][20] ), .QN(n2574) );
  DFFRX1 \register_reg[2][19]  ( .D(n159), .CK(clk), .RN(n2453), .Q(
        \register[2][19] ), .QN(n2573) );
  DFFRX1 \register_reg[2][18]  ( .D(n158), .CK(clk), .RN(n2453), .Q(
        \register[2][18] ), .QN(n2572) );
  DFFRX1 \register_reg[2][17]  ( .D(n157), .CK(clk), .RN(n2453), .Q(
        \register[2][17] ), .QN(n2571) );
  DFFRX1 \register_reg[2][16]  ( .D(n156), .CK(clk), .RN(n2453), .Q(
        \register[2][16] ), .QN(n2570) );
  DFFRX1 \register_reg[2][15]  ( .D(n155), .CK(clk), .RN(n2452), .Q(
        \register[2][15] ), .QN(n2569) );
  DFFRX1 \register_reg[2][14]  ( .D(n154), .CK(clk), .RN(n2452), .Q(
        \register[2][14] ), .QN(n2568) );
  DFFRX1 \register_reg[2][13]  ( .D(n153), .CK(clk), .RN(n2452), .Q(
        \register[2][13] ), .QN(n2567) );
  DFFRX1 \register_reg[2][12]  ( .D(n152), .CK(clk), .RN(n2452), .Q(
        \register[2][12] ), .QN(n2566) );
  DFFRX1 \register_reg[2][11]  ( .D(n151), .CK(clk), .RN(n2452), .Q(
        \register[2][11] ), .QN(n2565) );
  DFFRX1 \register_reg[2][10]  ( .D(n150), .CK(clk), .RN(n2452), .Q(
        \register[2][10] ), .QN(n2564) );
  DFFRX1 \register_reg[2][9]  ( .D(n149), .CK(clk), .RN(n2452), .Q(
        \register[2][9] ), .QN(n2563) );
  DFFRX1 \register_reg[2][8]  ( .D(n148), .CK(clk), .RN(n2452), .Q(
        \register[2][8] ), .QN(n2562) );
  DFFRX1 \register_reg[2][7]  ( .D(n147), .CK(clk), .RN(n2452), .Q(
        \register[2][7] ), .QN(n2561) );
  DFFRX1 \register_reg[2][6]  ( .D(n146), .CK(clk), .RN(n2452), .Q(
        \register[2][6] ), .QN(n2560) );
  DFFRX1 \register_reg[2][5]  ( .D(n145), .CK(clk), .RN(n2452), .Q(
        \register[2][5] ), .QN(n2559) );
  DFFRX1 \register_reg[2][4]  ( .D(n144), .CK(clk), .RN(n2452), .Q(
        \register[2][4] ), .QN(n2558) );
  DFFRX1 \register_reg[2][3]  ( .D(n143), .CK(clk), .RN(n2451), .Q(
        \register[2][3] ), .QN(n2557) );
  DFFRX1 \register_reg[2][2]  ( .D(n142), .CK(clk), .RN(n2451), .Q(
        \register[2][2] ), .QN(n2556) );
  DFFRX1 \register_reg[2][1]  ( .D(n141), .CK(clk), .RN(n2451), .Q(
        \register[2][1] ), .QN(n2555) );
  DFFRX1 \register_reg[2][0]  ( .D(n140), .CK(clk), .RN(n2451), .Q(
        \register[2][0] ), .QN(n2554) );
  DFFRX1 \register_reg[31][31]  ( .D(n1099), .CK(clk), .RN(n2531), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n1098), .CK(clk), .RN(n2531), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n1097), .CK(clk), .RN(n2531), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n1096), .CK(clk), .RN(n2531), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n1095), .CK(clk), .RN(n2531), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n1094), .CK(clk), .RN(n2531), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n1093), .CK(clk), .RN(n2531), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n1092), .CK(clk), .RN(n2531), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n1091), .CK(clk), .RN(n2530), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n1090), .CK(clk), .RN(n2530), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n1089), .CK(clk), .RN(n2530), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n1088), .CK(clk), .RN(n2530), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n1087), .CK(clk), .RN(n2530), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n1086), .CK(clk), .RN(n2530), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n1085), .CK(clk), .RN(n2530), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n1084), .CK(clk), .RN(n2530), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n1083), .CK(clk), .RN(n2530), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n1082), .CK(clk), .RN(n2530), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n1081), .CK(clk), .RN(n2530), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n1080), .CK(clk), .RN(n2530), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n1079), .CK(clk), .RN(n2529), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n1078), .CK(clk), .RN(n2529), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n1077), .CK(clk), .RN(n2529), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n1076), .CK(clk), .RN(n2529), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n1075), .CK(clk), .RN(n2529), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n1074), .CK(clk), .RN(n2529), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n1073), .CK(clk), .RN(n2529), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n1072), .CK(clk), .RN(n2529), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n1071), .CK(clk), .RN(n2529), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n1070), .CK(clk), .RN(n2529), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n1069), .CK(clk), .RN(n2529), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n1068), .CK(clk), .RN(n2529), .Q(
        \register[31][0] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n971), .CK(clk), .RN(n2520), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n970), .CK(clk), .RN(n2520), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n969), .CK(clk), .RN(n2520), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n968), .CK(clk), .RN(n2520), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n967), .CK(clk), .RN(n2520), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n966), .CK(clk), .RN(n2520), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n965), .CK(clk), .RN(n2520), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n964), .CK(clk), .RN(n2520), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n963), .CK(clk), .RN(n2520), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n962), .CK(clk), .RN(n2520), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n961), .CK(clk), .RN(n2520), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n960), .CK(clk), .RN(n2520), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n959), .CK(clk), .RN(n2519), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n958), .CK(clk), .RN(n2519), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n957), .CK(clk), .RN(n2519), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n956), .CK(clk), .RN(n2519), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n955), .CK(clk), .RN(n2519), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n954), .CK(clk), .RN(n2519), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n953), .CK(clk), .RN(n2519), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n952), .CK(clk), .RN(n2519), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n951), .CK(clk), .RN(n2519), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n950), .CK(clk), .RN(n2519), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n949), .CK(clk), .RN(n2519), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n948), .CK(clk), .RN(n2519), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n947), .CK(clk), .RN(n2518), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n946), .CK(clk), .RN(n2518), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n945), .CK(clk), .RN(n2518), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n944), .CK(clk), .RN(n2518), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n943), .CK(clk), .RN(n2518), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n942), .CK(clk), .RN(n2518), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n941), .CK(clk), .RN(n2518), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n940), .CK(clk), .RN(n2518), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n843), .CK(clk), .RN(n2510), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n842), .CK(clk), .RN(n2510), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n841), .CK(clk), .RN(n2510), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n840), .CK(clk), .RN(n2510), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n839), .CK(clk), .RN(n2509), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n838), .CK(clk), .RN(n2509), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n837), .CK(clk), .RN(n2509), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n836), .CK(clk), .RN(n2509), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n835), .CK(clk), .RN(n2509), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n834), .CK(clk), .RN(n2509), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n833), .CK(clk), .RN(n2509), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n832), .CK(clk), .RN(n2509), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n831), .CK(clk), .RN(n2509), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n830), .CK(clk), .RN(n2509), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n829), .CK(clk), .RN(n2509), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n828), .CK(clk), .RN(n2509), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n827), .CK(clk), .RN(n2508), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n826), .CK(clk), .RN(n2508), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n825), .CK(clk), .RN(n2508), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n824), .CK(clk), .RN(n2508), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n823), .CK(clk), .RN(n2508), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n822), .CK(clk), .RN(n2508), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n821), .CK(clk), .RN(n2508), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n820), .CK(clk), .RN(n2508), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n819), .CK(clk), .RN(n2508), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n818), .CK(clk), .RN(n2508), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n817), .CK(clk), .RN(n2508), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n816), .CK(clk), .RN(n2508), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n815), .CK(clk), .RN(n2507), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n814), .CK(clk), .RN(n2507), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n813), .CK(clk), .RN(n2507), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n812), .CK(clk), .RN(n2507), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n715), .CK(clk), .RN(n2499), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n714), .CK(clk), .RN(n2499), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n713), .CK(clk), .RN(n2499), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n712), .CK(clk), .RN(n2499), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n711), .CK(clk), .RN(n2499), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n710), .CK(clk), .RN(n2499), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n709), .CK(clk), .RN(n2499), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n708), .CK(clk), .RN(n2499), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n707), .CK(clk), .RN(n2498), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n706), .CK(clk), .RN(n2498), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n705), .CK(clk), .RN(n2498), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n704), .CK(clk), .RN(n2498), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n703), .CK(clk), .RN(n2498), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n702), .CK(clk), .RN(n2498), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n701), .CK(clk), .RN(n2498), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n700), .CK(clk), .RN(n2498), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n699), .CK(clk), .RN(n2498), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n698), .CK(clk), .RN(n2498), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n697), .CK(clk), .RN(n2498), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n696), .CK(clk), .RN(n2498), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n695), .CK(clk), .RN(n2497), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n694), .CK(clk), .RN(n2497), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n693), .CK(clk), .RN(n2497), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n692), .CK(clk), .RN(n2497), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n691), .CK(clk), .RN(n2497), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n690), .CK(clk), .RN(n2497), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n689), .CK(clk), .RN(n2497), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n688), .CK(clk), .RN(n2497), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n687), .CK(clk), .RN(n2497), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n686), .CK(clk), .RN(n2497), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n685), .CK(clk), .RN(n2497), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n684), .CK(clk), .RN(n2497), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n587), .CK(clk), .RN(n2488), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n586), .CK(clk), .RN(n2488), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n585), .CK(clk), .RN(n2488), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n584), .CK(clk), .RN(n2488), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n583), .CK(clk), .RN(n2488), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n582), .CK(clk), .RN(n2488), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n581), .CK(clk), .RN(n2488), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n580), .CK(clk), .RN(n2488), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n579), .CK(clk), .RN(n2488), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n578), .CK(clk), .RN(n2488), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n577), .CK(clk), .RN(n2488), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n576), .CK(clk), .RN(n2488), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n575), .CK(clk), .RN(n2487), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n574), .CK(clk), .RN(n2487), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n573), .CK(clk), .RN(n2487), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n572), .CK(clk), .RN(n2487), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n571), .CK(clk), .RN(n2487), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n570), .CK(clk), .RN(n2487), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n569), .CK(clk), .RN(n2487), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n568), .CK(clk), .RN(n2487), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n567), .CK(clk), .RN(n2487), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n566), .CK(clk), .RN(n2487), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n565), .CK(clk), .RN(n2487), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n564), .CK(clk), .RN(n2487), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n563), .CK(clk), .RN(n2486), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n562), .CK(clk), .RN(n2486), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n561), .CK(clk), .RN(n2486), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n560), .CK(clk), .RN(n2486), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n559), .CK(clk), .RN(n2486), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n558), .CK(clk), .RN(n2486), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n557), .CK(clk), .RN(n2486), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n556), .CK(clk), .RN(n2486), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n459), .CK(clk), .RN(n2478), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n458), .CK(clk), .RN(n2478), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n457), .CK(clk), .RN(n2478), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n456), .CK(clk), .RN(n2478), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n455), .CK(clk), .RN(n2477), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n454), .CK(clk), .RN(n2477), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n453), .CK(clk), .RN(n2477), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n452), .CK(clk), .RN(n2477), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n451), .CK(clk), .RN(n2477), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n450), .CK(clk), .RN(n2477), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n449), .CK(clk), .RN(n2477), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n448), .CK(clk), .RN(n2477), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n447), .CK(clk), .RN(n2477), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n446), .CK(clk), .RN(n2477), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n445), .CK(clk), .RN(n2477), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n444), .CK(clk), .RN(n2477), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n443), .CK(clk), .RN(n2476), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n442), .CK(clk), .RN(n2476), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n441), .CK(clk), .RN(n2476), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n440), .CK(clk), .RN(n2476), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n439), .CK(clk), .RN(n2476), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n438), .CK(clk), .RN(n2476), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n437), .CK(clk), .RN(n2476), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n436), .CK(clk), .RN(n2476), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n435), .CK(clk), .RN(n2476), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n434), .CK(clk), .RN(n2476), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n433), .CK(clk), .RN(n2476), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n432), .CK(clk), .RN(n2476), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n431), .CK(clk), .RN(n2475), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n430), .CK(clk), .RN(n2475), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n429), .CK(clk), .RN(n2475), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n428), .CK(clk), .RN(n2475), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n331), .CK(clk), .RN(n2467), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n330), .CK(clk), .RN(n2467), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n329), .CK(clk), .RN(n2467), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n328), .CK(clk), .RN(n2467), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n327), .CK(clk), .RN(n2467), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n326), .CK(clk), .RN(n2467), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n325), .CK(clk), .RN(n2467), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n324), .CK(clk), .RN(n2467), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n323), .CK(clk), .RN(n2466), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n322), .CK(clk), .RN(n2466), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n321), .CK(clk), .RN(n2466), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n320), .CK(clk), .RN(n2466), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n319), .CK(clk), .RN(n2466), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n318), .CK(clk), .RN(n2466), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n317), .CK(clk), .RN(n2466), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n316), .CK(clk), .RN(n2466), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n315), .CK(clk), .RN(n2466), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n314), .CK(clk), .RN(n2466), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n313), .CK(clk), .RN(n2466), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n312), .CK(clk), .RN(n2466), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n311), .CK(clk), .RN(n2465), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n310), .CK(clk), .RN(n2465), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n309), .CK(clk), .RN(n2465), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n308), .CK(clk), .RN(n2465), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n307), .CK(clk), .RN(n2465), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n306), .CK(clk), .RN(n2465), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n305), .CK(clk), .RN(n2465), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n304), .CK(clk), .RN(n2465), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n303), .CK(clk), .RN(n2465), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n302), .CK(clk), .RN(n2465), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n301), .CK(clk), .RN(n2465), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n300), .CK(clk), .RN(n2465), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n1035), .CK(clk), .RN(n2526), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n1034), .CK(clk), .RN(n2526), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n1033), .CK(clk), .RN(n2526), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n1032), .CK(clk), .RN(n2526), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n1031), .CK(clk), .RN(n2525), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n1030), .CK(clk), .RN(n2525), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n1029), .CK(clk), .RN(n2525), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n1028), .CK(clk), .RN(n2525), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n1027), .CK(clk), .RN(n2525), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n1026), .CK(clk), .RN(n2525), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n1025), .CK(clk), .RN(n2525), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n1024), .CK(clk), .RN(n2525), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n1023), .CK(clk), .RN(n2525), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n1022), .CK(clk), .RN(n2525), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n1021), .CK(clk), .RN(n2525), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n1020), .CK(clk), .RN(n2525), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n1019), .CK(clk), .RN(n2524), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n1018), .CK(clk), .RN(n2524), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n1017), .CK(clk), .RN(n2524), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n1016), .CK(clk), .RN(n2524), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n1015), .CK(clk), .RN(n2524), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n1014), .CK(clk), .RN(n2524), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n1013), .CK(clk), .RN(n2524), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n1012), .CK(clk), .RN(n2524), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n1011), .CK(clk), .RN(n2524), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n1010), .CK(clk), .RN(n2524), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n1009), .CK(clk), .RN(n2524), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n1008), .CK(clk), .RN(n2524), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n1007), .CK(clk), .RN(n2523), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n1006), .CK(clk), .RN(n2523), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n1005), .CK(clk), .RN(n2523), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n1004), .CK(clk), .RN(n2523), .Q(
        \register[29][0] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n907), .CK(clk), .RN(n2515), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n906), .CK(clk), .RN(n2515), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n905), .CK(clk), .RN(n2515), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n904), .CK(clk), .RN(n2515), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n903), .CK(clk), .RN(n2515), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n902), .CK(clk), .RN(n2515), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n901), .CK(clk), .RN(n2515), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n900), .CK(clk), .RN(n2515), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n899), .CK(clk), .RN(n2514), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n898), .CK(clk), .RN(n2514), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n897), .CK(clk), .RN(n2514), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n896), .CK(clk), .RN(n2514), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n895), .CK(clk), .RN(n2514), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n894), .CK(clk), .RN(n2514), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n893), .CK(clk), .RN(n2514), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n892), .CK(clk), .RN(n2514), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n891), .CK(clk), .RN(n2514), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n890), .CK(clk), .RN(n2514), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n889), .CK(clk), .RN(n2514), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n888), .CK(clk), .RN(n2514), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n887), .CK(clk), .RN(n2513), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n886), .CK(clk), .RN(n2513), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n885), .CK(clk), .RN(n2513), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n884), .CK(clk), .RN(n2513), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n883), .CK(clk), .RN(n2513), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n882), .CK(clk), .RN(n2513), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n881), .CK(clk), .RN(n2513), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n880), .CK(clk), .RN(n2513), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n879), .CK(clk), .RN(n2513), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n878), .CK(clk), .RN(n2513), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n877), .CK(clk), .RN(n2513), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n876), .CK(clk), .RN(n2513), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n779), .CK(clk), .RN(n2504), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n778), .CK(clk), .RN(n2504), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n777), .CK(clk), .RN(n2504), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n776), .CK(clk), .RN(n2504), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n775), .CK(clk), .RN(n2504), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n774), .CK(clk), .RN(n2504), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n773), .CK(clk), .RN(n2504), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n772), .CK(clk), .RN(n2504), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n771), .CK(clk), .RN(n2504), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n770), .CK(clk), .RN(n2504), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n769), .CK(clk), .RN(n2504), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n768), .CK(clk), .RN(n2504), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n767), .CK(clk), .RN(n2503), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n766), .CK(clk), .RN(n2503), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n765), .CK(clk), .RN(n2503), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n764), .CK(clk), .RN(n2503), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n763), .CK(clk), .RN(n2503), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n762), .CK(clk), .RN(n2503), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n761), .CK(clk), .RN(n2503), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n760), .CK(clk), .RN(n2503), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n759), .CK(clk), .RN(n2503), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n758), .CK(clk), .RN(n2503), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n757), .CK(clk), .RN(n2503), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n756), .CK(clk), .RN(n2503), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n755), .CK(clk), .RN(n2502), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n754), .CK(clk), .RN(n2502), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n753), .CK(clk), .RN(n2502), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n752), .CK(clk), .RN(n2502), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n751), .CK(clk), .RN(n2502), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n750), .CK(clk), .RN(n2502), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n749), .CK(clk), .RN(n2502), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n748), .CK(clk), .RN(n2502), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n651), .CK(clk), .RN(n2494), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n650), .CK(clk), .RN(n2494), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n649), .CK(clk), .RN(n2494), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n648), .CK(clk), .RN(n2494), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n647), .CK(clk), .RN(n2493), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n646), .CK(clk), .RN(n2493), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n645), .CK(clk), .RN(n2493), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n644), .CK(clk), .RN(n2493), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n643), .CK(clk), .RN(n2493), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n642), .CK(clk), .RN(n2493), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n641), .CK(clk), .RN(n2493), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n640), .CK(clk), .RN(n2493), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n639), .CK(clk), .RN(n2493), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n638), .CK(clk), .RN(n2493), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n637), .CK(clk), .RN(n2493), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n636), .CK(clk), .RN(n2493), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n635), .CK(clk), .RN(n2492), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n634), .CK(clk), .RN(n2492), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n633), .CK(clk), .RN(n2492), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n632), .CK(clk), .RN(n2492), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n631), .CK(clk), .RN(n2492), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n630), .CK(clk), .RN(n2492), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n629), .CK(clk), .RN(n2492), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n628), .CK(clk), .RN(n2492), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n627), .CK(clk), .RN(n2492), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n626), .CK(clk), .RN(n2492), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n625), .CK(clk), .RN(n2492), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n624), .CK(clk), .RN(n2492), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n623), .CK(clk), .RN(n2491), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n622), .CK(clk), .RN(n2491), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n621), .CK(clk), .RN(n2491), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n620), .CK(clk), .RN(n2491), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n523), .CK(clk), .RN(n2483), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n522), .CK(clk), .RN(n2483), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n521), .CK(clk), .RN(n2483), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n520), .CK(clk), .RN(n2483), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n519), .CK(clk), .RN(n2483), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n518), .CK(clk), .RN(n2483), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n517), .CK(clk), .RN(n2483), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n516), .CK(clk), .RN(n2483), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n515), .CK(clk), .RN(n2482), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n514), .CK(clk), .RN(n2482), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n513), .CK(clk), .RN(n2482), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n512), .CK(clk), .RN(n2482), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n511), .CK(clk), .RN(n2482), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n510), .CK(clk), .RN(n2482), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n509), .CK(clk), .RN(n2482), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n508), .CK(clk), .RN(n2482), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n507), .CK(clk), .RN(n2482), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n506), .CK(clk), .RN(n2482), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n505), .CK(clk), .RN(n2482), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n504), .CK(clk), .RN(n2482), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n503), .CK(clk), .RN(n2481), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n502), .CK(clk), .RN(n2481), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n501), .CK(clk), .RN(n2481), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n500), .CK(clk), .RN(n2481), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n499), .CK(clk), .RN(n2481), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n498), .CK(clk), .RN(n2481), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n497), .CK(clk), .RN(n2481), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n496), .CK(clk), .RN(n2481), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n495), .CK(clk), .RN(n2481), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n494), .CK(clk), .RN(n2481), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n493), .CK(clk), .RN(n2481), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n492), .CK(clk), .RN(n2481), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n395), .CK(clk), .RN(n2472), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n394), .CK(clk), .RN(n2472), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n393), .CK(clk), .RN(n2472), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n392), .CK(clk), .RN(n2472), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n391), .CK(clk), .RN(n2472), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n390), .CK(clk), .RN(n2472), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n389), .CK(clk), .RN(n2472), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n388), .CK(clk), .RN(n2472), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n387), .CK(clk), .RN(n2472), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n386), .CK(clk), .RN(n2472), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n385), .CK(clk), .RN(n2472), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n384), .CK(clk), .RN(n2472), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n383), .CK(clk), .RN(n2471), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n382), .CK(clk), .RN(n2471), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n381), .CK(clk), .RN(n2471), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n380), .CK(clk), .RN(n2471), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n379), .CK(clk), .RN(n2471), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n378), .CK(clk), .RN(n2471), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n377), .CK(clk), .RN(n2471), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n376), .CK(clk), .RN(n2471), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n375), .CK(clk), .RN(n2471), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n374), .CK(clk), .RN(n2471), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n373), .CK(clk), .RN(n2471), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n372), .CK(clk), .RN(n2471), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n371), .CK(clk), .RN(n2470), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n370), .CK(clk), .RN(n2470), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n369), .CK(clk), .RN(n2470), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n368), .CK(clk), .RN(n2470), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n367), .CK(clk), .RN(n2470), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n366), .CK(clk), .RN(n2470), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n365), .CK(clk), .RN(n2470), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n364), .CK(clk), .RN(n2470), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n267), .CK(clk), .RN(n2462), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n266), .CK(clk), .RN(n2462), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n265), .CK(clk), .RN(n2462), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n264), .CK(clk), .RN(n2462), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n263), .CK(clk), .RN(n2461), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n262), .CK(clk), .RN(n2461), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n261), .CK(clk), .RN(n2461), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n260), .CK(clk), .RN(n2461), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n259), .CK(clk), .RN(n2461), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n258), .CK(clk), .RN(n2461), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n257), .CK(clk), .RN(n2461), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n256), .CK(clk), .RN(n2461), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n255), .CK(clk), .RN(n2461), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n254), .CK(clk), .RN(n2461), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n253), .CK(clk), .RN(n2461), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n252), .CK(clk), .RN(n2461), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n251), .CK(clk), .RN(n2460), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n250), .CK(clk), .RN(n2460), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n249), .CK(clk), .RN(n2460), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n248), .CK(clk), .RN(n2460), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n247), .CK(clk), .RN(n2460), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n246), .CK(clk), .RN(n2460), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n245), .CK(clk), .RN(n2460), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n244), .CK(clk), .RN(n2460), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n243), .CK(clk), .RN(n2460), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n242), .CK(clk), .RN(n2460), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n241), .CK(clk), .RN(n2460), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n240), .CK(clk), .RN(n2460), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n239), .CK(clk), .RN(n2459), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n238), .CK(clk), .RN(n2459), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n237), .CK(clk), .RN(n2459), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n236), .CK(clk), .RN(n2459), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n1003), .CK(clk), .RN(n2523), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n1002), .CK(clk), .RN(n2523), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n1001), .CK(clk), .RN(n2523), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n1000), .CK(clk), .RN(n2523), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n999), .CK(clk), .RN(n2523), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n998), .CK(clk), .RN(n2523), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n997), .CK(clk), .RN(n2523), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n996), .CK(clk), .RN(n2523), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n995), .CK(clk), .RN(n2522), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n994), .CK(clk), .RN(n2522), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n993), .CK(clk), .RN(n2522), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n992), .CK(clk), .RN(n2522), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n991), .CK(clk), .RN(n2522), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n990), .CK(clk), .RN(n2522), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n989), .CK(clk), .RN(n2522), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n988), .CK(clk), .RN(n2522), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n987), .CK(clk), .RN(n2522), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n986), .CK(clk), .RN(n2522), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n985), .CK(clk), .RN(n2522), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n984), .CK(clk), .RN(n2522), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n983), .CK(clk), .RN(n2521), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n982), .CK(clk), .RN(n2521), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n981), .CK(clk), .RN(n2521), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n980), .CK(clk), .RN(n2521), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n979), .CK(clk), .RN(n2521), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n978), .CK(clk), .RN(n2521), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n977), .CK(clk), .RN(n2521), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n976), .CK(clk), .RN(n2521), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n975), .CK(clk), .RN(n2521), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n974), .CK(clk), .RN(n2521), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n973), .CK(clk), .RN(n2521), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][0]  ( .D(n972), .CK(clk), .RN(n2521), .Q(
        \register[28][0] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n875), .CK(clk), .RN(n2512), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n874), .CK(clk), .RN(n2512), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n873), .CK(clk), .RN(n2512), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n872), .CK(clk), .RN(n2512), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n871), .CK(clk), .RN(n2512), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n870), .CK(clk), .RN(n2512), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n869), .CK(clk), .RN(n2512), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n868), .CK(clk), .RN(n2512), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n867), .CK(clk), .RN(n2512), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n866), .CK(clk), .RN(n2512), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n865), .CK(clk), .RN(n2512), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n864), .CK(clk), .RN(n2512), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n863), .CK(clk), .RN(n2511), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n862), .CK(clk), .RN(n2511), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n861), .CK(clk), .RN(n2511), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n860), .CK(clk), .RN(n2511), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n859), .CK(clk), .RN(n2511), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n858), .CK(clk), .RN(n2511), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n857), .CK(clk), .RN(n2511), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n856), .CK(clk), .RN(n2511), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n855), .CK(clk), .RN(n2511), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n854), .CK(clk), .RN(n2511), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n853), .CK(clk), .RN(n2511), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n852), .CK(clk), .RN(n2511), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n851), .CK(clk), .RN(n2510), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n850), .CK(clk), .RN(n2510), .Q(
        \register[24][6] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n849), .CK(clk), .RN(n2510), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n848), .CK(clk), .RN(n2510), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n847), .CK(clk), .RN(n2510), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n846), .CK(clk), .RN(n2510), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n845), .CK(clk), .RN(n2510), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n844), .CK(clk), .RN(n2510), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n747), .CK(clk), .RN(n2502), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n746), .CK(clk), .RN(n2502), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n745), .CK(clk), .RN(n2502), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n744), .CK(clk), .RN(n2502), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n743), .CK(clk), .RN(n2501), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n742), .CK(clk), .RN(n2501), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n741), .CK(clk), .RN(n2501), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n740), .CK(clk), .RN(n2501), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n739), .CK(clk), .RN(n2501), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n738), .CK(clk), .RN(n2501), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n737), .CK(clk), .RN(n2501), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n736), .CK(clk), .RN(n2501), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n735), .CK(clk), .RN(n2501), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n734), .CK(clk), .RN(n2501), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n733), .CK(clk), .RN(n2501), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n732), .CK(clk), .RN(n2501), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n731), .CK(clk), .RN(n2500), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n730), .CK(clk), .RN(n2500), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n729), .CK(clk), .RN(n2500), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n728), .CK(clk), .RN(n2500), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n727), .CK(clk), .RN(n2500), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n726), .CK(clk), .RN(n2500), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n725), .CK(clk), .RN(n2500), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n724), .CK(clk), .RN(n2500), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n723), .CK(clk), .RN(n2500), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n722), .CK(clk), .RN(n2500), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n721), .CK(clk), .RN(n2500), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n720), .CK(clk), .RN(n2500), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n719), .CK(clk), .RN(n2499), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n718), .CK(clk), .RN(n2499), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n717), .CK(clk), .RN(n2499), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[20][0]  ( .D(n716), .CK(clk), .RN(n2499), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n619), .CK(clk), .RN(n2491), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n618), .CK(clk), .RN(n2491), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n617), .CK(clk), .RN(n2491), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n616), .CK(clk), .RN(n2491), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n615), .CK(clk), .RN(n2491), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n614), .CK(clk), .RN(n2491), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n613), .CK(clk), .RN(n2491), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n612), .CK(clk), .RN(n2491), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n611), .CK(clk), .RN(n2490), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n610), .CK(clk), .RN(n2490), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n609), .CK(clk), .RN(n2490), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n608), .CK(clk), .RN(n2490), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n607), .CK(clk), .RN(n2490), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n606), .CK(clk), .RN(n2490), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n605), .CK(clk), .RN(n2490), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n604), .CK(clk), .RN(n2490), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n603), .CK(clk), .RN(n2490), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n602), .CK(clk), .RN(n2490), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n601), .CK(clk), .RN(n2490), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n600), .CK(clk), .RN(n2490), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n599), .CK(clk), .RN(n2489), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n598), .CK(clk), .RN(n2489), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n597), .CK(clk), .RN(n2489), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n596), .CK(clk), .RN(n2489), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n595), .CK(clk), .RN(n2489), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n594), .CK(clk), .RN(n2489), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n593), .CK(clk), .RN(n2489), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n592), .CK(clk), .RN(n2489), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n591), .CK(clk), .RN(n2489), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n590), .CK(clk), .RN(n2489), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n589), .CK(clk), .RN(n2489), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n588), .CK(clk), .RN(n2489), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n491), .CK(clk), .RN(n2480), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n490), .CK(clk), .RN(n2480), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n489), .CK(clk), .RN(n2480), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n488), .CK(clk), .RN(n2480), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n487), .CK(clk), .RN(n2480), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n486), .CK(clk), .RN(n2480), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n485), .CK(clk), .RN(n2480), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n484), .CK(clk), .RN(n2480), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n483), .CK(clk), .RN(n2480), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n482), .CK(clk), .RN(n2480), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n481), .CK(clk), .RN(n2480), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n480), .CK(clk), .RN(n2480), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n479), .CK(clk), .RN(n2479), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n478), .CK(clk), .RN(n2479), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n477), .CK(clk), .RN(n2479), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n476), .CK(clk), .RN(n2479), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n475), .CK(clk), .RN(n2479), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n474), .CK(clk), .RN(n2479), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n473), .CK(clk), .RN(n2479), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n472), .CK(clk), .RN(n2479), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n471), .CK(clk), .RN(n2479), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n470), .CK(clk), .RN(n2479), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n469), .CK(clk), .RN(n2479), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n468), .CK(clk), .RN(n2479), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n467), .CK(clk), .RN(n2478), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n466), .CK(clk), .RN(n2478), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n465), .CK(clk), .RN(n2478), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n464), .CK(clk), .RN(n2478), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n463), .CK(clk), .RN(n2478), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n462), .CK(clk), .RN(n2478), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n461), .CK(clk), .RN(n2478), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n460), .CK(clk), .RN(n2478), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n363), .CK(clk), .RN(n2470), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n362), .CK(clk), .RN(n2470), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n361), .CK(clk), .RN(n2470), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n360), .CK(clk), .RN(n2470), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n359), .CK(clk), .RN(n2469), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n358), .CK(clk), .RN(n2469), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n357), .CK(clk), .RN(n2469), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n356), .CK(clk), .RN(n2469), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n355), .CK(clk), .RN(n2469), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n354), .CK(clk), .RN(n2469), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n353), .CK(clk), .RN(n2469), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n352), .CK(clk), .RN(n2469), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n351), .CK(clk), .RN(n2469), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n350), .CK(clk), .RN(n2469), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n349), .CK(clk), .RN(n2469), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n348), .CK(clk), .RN(n2469), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n347), .CK(clk), .RN(n2468), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n346), .CK(clk), .RN(n2468), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n345), .CK(clk), .RN(n2468), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n344), .CK(clk), .RN(n2468), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n343), .CK(clk), .RN(n2468), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n342), .CK(clk), .RN(n2468), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n341), .CK(clk), .RN(n2468), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n340), .CK(clk), .RN(n2468), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n339), .CK(clk), .RN(n2468), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n338), .CK(clk), .RN(n2468), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n337), .CK(clk), .RN(n2468), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n336), .CK(clk), .RN(n2468), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n335), .CK(clk), .RN(n2467), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n334), .CK(clk), .RN(n2467), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n333), .CK(clk), .RN(n2467), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n332), .CK(clk), .RN(n2467), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n235), .CK(clk), .RN(n2459), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n234), .CK(clk), .RN(n2459), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n233), .CK(clk), .RN(n2459), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n232), .CK(clk), .RN(n2459), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n231), .CK(clk), .RN(n2459), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n230), .CK(clk), .RN(n2459), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n229), .CK(clk), .RN(n2459), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n228), .CK(clk), .RN(n2459), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n227), .CK(clk), .RN(n2458), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n226), .CK(clk), .RN(n2458), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n225), .CK(clk), .RN(n2458), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n224), .CK(clk), .RN(n2458), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n223), .CK(clk), .RN(n2458), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n222), .CK(clk), .RN(n2458), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n221), .CK(clk), .RN(n2458), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n220), .CK(clk), .RN(n2458), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n219), .CK(clk), .RN(n2458), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n218), .CK(clk), .RN(n2458), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n217), .CK(clk), .RN(n2458), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n216), .CK(clk), .RN(n2458), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n215), .CK(clk), .RN(n2457), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n214), .CK(clk), .RN(n2457), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n213), .CK(clk), .RN(n2457), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n212), .CK(clk), .RN(n2457), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n211), .CK(clk), .RN(n2457), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n210), .CK(clk), .RN(n2457), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n209), .CK(clk), .RN(n2457), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n208), .CK(clk), .RN(n2457), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n207), .CK(clk), .RN(n2457), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n206), .CK(clk), .RN(n2457), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n205), .CK(clk), .RN(n2457), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n204), .CK(clk), .RN(n2457), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n1067), .CK(clk), .RN(n2528), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n1066), .CK(clk), .RN(n2528), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n1065), .CK(clk), .RN(n2528), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n1064), .CK(clk), .RN(n2528), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n1063), .CK(clk), .RN(n2528), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n1062), .CK(clk), .RN(n2528), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n1061), .CK(clk), .RN(n2528), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n1060), .CK(clk), .RN(n2528), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n1059), .CK(clk), .RN(n2528), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n1058), .CK(clk), .RN(n2528), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n1057), .CK(clk), .RN(n2528), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n1056), .CK(clk), .RN(n2528), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n1055), .CK(clk), .RN(n2527), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n1054), .CK(clk), .RN(n2527), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n1053), .CK(clk), .RN(n2527), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n1052), .CK(clk), .RN(n2527), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n1051), .CK(clk), .RN(n2527), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n1050), .CK(clk), .RN(n2527), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n1049), .CK(clk), .RN(n2527), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n1048), .CK(clk), .RN(n2527), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n1047), .CK(clk), .RN(n2527), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n1046), .CK(clk), .RN(n2527), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n1045), .CK(clk), .RN(n2527), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n1044), .CK(clk), .RN(n2527), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n1043), .CK(clk), .RN(n2526), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n1042), .CK(clk), .RN(n2526), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n1041), .CK(clk), .RN(n2526), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n1040), .CK(clk), .RN(n2526), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n1039), .CK(clk), .RN(n2526), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n1038), .CK(clk), .RN(n2526), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n1037), .CK(clk), .RN(n2526), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][0]  ( .D(n1036), .CK(clk), .RN(n2526), .Q(
        \register[30][0] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n939), .CK(clk), .RN(n2518), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n938), .CK(clk), .RN(n2518), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n937), .CK(clk), .RN(n2518), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n936), .CK(clk), .RN(n2518), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n935), .CK(clk), .RN(n2517), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n934), .CK(clk), .RN(n2517), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n933), .CK(clk), .RN(n2517), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n932), .CK(clk), .RN(n2517), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n931), .CK(clk), .RN(n2517), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n930), .CK(clk), .RN(n2517), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n929), .CK(clk), .RN(n2517), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n928), .CK(clk), .RN(n2517), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n927), .CK(clk), .RN(n2517), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n926), .CK(clk), .RN(n2517), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n925), .CK(clk), .RN(n2517), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n924), .CK(clk), .RN(n2517), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n923), .CK(clk), .RN(n2516), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n922), .CK(clk), .RN(n2516), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n921), .CK(clk), .RN(n2516), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n920), .CK(clk), .RN(n2516), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n919), .CK(clk), .RN(n2516), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n918), .CK(clk), .RN(n2516), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n917), .CK(clk), .RN(n2516), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n916), .CK(clk), .RN(n2516), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n915), .CK(clk), .RN(n2516), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n914), .CK(clk), .RN(n2516), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n913), .CK(clk), .RN(n2516), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n912), .CK(clk), .RN(n2516), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n911), .CK(clk), .RN(n2515), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n910), .CK(clk), .RN(n2515), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n909), .CK(clk), .RN(n2515), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n908), .CK(clk), .RN(n2515), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n811), .CK(clk), .RN(n2507), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n810), .CK(clk), .RN(n2507), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n809), .CK(clk), .RN(n2507), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n808), .CK(clk), .RN(n2507), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n807), .CK(clk), .RN(n2507), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n806), .CK(clk), .RN(n2507), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n805), .CK(clk), .RN(n2507), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n804), .CK(clk), .RN(n2507), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n803), .CK(clk), .RN(n2506), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n802), .CK(clk), .RN(n2506), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n801), .CK(clk), .RN(n2506), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n800), .CK(clk), .RN(n2506), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n799), .CK(clk), .RN(n2506), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n798), .CK(clk), .RN(n2506), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n797), .CK(clk), .RN(n2506), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n796), .CK(clk), .RN(n2506), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n795), .CK(clk), .RN(n2506), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n794), .CK(clk), .RN(n2506), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n793), .CK(clk), .RN(n2506), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n792), .CK(clk), .RN(n2506), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n791), .CK(clk), .RN(n2505), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n790), .CK(clk), .RN(n2505), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n789), .CK(clk), .RN(n2505), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n788), .CK(clk), .RN(n2505), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n787), .CK(clk), .RN(n2505), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n786), .CK(clk), .RN(n2505), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n785), .CK(clk), .RN(n2505), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n784), .CK(clk), .RN(n2505), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n783), .CK(clk), .RN(n2505), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n782), .CK(clk), .RN(n2505), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n781), .CK(clk), .RN(n2505), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n780), .CK(clk), .RN(n2505), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n683), .CK(clk), .RN(n2496), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n682), .CK(clk), .RN(n2496), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n681), .CK(clk), .RN(n2496), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n680), .CK(clk), .RN(n2496), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n679), .CK(clk), .RN(n2496), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n678), .CK(clk), .RN(n2496), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n677), .CK(clk), .RN(n2496), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n676), .CK(clk), .RN(n2496), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n675), .CK(clk), .RN(n2496), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n674), .CK(clk), .RN(n2496), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n673), .CK(clk), .RN(n2496), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n672), .CK(clk), .RN(n2496), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n671), .CK(clk), .RN(n2495), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n670), .CK(clk), .RN(n2495), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n669), .CK(clk), .RN(n2495), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n668), .CK(clk), .RN(n2495), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n667), .CK(clk), .RN(n2495), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n666), .CK(clk), .RN(n2495), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n665), .CK(clk), .RN(n2495), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n664), .CK(clk), .RN(n2495), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n663), .CK(clk), .RN(n2495), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n662), .CK(clk), .RN(n2495), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n661), .CK(clk), .RN(n2495), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n660), .CK(clk), .RN(n2495), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n659), .CK(clk), .RN(n2494), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n658), .CK(clk), .RN(n2494), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n657), .CK(clk), .RN(n2494), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n656), .CK(clk), .RN(n2494), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n655), .CK(clk), .RN(n2494), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n654), .CK(clk), .RN(n2494), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n653), .CK(clk), .RN(n2494), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n652), .CK(clk), .RN(n2494), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n555), .CK(clk), .RN(n2486), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n554), .CK(clk), .RN(n2486), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n553), .CK(clk), .RN(n2486), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n552), .CK(clk), .RN(n2486), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n551), .CK(clk), .RN(n2485), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n550), .CK(clk), .RN(n2485), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n549), .CK(clk), .RN(n2485), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n548), .CK(clk), .RN(n2485), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n547), .CK(clk), .RN(n2485), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n546), .CK(clk), .RN(n2485), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n545), .CK(clk), .RN(n2485), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n544), .CK(clk), .RN(n2485), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n543), .CK(clk), .RN(n2485), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n542), .CK(clk), .RN(n2485), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n541), .CK(clk), .RN(n2485), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n540), .CK(clk), .RN(n2485), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n539), .CK(clk), .RN(n2484), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n538), .CK(clk), .RN(n2484), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n537), .CK(clk), .RN(n2484), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n536), .CK(clk), .RN(n2484), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n535), .CK(clk), .RN(n2484), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n534), .CK(clk), .RN(n2484), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n533), .CK(clk), .RN(n2484), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n532), .CK(clk), .RN(n2484), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n531), .CK(clk), .RN(n2484), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n530), .CK(clk), .RN(n2484), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n529), .CK(clk), .RN(n2484), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n528), .CK(clk), .RN(n2484), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n527), .CK(clk), .RN(n2483), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n526), .CK(clk), .RN(n2483), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n525), .CK(clk), .RN(n2483), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n524), .CK(clk), .RN(n2483), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n427), .CK(clk), .RN(n2475), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n426), .CK(clk), .RN(n2475), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n425), .CK(clk), .RN(n2475), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n424), .CK(clk), .RN(n2475), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n423), .CK(clk), .RN(n2475), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n422), .CK(clk), .RN(n2475), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n421), .CK(clk), .RN(n2475), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n420), .CK(clk), .RN(n2475), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n419), .CK(clk), .RN(n2474), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n418), .CK(clk), .RN(n2474), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n417), .CK(clk), .RN(n2474), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n416), .CK(clk), .RN(n2474), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n415), .CK(clk), .RN(n2474), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n414), .CK(clk), .RN(n2474), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n413), .CK(clk), .RN(n2474), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n412), .CK(clk), .RN(n2474), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n411), .CK(clk), .RN(n2474), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n410), .CK(clk), .RN(n2474), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n409), .CK(clk), .RN(n2474), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n408), .CK(clk), .RN(n2474), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n407), .CK(clk), .RN(n2473), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n406), .CK(clk), .RN(n2473), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n405), .CK(clk), .RN(n2473), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n404), .CK(clk), .RN(n2473), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n403), .CK(clk), .RN(n2473), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n402), .CK(clk), .RN(n2473), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n401), .CK(clk), .RN(n2473), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n400), .CK(clk), .RN(n2473), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n399), .CK(clk), .RN(n2473), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n398), .CK(clk), .RN(n2473), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n397), .CK(clk), .RN(n2473), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n396), .CK(clk), .RN(n2473), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n299), .CK(clk), .RN(n2464), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n298), .CK(clk), .RN(n2464), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n297), .CK(clk), .RN(n2464), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n296), .CK(clk), .RN(n2464), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n295), .CK(clk), .RN(n2464), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n294), .CK(clk), .RN(n2464), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n293), .CK(clk), .RN(n2464), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n292), .CK(clk), .RN(n2464), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n291), .CK(clk), .RN(n2464), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n290), .CK(clk), .RN(n2464), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n289), .CK(clk), .RN(n2464), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n288), .CK(clk), .RN(n2464), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n287), .CK(clk), .RN(n2463), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n286), .CK(clk), .RN(n2463), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n285), .CK(clk), .RN(n2463), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n284), .CK(clk), .RN(n2463), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n283), .CK(clk), .RN(n2463), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n282), .CK(clk), .RN(n2463), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n281), .CK(clk), .RN(n2463), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n280), .CK(clk), .RN(n2463), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n279), .CK(clk), .RN(n2463), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n278), .CK(clk), .RN(n2463), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n277), .CK(clk), .RN(n2463), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n276), .CK(clk), .RN(n2463), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n275), .CK(clk), .RN(n2462), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n274), .CK(clk), .RN(n2462), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n273), .CK(clk), .RN(n2462), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n272), .CK(clk), .RN(n2462), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n271), .CK(clk), .RN(n2462), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n270), .CK(clk), .RN(n2462), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n269), .CK(clk), .RN(n2462), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n268), .CK(clk), .RN(n2462), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[3][31]  ( .D(n203), .CK(clk), .RN(n2456), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n202), .CK(clk), .RN(n2456), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n201), .CK(clk), .RN(n2456), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n200), .CK(clk), .RN(n2456), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n199), .CK(clk), .RN(n2456), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n198), .CK(clk), .RN(n2456), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n197), .CK(clk), .RN(n2456), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n196), .CK(clk), .RN(n2456), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n195), .CK(clk), .RN(n2456), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n194), .CK(clk), .RN(n2456), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n193), .CK(clk), .RN(n2456), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n192), .CK(clk), .RN(n2456), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n191), .CK(clk), .RN(n2455), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n190), .CK(clk), .RN(n2455), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n189), .CK(clk), .RN(n2455), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n188), .CK(clk), .RN(n2455), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n187), .CK(clk), .RN(n2455), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n186), .CK(clk), .RN(n2455), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n185), .CK(clk), .RN(n2455), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n184), .CK(clk), .RN(n2455), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n183), .CK(clk), .RN(n2455), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n182), .CK(clk), .RN(n2455), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n181), .CK(clk), .RN(n2455), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n180), .CK(clk), .RN(n2455), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n179), .CK(clk), .RN(n2454), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n178), .CK(clk), .RN(n2454), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n177), .CK(clk), .RN(n2454), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n176), .CK(clk), .RN(n2454), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n175), .CK(clk), .RN(n2454), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n174), .CK(clk), .RN(n2454), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n173), .CK(clk), .RN(n2454), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n172), .CK(clk), .RN(n2454), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n139), .CK(clk), .RN(n2451), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n138), .CK(clk), .RN(n2451), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n137), .CK(clk), .RN(n2451), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n136), .CK(clk), .RN(n2451), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n135), .CK(clk), .RN(n2451), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n134), .CK(clk), .RN(n2451), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n133), .CK(clk), .RN(n2451), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n132), .CK(clk), .RN(n2451), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n131), .CK(clk), .RN(n2450), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n130), .CK(clk), .RN(n2450), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n129), .CK(clk), .RN(n2450), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n128), .CK(clk), .RN(n2450), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n127), .CK(clk), .RN(n2450), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n126), .CK(clk), .RN(n2450), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n125), .CK(clk), .RN(n2450), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n124), .CK(clk), .RN(n2450), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n123), .CK(clk), .RN(n2450), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n122), .CK(clk), .RN(n2450), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n121), .CK(clk), .RN(n2450), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n120), .CK(clk), .RN(n2450), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n119), .CK(clk), .RN(n2449), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n118), .CK(clk), .RN(n2449), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n117), .CK(clk), .RN(n2449), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n116), .CK(clk), .RN(n2449), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n115), .CK(clk), .RN(n2449), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n114), .CK(clk), .RN(n2449), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n113), .CK(clk), .RN(n2449), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n112), .CK(clk), .RN(n2449), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n111), .CK(clk), .RN(n2449), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n110), .CK(clk), .RN(n2449), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][1]  ( .D(n109), .CK(clk), .RN(n2449), .Q(
        \register[1][1] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n108), .CK(clk), .RN(n2449), .Q(
        \register[1][0] ) );
  INVX4 U3 ( .A(wdata[7]), .Y(n2610) );
  CLKINVX4 U4 ( .A(n4), .Y(n11) );
  INVX4 U5 ( .A(wsel[1]), .Y(n10) );
  INVX4 U6 ( .A(wsel[2]), .Y(n2619) );
  INVX4 U7 ( .A(wsel[0]), .Y(n2620) );
  BUFX4 U8 ( .A(n2114), .Y(n2124) );
  OAI2BB2XL U9 ( .B0(n2240), .B1(n2430), .A0N(N53), .A1N(n2433), .Y(rdata1[3])
         );
  OAI2BB2XL U10 ( .B0(n2238), .B1(n2430), .A0N(N52), .A1N(n2433), .Y(rdata1[4]) );
  OAI2BB2XL U11 ( .B0(n2193), .B1(n2431), .A0N(N37), .A1N(n2432), .Y(
        rdata1[19]) );
  OAI2BB2XL U12 ( .B0(n2175), .B1(n2431), .A0N(N31), .A1N(n2433), .Y(
        rdata1[25]) );
  OAI2BB2XL U13 ( .B0(n2172), .B1(n2431), .A0N(N30), .A1N(n2433), .Y(
        rdata1[26]) );
  OAI2BB2XL U14 ( .B0(n2169), .B1(n2430), .A0N(N29), .A1N(n2433), .Y(
        rdata1[27]) );
  OAI2BB2XL U15 ( .B0(n2163), .B1(n2430), .A0N(N27), .A1N(n2433), .Y(
        rdata1[29]) );
  OAI2BB2XL U16 ( .B0(n2160), .B1(n2430), .A0N(N26), .A1N(n2433), .Y(
        rdata1[30]) );
  OAI2BB2XL U17 ( .B0(n2157), .B1(n2430), .A0N(N25), .A1N(n2433), .Y(
        rdata1[31]) );
  OAI2BB2XL U18 ( .B0(n2243), .B1(n2430), .A0N(N54), .A1N(n2433), .Y(rdata1[2]) );
  OAI2BB2XL U19 ( .B0(n2166), .B1(n2430), .A0N(N28), .A1N(n2433), .Y(
        rdata1[28]) );
  CLKBUFX3 U20 ( .A(N12), .Y(n2443) );
  BUFX2 U21 ( .A(n2135), .Y(n2138) );
  BUFX2 U22 ( .A(n1590), .Y(n1594) );
  CLKBUFX3 U23 ( .A(N13), .Y(n1589) );
  BUFX4 U24 ( .A(n1569), .Y(n1583) );
  BUFX2 U25 ( .A(n90), .Y(n2338) );
  NAND2X1 U26 ( .A(n100), .B(n11), .Y(n105) );
  CLKBUFX3 U27 ( .A(n1589), .Y(n1567) );
  BUFX4 U28 ( .A(n2136), .Y(n2151) );
  BUFX2 U29 ( .A(n2343), .Y(n2342) );
  BUFX4 U30 ( .A(n2343), .Y(n2346) );
  BUFX2 U31 ( .A(n2389), .Y(n2390) );
  OR3XL U32 ( .A(wsel[1]), .B(wsel[2]), .C(n2620), .Y(n1) );
  OR3XL U33 ( .A(wsel[0]), .B(wsel[1]), .C(n2619), .Y(n2) );
  CLKBUFX3 U34 ( .A(n87), .Y(n2353) );
  CLKBUFX3 U35 ( .A(n96), .Y(n2309) );
  CLKBUFX3 U36 ( .A(n74), .Y(n2398) );
  OR3XL U37 ( .A(wsel[1]), .B(wsel[2]), .C(wsel[0]), .Y(n3) );
  BUFX2 U38 ( .A(n1567), .Y(n1572) );
  CLKBUFX3 U39 ( .A(n2441), .Y(n2099) );
  OR3XL U40 ( .A(n2620), .B(wsel[1]), .C(n2619), .Y(n4) );
  CLKBUFX3 U41 ( .A(n1566), .Y(n1560) );
  NAND2X1 U42 ( .A(n91), .B(n9), .Y(n92) );
  NAND2X1 U43 ( .A(n100), .B(n9), .Y(n101) );
  BUFX2 U44 ( .A(n88), .Y(n2347) );
  BUFX2 U45 ( .A(n78), .Y(n2389) );
  BUFX2 U46 ( .A(N17), .Y(n2439) );
  INVX1 U47 ( .A(wdata[3]), .Y(n2614) );
  BUFX2 U48 ( .A(n2446), .Y(n1549) );
  BUFX4 U49 ( .A(n70), .Y(n2411) );
  BUFX2 U50 ( .A(n2442), .Y(n2093) );
  BUFX2 U51 ( .A(n2106), .Y(n2100) );
  BUFX2 U52 ( .A(n86), .Y(n2359) );
  BUFX2 U53 ( .A(n95), .Y(n2315) );
  BUFX2 U54 ( .A(n72), .Y(n2404) );
  BUFX2 U55 ( .A(n97), .Y(n2303) );
  BUFX4 U56 ( .A(n56), .Y(n2429) );
  BUFX4 U57 ( .A(n84), .Y(n2371) );
  BUFX4 U58 ( .A(n85), .Y(n2365) );
  BUFX4 U59 ( .A(n93), .Y(n2327) );
  BUFX4 U60 ( .A(n94), .Y(n2321) );
  BUFX4 U61 ( .A(n102), .Y(n2279) );
  BUFX4 U62 ( .A(n103), .Y(n2273) );
  BUFX4 U63 ( .A(n83), .Y(n2377) );
  BUFX4 U64 ( .A(n68), .Y(n2418) );
  BUFX4 U65 ( .A(n65), .Y(n2424) );
  BUFX2 U66 ( .A(n47), .Y(n2434) );
  CLKBUFX4 U67 ( .A(n2140), .Y(n2141) );
  MXI4X1 U68 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n2145), .S1(n2118), .Y(
        n1840) );
  MXI4X1 U69 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n2145), .S1(n2118), 
        .Y(n1838) );
  MXI4X1 U70 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n2145), .S1(n2118), 
        .Y(n1836) );
  MXI4X1 U71 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n2145), .S1(n2118), 
        .Y(n1837) );
  MXI4X1 U72 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n2145), .S1(n2118), 
        .Y(n1839) );
  CLKBUFX4 U73 ( .A(n2108), .Y(n2127) );
  BUFX20 U74 ( .A(n2136), .Y(n2145) );
  BUFX20 U75 ( .A(n2443), .Y(n1599) );
  INVX6 U76 ( .A(wsel[4]), .Y(n14) );
  NOR3XL U77 ( .A(wsel[3]), .B(wsel[4]), .C(n2621), .Y(n67) );
  NOR3XL U78 ( .A(n2618), .B(wsel[4]), .C(n2621), .Y(n81) );
  CLKINVX4 U79 ( .A(n3), .Y(n5) );
  INVX3 U80 ( .A(n67), .Y(n6) );
  CLKINVX8 U81 ( .A(n6), .Y(n7) );
  CLKINVX4 U82 ( .A(n2), .Y(n8) );
  NOR3X4 U83 ( .A(wsel[0]), .B(wsel[2]), .C(n10), .Y(n69) );
  CLKINVX4 U84 ( .A(n1), .Y(n9) );
  NOR3X6 U85 ( .A(n10), .B(n2620), .C(n2619), .Y(n79) );
  NOR3X2 U86 ( .A(n10), .B(wsel[0]), .C(n2619), .Y(n77) );
  NOR3X1 U87 ( .A(n2620), .B(wsel[2]), .C(n10), .Y(n71) );
  INVX2 U88 ( .A(n77), .Y(n12) );
  CLKINVX6 U89 ( .A(n12), .Y(n13) );
  INVX3 U90 ( .A(n81), .Y(n15) );
  CLKINVX8 U91 ( .A(n15), .Y(n16) );
  INVX8 U92 ( .A(wen), .Y(n2621) );
  INVX2 U93 ( .A(wsel[3]), .Y(n2618) );
  NAND2XL U94 ( .A(n69), .B(n7), .Y(n68) );
  NAND2XL U95 ( .A(n71), .B(n7), .Y(n70) );
  NAND2XL U96 ( .A(n100), .B(n13), .Y(n106) );
  NAND2XL U97 ( .A(n8), .B(n7), .Y(n72) );
  NAND2XL U98 ( .A(n100), .B(n8), .Y(n104) );
  NAND2XL U99 ( .A(n91), .B(n8), .Y(n95) );
  NAND2XL U100 ( .A(n16), .B(n8), .Y(n86) );
  NAND2XL U101 ( .A(n9), .B(n7), .Y(n65) );
  BUFX2 U102 ( .A(n2111), .Y(n2131) );
  CLKBUFX4 U103 ( .A(n2251), .Y(n2255) );
  BUFX2 U104 ( .A(n2439), .Y(n2140) );
  BUFX8 U105 ( .A(n2099), .Y(n2094) );
  BUFX8 U106 ( .A(n1551), .Y(n1553) );
  BUFX6 U107 ( .A(n2100), .Y(n2101) );
  CLKBUFX2 U108 ( .A(n1551), .Y(n1552) );
  CLKBUFX4 U109 ( .A(n2297), .Y(n2301) );
  MXI4XL U110 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1606), .S1(n1582), 
        .Y(n1246) );
  MXI4XL U111 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1599), .S1(n1578), .Y(
        n1138) );
  MXI4XL U112 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1600), .S1(n1578), .Y(
        n1142) );
  MXI4XL U113 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1606), .S1(n1582), 
        .Y(n1244) );
  MXI4XL U114 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1600), .S1(n1578), .Y(
        n1140) );
  MXI4XL U115 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n2148), .S1(n2124), .Y(
        n1730) );
  MXI4XL U116 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n2149), .S1(n2124), .Y(
        n1736) );
  BUFX3 U117 ( .A(n1593), .Y(n1606) );
  XNOR2X1 U118 ( .A(n14), .B(n2446), .Y(n62) );
  XNOR2X1 U119 ( .A(n2618), .B(n2445), .Y(n63) );
  MXI2X1 U120 ( .A(n2555), .B(n1536), .S0(n1606), .Y(n1539) );
  BUFX2 U121 ( .A(n1569), .Y(n1587) );
  NOR2X1 U122 ( .A(n2131), .B(\register[1][20] ), .Y(n1987) );
  MXI2X1 U123 ( .A(n2574), .B(n1985), .S0(n2153), .Y(n1988) );
  OR2XL U124 ( .A(n2443), .B(N13), .Y(n64) );
  BUFX4 U125 ( .A(n2445), .Y(n1558) );
  INVXL U126 ( .A(wdata[24]), .Y(n2593) );
  OAI2BB2X1 U127 ( .B0(n2196), .B1(n2431), .A0N(N38), .A1N(n2433), .Y(
        rdata1[18]) );
  OAI2BB2X1 U128 ( .B0(n2178), .B1(n2431), .A0N(N32), .A1N(n2432), .Y(
        rdata1[24]) );
  MXI2X1 U129 ( .A(n2561), .B(n2050), .S0(n2152), .Y(n2053) );
  MXI2X1 U130 ( .A(n2568), .B(n1471), .S0(n1607), .Y(n1474) );
  NOR2BX1 U131 ( .AN(n2127), .B(\register[3][20] ), .Y(n1985) );
  NOR2BX1 U132 ( .AN(n2127), .B(\register[3][7] ), .Y(n2050) );
  NOR2BX1 U133 ( .AN(n1583), .B(\register[3][14] ), .Y(n1471) );
  MXI4X1 U134 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1605), .S1(n1582), 
        .Y(n1242) );
  CLKBUFX3 U135 ( .A(n2136), .Y(n2154) );
  CLKBUFX3 U136 ( .A(n1592), .Y(n1609) );
  BUFX4 U137 ( .A(n1560), .Y(n1561) );
  BUFX4 U138 ( .A(n107), .Y(n2251) );
  NAND2XL U139 ( .A(n100), .B(n79), .Y(n107) );
  BUFX8 U140 ( .A(N18), .Y(n2134) );
  BUFX4 U141 ( .A(n101), .Y(n2284) );
  BUFX4 U142 ( .A(n2411), .Y(n2409) );
  CLKBUFX2 U143 ( .A(n92), .Y(n2332) );
  BUFX2 U144 ( .A(n1549), .Y(n1546) );
  CLKBUFX2 U145 ( .A(n2424), .Y(n2423) );
  BUFX2 U146 ( .A(n2410), .Y(n2416) );
  CLKBUFX2 U147 ( .A(n2411), .Y(n2410) );
  CLKBUFX2 U148 ( .A(n2418), .Y(n2417) );
  CLKBUFX2 U149 ( .A(n2440), .Y(n2106) );
  CLKBUFX2 U150 ( .A(n2444), .Y(n1566) );
  BUFX4 U151 ( .A(n104), .Y(n2266) );
  BUFX4 U152 ( .A(n106), .Y(n2256) );
  BUFX4 U153 ( .A(n90), .Y(n2337) );
  CLKBUFX2 U154 ( .A(n104), .Y(n2267) );
  CLKBUFX2 U155 ( .A(n106), .Y(n2257) );
  CLKBUFX2 U156 ( .A(n2353), .Y(n2352) );
  CLKBUFX2 U157 ( .A(n2309), .Y(n2308) );
  CLKBUFX2 U158 ( .A(n2398), .Y(n2397) );
  CLKBUFX2 U159 ( .A(n2404), .Y(n2403) );
  CLKBUFX2 U160 ( .A(n2359), .Y(n2358) );
  CLKBUFX2 U161 ( .A(n2315), .Y(n2314) );
  CLKBUFX2 U162 ( .A(n2303), .Y(n2302) );
  CLKBUFX2 U163 ( .A(n2291), .Y(n2290) );
  CLKBUFX2 U164 ( .A(n2383), .Y(n2382) );
  CLKBUFX2 U165 ( .A(n2377), .Y(n2376) );
  CLKBUFX2 U166 ( .A(n2365), .Y(n2364) );
  CLKBUFX2 U167 ( .A(n2321), .Y(n2320) );
  CLKBUFX2 U168 ( .A(n2371), .Y(n2370) );
  CLKBUFX2 U169 ( .A(n2327), .Y(n2326) );
  CLKBUFX2 U170 ( .A(n101), .Y(n2285) );
  CLKBUFX2 U171 ( .A(n2273), .Y(n2272) );
  CLKBUFX2 U172 ( .A(n2279), .Y(n2278) );
  CLKBUFX2 U173 ( .A(rst_n), .Y(n2448) );
  CLKBUFX2 U174 ( .A(rst_n), .Y(n2447) );
  BUFX4 U175 ( .A(n89), .Y(n2343) );
  NAND2XL U176 ( .A(n16), .B(n79), .Y(n89) );
  BUFX4 U177 ( .A(n98), .Y(n2297) );
  NAND2XL U178 ( .A(n91), .B(n79), .Y(n98) );
  CLKBUFX2 U179 ( .A(N21), .Y(n2442) );
  NAND2XL U180 ( .A(n100), .B(n71), .Y(n103) );
  NAND2XL U181 ( .A(n100), .B(n69), .Y(n102) );
  INVXL U182 ( .A(wdata[12]), .Y(n2605) );
  INVXL U183 ( .A(wdata[14]), .Y(n2603) );
  INVXL U184 ( .A(wdata[22]), .Y(n2595) );
  INVXL U185 ( .A(wdata[25]), .Y(n2592) );
  INVXL U186 ( .A(wdata[27]), .Y(n2590) );
  INVXL U187 ( .A(wdata[31]), .Y(n2586) );
  INVXL U188 ( .A(wdata[1]), .Y(n2616) );
  INVXL U189 ( .A(wdata[5]), .Y(n2612) );
  INVXL U190 ( .A(wdata[15]), .Y(n2602) );
  INVXL U191 ( .A(wdata[29]), .Y(n2588) );
  INVXL U192 ( .A(wdata[30]), .Y(n2587) );
  INVXL U193 ( .A(wdata[11]), .Y(n2606) );
  INVXL U194 ( .A(wdata[18]), .Y(n2599) );
  INVXL U195 ( .A(wdata[2]), .Y(n2615) );
  INVXL U196 ( .A(wdata[23]), .Y(n2594) );
  INVXL U197 ( .A(wdata[13]), .Y(n2604) );
  INVXL U198 ( .A(wdata[17]), .Y(n2600) );
  INVXL U199 ( .A(wdata[16]), .Y(n2601) );
  INVXL U200 ( .A(wdata[19]), .Y(n2598) );
  INVXL U201 ( .A(wdata[21]), .Y(n2596) );
  INVXL U202 ( .A(wdata[26]), .Y(n2591) );
  INVXL U203 ( .A(wdata[28]), .Y(n2589) );
  INVXL U204 ( .A(wdata[20]), .Y(n2597) );
  INVXL U205 ( .A(wdata[0]), .Y(n2617) );
  INVXL U206 ( .A(wdata[4]), .Y(n2613) );
  INVXL U207 ( .A(wdata[6]), .Y(n2611) );
  INVXL U208 ( .A(wdata[8]), .Y(n2609) );
  INVXL U209 ( .A(wdata[9]), .Y(n2608) );
  INVXL U210 ( .A(wdata[10]), .Y(n2607) );
  MXI4XL U211 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n2151), .S1(n2126), 
        .Y(n1797) );
  MXI4XL U212 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n2148), .S1(n2124), .Y(
        n1733) );
  MXI4XL U213 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1600), .S1(n1578), .Y(
        n1143) );
  NOR2BXL U214 ( .AN(n1584), .B(\register[3][1] ), .Y(n1536) );
  MXI4XL U215 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n2151), .S1(n2127), .Y(
        n1738) );
  MXI4XL U216 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n2151), .S1(n2127), 
        .Y(n1798) );
  MXI4XL U217 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n2151), .S1(n2127), .Y(
        n1928) );
  MXI4XL U218 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n2151), .S1(n2127), 
        .Y(n1799) );
  MXI4XL U219 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n2148), .S1(n2124), .Y(
        n1734) );
  MXI4XL U220 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n2142), .S1(n2118), 
        .Y(n1834) );
  MXI4XL U221 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1606), .S1(n1582), 
        .Y(n1245) );
  MXI4XL U222 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1600), .S1(n1578), .Y(
        n1141) );
  MXI4XL U223 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n2148), .S1(n2124), .Y(
        n1732) );
  MXI4XL U224 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n1600), .S1(n1578), .Y(
        n1144) );
  MXI4XL U225 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1606), .S1(n1582), .Y(
        n1248) );
  MXI4XL U226 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n2148), .S1(n2124), .Y(
        n1731) );
  MXI4XL U227 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n2149), .S1(n2124), .Y(
        n1735) );
  MXI4XL U228 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n2142), .S1(n2118), 
        .Y(n1835) );
  MXI4XL U229 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1606), .S1(n1582), 
        .Y(n1243) );
  MXI4XL U230 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1606), .S1(n1582), 
        .Y(n1247) );
  MXI4XL U231 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1599), .S1(n1578), .Y(
        n1139) );
  NOR2X1 U232 ( .A(n2131), .B(n2151), .Y(n2006) );
  NOR2X1 U233 ( .A(n2131), .B(n2151), .Y(n2001) );
  NOR2X1 U234 ( .A(n2131), .B(n2151), .Y(n1991) );
  NOR2X1 U235 ( .A(n2132), .B(n2151), .Y(n1986) );
  NOR2X1 U236 ( .A(n2132), .B(n2145), .Y(n1981) );
  NOR2X1 U237 ( .A(n2132), .B(n2145), .Y(n1976) );
  NOR2X1 U238 ( .A(n2132), .B(n2145), .Y(n1971) );
  NOR2X1 U239 ( .A(n2132), .B(n2145), .Y(n1966) );
  NOR2X1 U240 ( .A(n1587), .B(n1599), .Y(n1462) );
  NOR2X1 U241 ( .A(n1587), .B(n1599), .Y(n1457) );
  NOR2X1 U242 ( .A(n1587), .B(n1599), .Y(n1447) );
  NOR2X1 U243 ( .A(n1574), .B(n1599), .Y(n1442) );
  NOR2X1 U244 ( .A(n1574), .B(n1599), .Y(n1437) );
  NOR2X1 U245 ( .A(n1574), .B(n1599), .Y(n1432) );
  NOR2X1 U246 ( .A(n1574), .B(n1599), .Y(n1427) );
  NOR2X1 U247 ( .A(n1573), .B(n1599), .Y(n1422) );
  NOR2X1 U248 ( .A(n2128), .B(n2154), .Y(n2086) );
  NOR2X1 U249 ( .A(n2128), .B(n2154), .Y(n2061) );
  NOR2X1 U250 ( .A(n1584), .B(n1599), .Y(n1542) );
  NOR2X1 U251 ( .A(n1584), .B(n1599), .Y(n1517) );
  NOR2X1 U252 ( .A(n2130), .B(n2145), .Y(n2081) );
  NOR2X1 U253 ( .A(n2129), .B(n2154), .Y(n2076) );
  NOR2X1 U254 ( .A(n2129), .B(n2145), .Y(n2071) );
  NOR2X1 U255 ( .A(n2129), .B(n2145), .Y(n2066) );
  NOR2X1 U256 ( .A(n2130), .B(n2153), .Y(n2056) );
  NOR2X1 U257 ( .A(n2129), .B(n2145), .Y(n2051) );
  NOR2X1 U258 ( .A(n2129), .B(n2154), .Y(n2046) );
  NOR2X1 U259 ( .A(n2129), .B(n2154), .Y(n2041) );
  NOR2X1 U260 ( .A(n2129), .B(n2154), .Y(n2036) );
  NOR2X1 U261 ( .A(n2130), .B(n2154), .Y(n2031) );
  NOR2X1 U262 ( .A(n2130), .B(n2154), .Y(n2026) );
  NOR2X1 U263 ( .A(n2130), .B(n2154), .Y(n2021) );
  NOR2X1 U264 ( .A(n2131), .B(n2154), .Y(n2016) );
  NOR2X1 U265 ( .A(n2131), .B(n2154), .Y(n2011) );
  NOR2X1 U266 ( .A(n2131), .B(n2154), .Y(n1996) );
  NOR2X1 U267 ( .A(n2132), .B(n2154), .Y(n1961) );
  NOR2X1 U268 ( .A(n1586), .B(n1599), .Y(n1537) );
  NOR2X1 U269 ( .A(n1585), .B(n1599), .Y(n1532) );
  NOR2X1 U270 ( .A(n1585), .B(n1599), .Y(n1527) );
  NOR2X1 U271 ( .A(n1585), .B(n1599), .Y(n1522) );
  NOR2X1 U272 ( .A(n1586), .B(n1599), .Y(n1512) );
  NOR2X1 U273 ( .A(n1585), .B(n1599), .Y(n1507) );
  NOR2X1 U274 ( .A(n1585), .B(n1609), .Y(n1502) );
  NOR2X1 U275 ( .A(n1585), .B(n1609), .Y(n1497) );
  NOR2X1 U276 ( .A(n1585), .B(n1609), .Y(n1492) );
  NOR2X1 U277 ( .A(n1586), .B(n1609), .Y(n1487) );
  NOR2X1 U278 ( .A(n1586), .B(n1609), .Y(n1482) );
  NOR2X1 U279 ( .A(n1586), .B(n1609), .Y(n1477) );
  NOR2X1 U280 ( .A(n1587), .B(n1609), .Y(n1472) );
  NOR2X1 U281 ( .A(n1587), .B(n1609), .Y(n1467) );
  NOR2X1 U282 ( .A(n1587), .B(n1609), .Y(n1452) );
  NOR2X1 U283 ( .A(n1577), .B(n1609), .Y(n1417) );
  CLKBUFX3 U284 ( .A(n2547), .Y(n2460) );
  CLKBUFX3 U285 ( .A(n2547), .Y(n2461) );
  CLKBUFX3 U286 ( .A(n2547), .Y(n2462) );
  CLKBUFX3 U287 ( .A(n2547), .Y(n2463) );
  CLKBUFX3 U288 ( .A(n2546), .Y(n2464) );
  CLKBUFX3 U289 ( .A(n2546), .Y(n2465) );
  CLKBUFX3 U290 ( .A(n2546), .Y(n2466) );
  CLKBUFX3 U291 ( .A(n2546), .Y(n2467) );
  CLKBUFX3 U292 ( .A(n2545), .Y(n2468) );
  CLKBUFX3 U293 ( .A(n2545), .Y(n2469) );
  CLKBUFX3 U294 ( .A(n2545), .Y(n2470) );
  CLKBUFX3 U295 ( .A(n2545), .Y(n2471) );
  CLKBUFX3 U296 ( .A(n2544), .Y(n2472) );
  CLKBUFX3 U297 ( .A(n2544), .Y(n2473) );
  CLKBUFX3 U298 ( .A(n2544), .Y(n2474) );
  CLKBUFX3 U299 ( .A(n2544), .Y(n2475) );
  CLKBUFX3 U300 ( .A(n2543), .Y(n2476) );
  CLKBUFX3 U301 ( .A(n2543), .Y(n2477) );
  CLKBUFX3 U302 ( .A(n2543), .Y(n2478) );
  CLKBUFX3 U303 ( .A(n2543), .Y(n2479) );
  CLKBUFX3 U304 ( .A(n2542), .Y(n2480) );
  CLKBUFX3 U305 ( .A(n2542), .Y(n2481) );
  CLKBUFX3 U306 ( .A(n2542), .Y(n2482) );
  CLKBUFX3 U307 ( .A(n2542), .Y(n2483) );
  CLKBUFX3 U308 ( .A(n2541), .Y(n2484) );
  CLKBUFX3 U309 ( .A(n2541), .Y(n2485) );
  CLKBUFX3 U310 ( .A(n2541), .Y(n2486) );
  CLKBUFX3 U311 ( .A(n2541), .Y(n2487) );
  CLKBUFX3 U312 ( .A(n2540), .Y(n2488) );
  CLKBUFX3 U313 ( .A(n2540), .Y(n2489) );
  CLKBUFX3 U314 ( .A(n2540), .Y(n2490) );
  CLKBUFX3 U315 ( .A(n2540), .Y(n2491) );
  CLKBUFX3 U316 ( .A(n2539), .Y(n2492) );
  CLKBUFX3 U317 ( .A(n2539), .Y(n2493) );
  CLKBUFX3 U318 ( .A(n2539), .Y(n2494) );
  CLKBUFX3 U319 ( .A(n2539), .Y(n2495) );
  CLKBUFX3 U320 ( .A(n2538), .Y(n2496) );
  CLKBUFX3 U321 ( .A(n2538), .Y(n2497) );
  CLKBUFX3 U322 ( .A(n2538), .Y(n2498) );
  CLKBUFX3 U323 ( .A(n2538), .Y(n2499) );
  CLKBUFX3 U324 ( .A(n2537), .Y(n2500) );
  CLKBUFX3 U325 ( .A(n2537), .Y(n2501) );
  CLKBUFX3 U326 ( .A(n2537), .Y(n2502) );
  CLKBUFX3 U327 ( .A(n2537), .Y(n2503) );
  CLKBUFX3 U328 ( .A(n2536), .Y(n2504) );
  CLKBUFX3 U329 ( .A(n2536), .Y(n2505) );
  CLKBUFX3 U330 ( .A(n2536), .Y(n2506) );
  CLKBUFX3 U331 ( .A(n2536), .Y(n2507) );
  CLKBUFX3 U332 ( .A(n2535), .Y(n2508) );
  CLKBUFX3 U333 ( .A(n2535), .Y(n2509) );
  CLKBUFX3 U334 ( .A(n2535), .Y(n2510) );
  CLKBUFX3 U335 ( .A(n2535), .Y(n2511) );
  CLKBUFX3 U336 ( .A(n2534), .Y(n2512) );
  CLKBUFX3 U337 ( .A(n2534), .Y(n2513) );
  CLKBUFX3 U338 ( .A(n2534), .Y(n2514) );
  CLKBUFX3 U339 ( .A(n2534), .Y(n2515) );
  CLKBUFX3 U340 ( .A(n2551), .Y(n2516) );
  CLKBUFX3 U341 ( .A(n2551), .Y(n2517) );
  CLKBUFX3 U342 ( .A(n2535), .Y(n2518) );
  CLKBUFX3 U343 ( .A(n2552), .Y(n2519) );
  CLKBUFX3 U344 ( .A(n2533), .Y(n2520) );
  CLKBUFX3 U345 ( .A(n2533), .Y(n2521) );
  CLKBUFX3 U346 ( .A(n2533), .Y(n2522) );
  CLKBUFX3 U347 ( .A(n2533), .Y(n2523) );
  CLKBUFX3 U348 ( .A(n2532), .Y(n2524) );
  CLKBUFX3 U349 ( .A(n2532), .Y(n2525) );
  CLKBUFX3 U350 ( .A(n2532), .Y(n2526) );
  CLKBUFX3 U351 ( .A(n2532), .Y(n2527) );
  CLKBUFX3 U352 ( .A(n2553), .Y(n2528) );
  CLKBUFX3 U353 ( .A(n2553), .Y(n2529) );
  CLKBUFX3 U354 ( .A(n2533), .Y(n2530) );
  CLKBUFX3 U355 ( .A(n2548), .Y(n2531) );
  CLKBUFX3 U356 ( .A(n2136), .Y(n2152) );
  CLKBUFX3 U357 ( .A(n2136), .Y(n2153) );
  CLKBUFX3 U358 ( .A(n1593), .Y(n1607) );
  CLKBUFX3 U359 ( .A(n1592), .Y(n1608) );
  NOR2X1 U360 ( .A(n2133), .B(n2154), .Y(n1956) );
  NOR2X1 U361 ( .A(n2133), .B(n2154), .Y(n1951) );
  NOR2X1 U362 ( .A(n2133), .B(n2145), .Y(n1946) );
  NOR2X1 U363 ( .A(n2133), .B(n2145), .Y(n1941) );
  NOR2X1 U364 ( .A(n2133), .B(n2145), .Y(n1936) );
  NOR2X1 U365 ( .A(n2133), .B(n2154), .Y(n1931) );
  NOR2X1 U366 ( .A(n1588), .B(n1609), .Y(n1407) );
  NOR2X1 U367 ( .A(n1588), .B(n1599), .Y(n1402) );
  NOR2X1 U368 ( .A(n1588), .B(n1599), .Y(n1397) );
  NOR2X1 U369 ( .A(n1588), .B(n1599), .Y(n1392) );
  NOR2X1 U370 ( .A(n1588), .B(n1599), .Y(n1387) );
  CLKBUFX3 U371 ( .A(n2138), .Y(n2146) );
  CLKBUFX3 U372 ( .A(n2138), .Y(n2147) );
  CLKBUFX3 U373 ( .A(n2137), .Y(n2148) );
  CLKBUFX3 U374 ( .A(n2136), .Y(n2150) );
  CLKBUFX3 U375 ( .A(n2137), .Y(n2149) );
  CLKBUFX3 U376 ( .A(n2140), .Y(n2142) );
  CLKBUFX3 U377 ( .A(n2139), .Y(n2143) );
  CLKBUFX3 U378 ( .A(n2139), .Y(n2144) );
  CLKBUFX3 U379 ( .A(n1591), .Y(n1600) );
  CLKBUFX3 U380 ( .A(n1594), .Y(n1601) );
  CLKBUFX3 U381 ( .A(n1594), .Y(n1602) );
  CLKBUFX3 U382 ( .A(n1591), .Y(n1604) );
  CLKBUFX3 U383 ( .A(n1591), .Y(n1605) );
  CLKBUFX3 U384 ( .A(n1594), .Y(n1603) );
  CLKBUFX3 U385 ( .A(n1594), .Y(n1595) );
  CLKBUFX3 U386 ( .A(n1591), .Y(n1597) );
  CLKBUFX3 U387 ( .A(n1591), .Y(n1598) );
  CLKBUFX3 U388 ( .A(n1590), .Y(n1596) );
  BUFX4 U389 ( .A(n2114), .Y(n2123) );
  BUFX4 U390 ( .A(n2113), .Y(n2125) );
  BUFX4 U391 ( .A(n2113), .Y(n2126) );
  BUFX4 U392 ( .A(n2107), .Y(n2117) );
  BUFX4 U393 ( .A(n2107), .Y(n2118) );
  BUFX4 U394 ( .A(n2116), .Y(n2120) );
  BUFX4 U395 ( .A(n2115), .Y(n2122) );
  BUFX4 U396 ( .A(n2116), .Y(n2119) );
  BUFX4 U397 ( .A(n2115), .Y(n2121) );
  BUFX4 U398 ( .A(n1571), .Y(n1579) );
  BUFX4 U399 ( .A(n1570), .Y(n1581) );
  BUFX4 U400 ( .A(n1571), .Y(n1580) );
  BUFX4 U401 ( .A(n1570), .Y(n1582) );
  BUFX4 U402 ( .A(n1572), .Y(n1573) );
  BUFX4 U403 ( .A(n1567), .Y(n1574) );
  BUFX4 U404 ( .A(n1570), .Y(n1576) );
  BUFX4 U405 ( .A(n1572), .Y(n1578) );
  BUFX4 U406 ( .A(n1570), .Y(n1575) );
  BUFX4 U407 ( .A(n1572), .Y(n1577) );
  CLKBUFX3 U408 ( .A(n2134), .Y(n2128) );
  CLKBUFX3 U409 ( .A(n1569), .Y(n1584) );
  CLKBUFX3 U410 ( .A(n2112), .Y(n2129) );
  CLKBUFX3 U411 ( .A(n2112), .Y(n2130) );
  CLKBUFX3 U412 ( .A(n2111), .Y(n2132) );
  CLKBUFX3 U413 ( .A(n1568), .Y(n1585) );
  CLKBUFX3 U414 ( .A(n1568), .Y(n1586) );
  CLKBUFX3 U415 ( .A(n2549), .Y(n2452) );
  CLKBUFX3 U416 ( .A(n2549), .Y(n2453) );
  CLKBUFX3 U417 ( .A(n2448), .Y(n2454) );
  CLKBUFX3 U418 ( .A(n2447), .Y(n2455) );
  CLKBUFX3 U419 ( .A(n2548), .Y(n2456) );
  CLKBUFX3 U420 ( .A(n2548), .Y(n2457) );
  CLKBUFX3 U421 ( .A(n2548), .Y(n2458) );
  CLKBUFX3 U422 ( .A(n2548), .Y(n2459) );
  CLKBUFX3 U423 ( .A(n2549), .Y(n2449) );
  CLKBUFX3 U424 ( .A(n2549), .Y(n2450) );
  CLKBUFX3 U425 ( .A(n2447), .Y(n2451) );
  CLKBUFX3 U426 ( .A(n2550), .Y(n2547) );
  CLKBUFX3 U427 ( .A(n2550), .Y(n2546) );
  CLKBUFX3 U428 ( .A(n2550), .Y(n2545) );
  CLKBUFX3 U429 ( .A(n2551), .Y(n2544) );
  CLKBUFX3 U430 ( .A(n2551), .Y(n2543) );
  CLKBUFX3 U431 ( .A(n2551), .Y(n2542) );
  CLKBUFX3 U432 ( .A(n2552), .Y(n2541) );
  CLKBUFX3 U433 ( .A(n2552), .Y(n2540) );
  CLKBUFX3 U434 ( .A(n2552), .Y(n2539) );
  CLKBUFX3 U435 ( .A(n2553), .Y(n2538) );
  CLKBUFX3 U436 ( .A(n2553), .Y(n2537) );
  CLKBUFX3 U437 ( .A(n2553), .Y(n2536) );
  CLKBUFX3 U438 ( .A(n2447), .Y(n2535) );
  CLKBUFX3 U439 ( .A(n2550), .Y(n2534) );
  CLKBUFX3 U440 ( .A(n2448), .Y(n2533) );
  CLKBUFX3 U441 ( .A(n2552), .Y(n2532) );
  CLKBUFX3 U442 ( .A(n2099), .Y(n2095) );
  CLKBUFX3 U443 ( .A(n2099), .Y(n2096) );
  CLKBUFX3 U444 ( .A(n2099), .Y(n2097) );
  CLKBUFX3 U445 ( .A(n2099), .Y(n2098) );
  CLKBUFX3 U446 ( .A(n1558), .Y(n1554) );
  CLKBUFX3 U447 ( .A(n1558), .Y(n1555) );
  CLKBUFX3 U448 ( .A(n1550), .Y(n1556) );
  CLKBUFX3 U449 ( .A(n1550), .Y(n1557) );
  CLKBUFX3 U450 ( .A(n2110), .Y(n2133) );
  CLKBUFX3 U451 ( .A(n2109), .Y(n2110) );
  CLKBUFX3 U452 ( .A(n1571), .Y(n1588) );
  CLKBUFX3 U453 ( .A(n2251), .Y(n2254) );
  CLKBUFX3 U454 ( .A(n2251), .Y(n2252) );
  CLKBUFX3 U455 ( .A(n2251), .Y(n2253) );
  CLKBUFX3 U456 ( .A(n2106), .Y(n2102) );
  CLKBUFX3 U457 ( .A(n2106), .Y(n2103) );
  CLKBUFX3 U458 ( .A(n2100), .Y(n2104) );
  CLKBUFX3 U459 ( .A(n2106), .Y(n2105) );
  CLKBUFX3 U460 ( .A(n1559), .Y(n1562) );
  CLKBUFX3 U461 ( .A(n1559), .Y(n1563) );
  CLKBUFX3 U462 ( .A(n1560), .Y(n1564) );
  CLKBUFX3 U463 ( .A(n1560), .Y(n1565) );
  CLKBUFX3 U464 ( .A(N13), .Y(n1569) );
  CLKBUFX3 U465 ( .A(n2109), .Y(n2112) );
  CLKBUFX3 U466 ( .A(n2109), .Y(n2111) );
  CLKBUFX3 U467 ( .A(n1589), .Y(n1568) );
  CLKBUFX3 U468 ( .A(n2108), .Y(n2114) );
  CLKBUFX3 U469 ( .A(n2108), .Y(n2113) );
  CLKBUFX3 U470 ( .A(n2107), .Y(n2116) );
  CLKBUFX3 U471 ( .A(n2107), .Y(n2115) );
  CLKBUFX3 U472 ( .A(n1567), .Y(n1571) );
  CLKBUFX3 U473 ( .A(n1567), .Y(n1570) );
  CLKBUFX3 U474 ( .A(n2135), .Y(n2137) );
  CLKBUFX3 U475 ( .A(n2136), .Y(n2139) );
  CLKBUFX3 U476 ( .A(n1591), .Y(n1593) );
  CLKBUFX3 U477 ( .A(n2448), .Y(n2550) );
  CLKBUFX3 U478 ( .A(n2448), .Y(n2551) );
  CLKBUFX3 U479 ( .A(n2447), .Y(n2552) );
  CLKBUFX3 U480 ( .A(n2447), .Y(n2553) );
  CLKBUFX3 U481 ( .A(n2549), .Y(n2548) );
  CLKBUFX3 U482 ( .A(n2093), .Y(n2091) );
  CLKBUFX3 U483 ( .A(n2093), .Y(n2092) );
  CLKBUFX3 U484 ( .A(n1549), .Y(n1547) );
  CLKBUFX3 U485 ( .A(n1549), .Y(n1548) );
  CLKBUFX3 U486 ( .A(n2418), .Y(n2421) );
  CLKBUFX3 U487 ( .A(n2409), .Y(n2414) );
  CLKBUFX3 U488 ( .A(n2371), .Y(n2374) );
  CLKBUFX3 U489 ( .A(n2365), .Y(n2368) );
  CLKBUFX3 U490 ( .A(n2327), .Y(n2330) );
  CLKBUFX3 U491 ( .A(n2321), .Y(n2324) );
  CLKBUFX3 U492 ( .A(n2279), .Y(n2282) );
  CLKBUFX3 U493 ( .A(n2273), .Y(n2276) );
  CLKBUFX3 U494 ( .A(n2424), .Y(n2427) );
  CLKBUFX3 U495 ( .A(n2377), .Y(n2380) );
  CLKBUFX3 U496 ( .A(n92), .Y(n2335) );
  CLKBUFX3 U497 ( .A(n2284), .Y(n2288) );
  CLKBUFX3 U498 ( .A(n2359), .Y(n2362) );
  CLKBUFX3 U499 ( .A(n88), .Y(n2350) );
  CLKBUFX3 U500 ( .A(n2315), .Y(n2318) );
  CLKBUFX3 U501 ( .A(n97), .Y(n2306) );
  CLKBUFX3 U502 ( .A(n2266), .Y(n2270) );
  CLKBUFX3 U503 ( .A(n2256), .Y(n2260) );
  CLKBUFX3 U504 ( .A(n2404), .Y(n2407) );
  CLKBUFX3 U505 ( .A(n76), .Y(n2395) );
  CLKBUFX3 U506 ( .A(n2383), .Y(n2386) );
  CLKBUFX3 U507 ( .A(n2337), .Y(n2340) );
  CLKBUFX3 U508 ( .A(n2291), .Y(n2294) );
  CLKBUFX3 U509 ( .A(n87), .Y(n2356) );
  CLKBUFX3 U510 ( .A(n96), .Y(n2312) );
  CLKBUFX3 U511 ( .A(n98), .Y(n2300) );
  CLKBUFX3 U512 ( .A(n105), .Y(n2264) );
  CLKBUFX3 U513 ( .A(n74), .Y(n2401) );
  CLKBUFX3 U514 ( .A(n2418), .Y(n2422) );
  CLKBUFX3 U515 ( .A(n2409), .Y(n2415) );
  CLKBUFX3 U516 ( .A(n2371), .Y(n2375) );
  CLKBUFX3 U517 ( .A(n2365), .Y(n2369) );
  CLKBUFX3 U518 ( .A(n2327), .Y(n2331) );
  CLKBUFX3 U519 ( .A(n2321), .Y(n2325) );
  CLKBUFX3 U520 ( .A(n2279), .Y(n2283) );
  CLKBUFX3 U521 ( .A(n2273), .Y(n2277) );
  CLKBUFX3 U522 ( .A(n2424), .Y(n2428) );
  CLKBUFX3 U523 ( .A(n2377), .Y(n2381) );
  CLKBUFX3 U524 ( .A(n92), .Y(n2336) );
  CLKBUFX3 U525 ( .A(n2284), .Y(n2289) );
  CLKBUFX3 U526 ( .A(n2359), .Y(n2363) );
  CLKBUFX3 U527 ( .A(n2347), .Y(n2351) );
  CLKBUFX3 U528 ( .A(n2315), .Y(n2319) );
  CLKBUFX3 U529 ( .A(n2303), .Y(n2307) );
  CLKBUFX3 U530 ( .A(n2266), .Y(n2271) );
  CLKBUFX3 U531 ( .A(n2256), .Y(n2261) );
  CLKBUFX3 U532 ( .A(n2404), .Y(n2408) );
  CLKBUFX3 U533 ( .A(n76), .Y(n2396) );
  CLKBUFX3 U534 ( .A(n2383), .Y(n2387) );
  CLKBUFX3 U535 ( .A(n2337), .Y(n2341) );
  CLKBUFX3 U536 ( .A(n2291), .Y(n2295) );
  CLKBUFX3 U537 ( .A(n2353), .Y(n2357) );
  CLKBUFX3 U538 ( .A(n2309), .Y(n2313) );
  CLKBUFX3 U539 ( .A(n105), .Y(n2265) );
  CLKBUFX3 U540 ( .A(n2398), .Y(n2402) );
  CLKBUFX3 U541 ( .A(n2389), .Y(n2392) );
  CLKBUFX3 U542 ( .A(n2418), .Y(n2419) );
  CLKBUFX3 U543 ( .A(n2418), .Y(n2420) );
  CLKBUFX3 U544 ( .A(n2410), .Y(n2412) );
  CLKBUFX3 U545 ( .A(n2409), .Y(n2413) );
  CLKBUFX3 U546 ( .A(n2371), .Y(n2372) );
  CLKBUFX3 U547 ( .A(n2371), .Y(n2373) );
  CLKBUFX3 U548 ( .A(n2365), .Y(n2366) );
  CLKBUFX3 U549 ( .A(n2365), .Y(n2367) );
  CLKBUFX3 U550 ( .A(n2327), .Y(n2328) );
  CLKBUFX3 U551 ( .A(n2327), .Y(n2329) );
  CLKBUFX3 U552 ( .A(n2321), .Y(n2322) );
  CLKBUFX3 U553 ( .A(n2321), .Y(n2323) );
  CLKBUFX3 U554 ( .A(n2279), .Y(n2280) );
  CLKBUFX3 U555 ( .A(n2279), .Y(n2281) );
  CLKBUFX3 U556 ( .A(n2273), .Y(n2274) );
  CLKBUFX3 U557 ( .A(n2273), .Y(n2275) );
  CLKBUFX3 U558 ( .A(n2424), .Y(n2425) );
  CLKBUFX3 U559 ( .A(n2424), .Y(n2426) );
  CLKBUFX3 U560 ( .A(n2377), .Y(n2378) );
  CLKBUFX3 U561 ( .A(n2377), .Y(n2379) );
  CLKBUFX3 U562 ( .A(n2332), .Y(n2333) );
  CLKBUFX3 U563 ( .A(n2332), .Y(n2334) );
  CLKBUFX3 U564 ( .A(n2284), .Y(n2286) );
  CLKBUFX3 U565 ( .A(n2284), .Y(n2287) );
  CLKBUFX3 U566 ( .A(n2383), .Y(n2384) );
  CLKBUFX3 U567 ( .A(n2383), .Y(n2385) );
  CLKBUFX3 U568 ( .A(n2337), .Y(n2339) );
  CLKBUFX3 U569 ( .A(n2291), .Y(n2292) );
  CLKBUFX3 U570 ( .A(n2291), .Y(n2293) );
  CLKBUFX3 U571 ( .A(n2359), .Y(n2360) );
  CLKBUFX3 U572 ( .A(n2359), .Y(n2361) );
  CLKBUFX3 U573 ( .A(n2347), .Y(n2348) );
  CLKBUFX3 U574 ( .A(n2347), .Y(n2349) );
  CLKBUFX3 U575 ( .A(n2315), .Y(n2316) );
  CLKBUFX3 U576 ( .A(n2315), .Y(n2317) );
  CLKBUFX3 U577 ( .A(n2303), .Y(n2304) );
  CLKBUFX3 U578 ( .A(n2303), .Y(n2305) );
  CLKBUFX3 U579 ( .A(n2266), .Y(n2268) );
  CLKBUFX3 U580 ( .A(n2266), .Y(n2269) );
  CLKBUFX3 U581 ( .A(n2256), .Y(n2258) );
  CLKBUFX3 U582 ( .A(n2256), .Y(n2259) );
  CLKBUFX3 U583 ( .A(n2404), .Y(n2405) );
  CLKBUFX3 U584 ( .A(n2404), .Y(n2406) );
  CLKBUFX3 U585 ( .A(n76), .Y(n2393) );
  CLKBUFX3 U586 ( .A(n76), .Y(n2394) );
  CLKBUFX3 U587 ( .A(n2353), .Y(n2354) );
  CLKBUFX3 U588 ( .A(n2353), .Y(n2355) );
  CLKBUFX3 U589 ( .A(n2343), .Y(n2344) );
  CLKBUFX3 U590 ( .A(n2343), .Y(n2345) );
  CLKBUFX3 U591 ( .A(n2309), .Y(n2310) );
  CLKBUFX3 U592 ( .A(n2309), .Y(n2311) );
  CLKBUFX3 U593 ( .A(n2297), .Y(n2298) );
  CLKBUFX3 U594 ( .A(n2297), .Y(n2299) );
  CLKBUFX3 U595 ( .A(n105), .Y(n2263) );
  CLKBUFX3 U596 ( .A(n2398), .Y(n2399) );
  CLKBUFX3 U597 ( .A(n2398), .Y(n2400) );
  CLKBUFX3 U598 ( .A(n2389), .Y(n2391) );
  CLKBUFX3 U599 ( .A(N17), .Y(n2135) );
  CLKBUFX3 U600 ( .A(N12), .Y(n1590) );
  CLKBUFX3 U601 ( .A(N17), .Y(n2136) );
  CLKBUFX3 U602 ( .A(N12), .Y(n1591) );
  CLKBUFX3 U603 ( .A(n2443), .Y(n1592) );
  CLKBUFX3 U604 ( .A(n2134), .Y(n2108) );
  CLKBUFX3 U605 ( .A(n2134), .Y(n2109) );
  CLKBUFX3 U606 ( .A(n2134), .Y(n2107) );
  CLKBUFX3 U607 ( .A(n1558), .Y(n1551) );
  CLKBUFX3 U608 ( .A(n1566), .Y(n1559) );
  CLKBUFX3 U609 ( .A(n1558), .Y(n1550) );
  CLKBUFX3 U610 ( .A(n2251), .Y(n2250) );
  CLKBUFX3 U611 ( .A(n2448), .Y(n2549) );
  NOR4X1 U612 ( .A(n55), .B(n2440), .C(n2442), .D(n2441), .Y(n52) );
  OR2X1 U613 ( .A(n2439), .B(N18), .Y(n55) );
  NOR4X1 U614 ( .A(n64), .B(n2444), .C(n2446), .D(n2445), .Y(n61) );
  CLKBUFX3 U615 ( .A(n2434), .Y(n2437) );
  CLKBUFX3 U616 ( .A(n2617), .Y(n2248) );
  CLKBUFX3 U617 ( .A(n2616), .Y(n2245) );
  CLKBUFX3 U618 ( .A(n2614), .Y(n2240) );
  CLKBUFX3 U619 ( .A(n2613), .Y(n2237) );
  CLKBUFX3 U620 ( .A(n2612), .Y(n2234) );
  CLKBUFX3 U621 ( .A(n2611), .Y(n2231) );
  CLKBUFX3 U622 ( .A(n2610), .Y(n2228) );
  CLKBUFX3 U623 ( .A(n2609), .Y(n2225) );
  CLKBUFX3 U624 ( .A(n2608), .Y(n2222) );
  CLKBUFX3 U625 ( .A(n2606), .Y(n2216) );
  CLKBUFX3 U626 ( .A(n2605), .Y(n2213) );
  CLKBUFX3 U627 ( .A(n2604), .Y(n2210) );
  CLKBUFX3 U628 ( .A(n2603), .Y(n2207) );
  CLKBUFX3 U629 ( .A(n2601), .Y(n2201) );
  CLKBUFX3 U630 ( .A(n2600), .Y(n2198) );
  CLKBUFX3 U631 ( .A(n2598), .Y(n2192) );
  CLKBUFX3 U632 ( .A(n2597), .Y(n2189) );
  CLKBUFX3 U633 ( .A(n2595), .Y(n2183) );
  CLKBUFX3 U634 ( .A(n2593), .Y(n2177) );
  CLKBUFX3 U635 ( .A(n2592), .Y(n2174) );
  CLKBUFX3 U636 ( .A(n2590), .Y(n2168) );
  CLKBUFX3 U637 ( .A(n2586), .Y(n2156) );
  CLKBUFX3 U638 ( .A(n2617), .Y(n2247) );
  CLKBUFX3 U639 ( .A(n2616), .Y(n2244) );
  CLKBUFX3 U640 ( .A(n2614), .Y(n2239) );
  CLKBUFX3 U641 ( .A(n2613), .Y(n2236) );
  CLKBUFX3 U642 ( .A(n2612), .Y(n2233) );
  CLKBUFX3 U643 ( .A(n2611), .Y(n2230) );
  CLKBUFX3 U644 ( .A(n2610), .Y(n2227) );
  CLKBUFX3 U645 ( .A(n2609), .Y(n2224) );
  CLKBUFX3 U646 ( .A(n2608), .Y(n2221) );
  CLKBUFX3 U647 ( .A(n2606), .Y(n2215) );
  CLKBUFX3 U648 ( .A(n2605), .Y(n2212) );
  CLKBUFX3 U649 ( .A(n2604), .Y(n2209) );
  CLKBUFX3 U650 ( .A(n2603), .Y(n2206) );
  CLKBUFX3 U651 ( .A(n2601), .Y(n2200) );
  CLKBUFX3 U652 ( .A(n2600), .Y(n2197) );
  CLKBUFX3 U653 ( .A(n2598), .Y(n2191) );
  CLKBUFX3 U654 ( .A(n2597), .Y(n2188) );
  CLKBUFX3 U655 ( .A(n2595), .Y(n2182) );
  CLKBUFX3 U656 ( .A(n2593), .Y(n2176) );
  CLKBUFX3 U657 ( .A(n2592), .Y(n2173) );
  CLKBUFX3 U658 ( .A(n2590), .Y(n2167) );
  CLKBUFX3 U659 ( .A(n2586), .Y(n2155) );
  CLKBUFX3 U660 ( .A(n2615), .Y(n2242) );
  CLKBUFX3 U661 ( .A(n2607), .Y(n2219) );
  CLKBUFX3 U662 ( .A(n2602), .Y(n2204) );
  CLKBUFX3 U663 ( .A(n2599), .Y(n2195) );
  CLKBUFX3 U664 ( .A(n2596), .Y(n2186) );
  CLKBUFX3 U665 ( .A(n2594), .Y(n2180) );
  CLKBUFX3 U666 ( .A(n2591), .Y(n2171) );
  CLKBUFX3 U667 ( .A(n2589), .Y(n2165) );
  CLKBUFX3 U668 ( .A(n2588), .Y(n2162) );
  CLKBUFX3 U669 ( .A(n2587), .Y(n2159) );
  CLKBUFX3 U670 ( .A(n2615), .Y(n2241) );
  CLKBUFX3 U671 ( .A(n2607), .Y(n2218) );
  CLKBUFX3 U672 ( .A(n2602), .Y(n2203) );
  CLKBUFX3 U673 ( .A(n2599), .Y(n2194) );
  CLKBUFX3 U674 ( .A(n2596), .Y(n2185) );
  CLKBUFX3 U675 ( .A(n2594), .Y(n2179) );
  CLKBUFX3 U676 ( .A(n2591), .Y(n2170) );
  CLKBUFX3 U677 ( .A(n2589), .Y(n2164) );
  CLKBUFX3 U678 ( .A(n2588), .Y(n2161) );
  CLKBUFX3 U679 ( .A(n2587), .Y(n2158) );
  CLKBUFX3 U680 ( .A(n2429), .Y(n2432) );
  CLKBUFX3 U681 ( .A(n2434), .Y(n2436) );
  CLKBUFX3 U682 ( .A(n2434), .Y(n2435) );
  CLKBUFX3 U683 ( .A(n2429), .Y(n2433) );
  CLKBUFX3 U684 ( .A(n2429), .Y(n2431) );
  CLKBUFX3 U685 ( .A(n2429), .Y(n2430) );
  CLKBUFX3 U686 ( .A(n2617), .Y(n2249) );
  CLKBUFX3 U687 ( .A(n2616), .Y(n2246) );
  CLKBUFX3 U688 ( .A(n2613), .Y(n2238) );
  CLKBUFX3 U689 ( .A(n2612), .Y(n2235) );
  CLKBUFX3 U690 ( .A(n2611), .Y(n2232) );
  CLKBUFX3 U691 ( .A(n2610), .Y(n2229) );
  CLKBUFX3 U692 ( .A(n2609), .Y(n2226) );
  CLKBUFX3 U693 ( .A(n2608), .Y(n2223) );
  CLKBUFX3 U694 ( .A(n2606), .Y(n2217) );
  CLKBUFX3 U695 ( .A(n2605), .Y(n2214) );
  CLKBUFX3 U696 ( .A(n2604), .Y(n2211) );
  CLKBUFX3 U697 ( .A(n2603), .Y(n2208) );
  CLKBUFX3 U698 ( .A(n2601), .Y(n2202) );
  CLKBUFX3 U699 ( .A(n2600), .Y(n2199) );
  CLKBUFX3 U700 ( .A(n2598), .Y(n2193) );
  CLKBUFX3 U701 ( .A(n2597), .Y(n2190) );
  CLKBUFX3 U702 ( .A(n2595), .Y(n2184) );
  CLKBUFX3 U703 ( .A(n2593), .Y(n2178) );
  CLKBUFX3 U704 ( .A(n2592), .Y(n2175) );
  CLKBUFX3 U705 ( .A(n2590), .Y(n2169) );
  CLKBUFX3 U706 ( .A(n2586), .Y(n2157) );
  CLKBUFX3 U707 ( .A(n2602), .Y(n2205) );
  CLKBUFX3 U708 ( .A(n2589), .Y(n2166) );
  CLKBUFX3 U709 ( .A(n2588), .Y(n2163) );
  CLKBUFX3 U710 ( .A(n2587), .Y(n2160) );
  CLKBUFX3 U711 ( .A(n2615), .Y(n2243) );
  CLKBUFX3 U712 ( .A(n2607), .Y(n2220) );
  CLKBUFX3 U713 ( .A(n2599), .Y(n2196) );
  CLKBUFX3 U714 ( .A(n2596), .Y(n2187) );
  CLKBUFX3 U715 ( .A(n2594), .Y(n2181) );
  CLKBUFX3 U716 ( .A(n2591), .Y(n2172) );
  CLKBUFX3 U717 ( .A(n2093), .Y(n2090) );
  CLKBUFX3 U718 ( .A(n2389), .Y(n2388) );
  CLKBUFX3 U719 ( .A(n2297), .Y(n2296) );
  CLKBUFX3 U720 ( .A(n105), .Y(n2262) );
  NOR3X2 U721 ( .A(n2618), .B(n14), .C(n2621), .Y(n100) );
  XNOR2X1 U722 ( .A(n2618), .B(n2441), .Y(n54) );
  XNOR2X1 U723 ( .A(n14), .B(n2442), .Y(n53) );
  NAND2XL U724 ( .A(n16), .B(n69), .Y(n84) );
  NAND2XL U725 ( .A(n16), .B(n71), .Y(n85) );
  NAND2XL U726 ( .A(n91), .B(n69), .Y(n93) );
  NAND2XL U727 ( .A(n91), .B(n71), .Y(n94) );
  NAND2XL U728 ( .A(n16), .B(n9), .Y(n83) );
  CLKBUFX3 U729 ( .A(N16), .Y(n2446) );
  BUFX2 U730 ( .A(n80), .Y(n2383) );
  NAND2X1 U731 ( .A(n16), .B(n5), .Y(n80) );
  NAND2X1 U732 ( .A(n91), .B(n5), .Y(n90) );
  BUFX2 U733 ( .A(n99), .Y(n2291) );
  NAND2X1 U734 ( .A(n100), .B(n5), .Y(n99) );
  NAND2X1 U735 ( .A(n16), .B(n13), .Y(n88) );
  NAND2X1 U736 ( .A(n91), .B(n13), .Y(n97) );
  NAND2X1 U737 ( .A(n13), .B(n7), .Y(n76) );
  NAND2X1 U738 ( .A(n16), .B(n11), .Y(n87) );
  NAND2X1 U739 ( .A(n91), .B(n11), .Y(n96) );
  NAND2X1 U740 ( .A(n11), .B(n7), .Y(n74) );
  NAND2X1 U741 ( .A(n79), .B(n7), .Y(n78) );
  CLKBUFX3 U742 ( .A(N20), .Y(n2441) );
  CLKBUFX3 U743 ( .A(N15), .Y(n2445) );
  CLKBUFX3 U744 ( .A(N19), .Y(n2440) );
  CLKBUFX3 U745 ( .A(N14), .Y(n2444) );
  CLKBUFX3 U746 ( .A(n2434), .Y(n2438) );
  OAI2BB2XL U747 ( .B0(n2437), .B1(n2249), .A0N(N91), .A1N(n2438), .Y(
        rdata2[0]) );
  OAI2BB2XL U748 ( .B0(n2436), .B1(n2246), .A0N(N90), .A1N(n2437), .Y(
        rdata2[1]) );
  OAI2BB2XL U749 ( .B0(n2435), .B1(n2243), .A0N(N89), .A1N(n2438), .Y(
        rdata2[2]) );
  OAI2BB2XL U750 ( .B0(n2435), .B1(n2614), .A0N(N88), .A1N(n2438), .Y(
        rdata2[3]) );
  OAI2BB2XL U751 ( .B0(n2435), .B1(n2238), .A0N(N87), .A1N(n2438), .Y(
        rdata2[4]) );
  OAI2BB2XL U752 ( .B0(n2435), .B1(n2235), .A0N(N86), .A1N(n2438), .Y(
        rdata2[5]) );
  OAI2BB2XL U753 ( .B0(n2435), .B1(n2232), .A0N(N85), .A1N(n2438), .Y(
        rdata2[6]) );
  OAI2BB2XL U754 ( .B0(n2435), .B1(n2229), .A0N(N84), .A1N(n2438), .Y(
        rdata2[7]) );
  OAI2BB2XL U755 ( .B0(n2435), .B1(n2226), .A0N(N83), .A1N(n2438), .Y(
        rdata2[8]) );
  OAI2BB2XL U756 ( .B0(n2436), .B1(n2223), .A0N(N82), .A1N(n2438), .Y(
        rdata2[9]) );
  OAI2BB2XL U757 ( .B0(n2437), .B1(n2220), .A0N(N81), .A1N(n2438), .Y(
        rdata2[10]) );
  OAI2BB2XL U758 ( .B0(n2437), .B1(n2217), .A0N(N80), .A1N(n2438), .Y(
        rdata2[11]) );
  OAI2BB2XL U759 ( .B0(n2437), .B1(n2214), .A0N(N79), .A1N(n2436), .Y(
        rdata2[12]) );
  OAI2BB2XL U760 ( .B0(n2437), .B1(n2211), .A0N(N78), .A1N(n2436), .Y(
        rdata2[13]) );
  OAI2BB2XL U761 ( .B0(n2437), .B1(n2208), .A0N(N77), .A1N(n2435), .Y(
        rdata2[14]) );
  OAI2BB2XL U762 ( .B0(n2437), .B1(n2205), .A0N(N76), .A1N(n2435), .Y(
        rdata2[15]) );
  OAI2BB2XL U763 ( .B0(n2436), .B1(n2202), .A0N(N75), .A1N(n2438), .Y(
        rdata2[16]) );
  OAI2BB2XL U764 ( .B0(n2437), .B1(n2199), .A0N(N74), .A1N(n2437), .Y(
        rdata2[17]) );
  OAI2BB2XL U765 ( .B0(n2436), .B1(n2196), .A0N(N73), .A1N(n2438), .Y(
        rdata2[18]) );
  OAI2BB2XL U766 ( .B0(n2436), .B1(n2193), .A0N(N72), .A1N(n2437), .Y(
        rdata2[19]) );
  OAI2BB2XL U767 ( .B0(n2436), .B1(n2190), .A0N(N71), .A1N(n2437), .Y(
        rdata2[20]) );
  OAI2BB2XL U768 ( .B0(n2436), .B1(n2187), .A0N(N70), .A1N(n2437), .Y(
        rdata2[21]) );
  OAI2BB2XL U769 ( .B0(n2436), .B1(n2184), .A0N(N69), .A1N(n2437), .Y(
        rdata2[22]) );
  OAI2BB2XL U770 ( .B0(n2436), .B1(n2181), .A0N(N68), .A1N(n2435), .Y(
        rdata2[23]) );
  OAI2BB2XL U771 ( .B0(n2436), .B1(n2178), .A0N(N67), .A1N(n2437), .Y(
        rdata2[24]) );
  OAI2BB2XL U772 ( .B0(n2436), .B1(n2175), .A0N(N66), .A1N(n2438), .Y(
        rdata2[25]) );
  OAI2BB2XL U773 ( .B0(n2436), .B1(n2172), .A0N(N65), .A1N(n2436), .Y(
        rdata2[26]) );
  OAI2BB2XL U774 ( .B0(n2435), .B1(n2169), .A0N(N64), .A1N(n2435), .Y(
        rdata2[27]) );
  OAI2BB2XL U775 ( .B0(n2435), .B1(n2166), .A0N(N63), .A1N(n2438), .Y(
        rdata2[28]) );
  OAI2BB2XL U776 ( .B0(n2435), .B1(n2163), .A0N(N62), .A1N(n2436), .Y(
        rdata2[29]) );
  OAI2BB2XL U777 ( .B0(n2435), .B1(n2160), .A0N(N61), .A1N(n2438), .Y(
        rdata2[30]) );
  OAI2BB2XL U778 ( .B0(n2435), .B1(n2157), .A0N(N60), .A1N(n2438), .Y(
        rdata2[31]) );
  OAI2BB2XL U779 ( .B0(n2249), .B1(n2432), .A0N(N56), .A1N(n2429), .Y(
        rdata1[0]) );
  OAI2BB2XL U780 ( .B0(n2246), .B1(n2431), .A0N(N55), .A1N(n2432), .Y(
        rdata1[1]) );
  OAI2BB2XL U781 ( .B0(n2235), .B1(n2430), .A0N(N51), .A1N(n2430), .Y(
        rdata1[5]) );
  OAI2BB2XL U782 ( .B0(n2232), .B1(n2430), .A0N(N50), .A1N(n2433), .Y(
        rdata1[6]) );
  OAI2BB2XL U783 ( .B0(n2229), .B1(n2430), .A0N(N49), .A1N(n2431), .Y(
        rdata1[7]) );
  OAI2BB2XL U784 ( .B0(n2226), .B1(n2430), .A0N(N48), .A1N(n2429), .Y(
        rdata1[8]) );
  OAI2BB2XL U785 ( .B0(n2223), .B1(n2431), .A0N(N47), .A1N(n2433), .Y(
        rdata1[9]) );
  OAI2BB2XL U786 ( .B0(n2220), .B1(n2432), .A0N(N46), .A1N(n2429), .Y(
        rdata1[10]) );
  OAI2BB2XL U787 ( .B0(n2217), .B1(n2432), .A0N(N45), .A1N(n2433), .Y(
        rdata1[11]) );
  OAI2BB2XL U788 ( .B0(n2214), .B1(n2432), .A0N(N44), .A1N(n2433), .Y(
        rdata1[12]) );
  OAI2BB2XL U789 ( .B0(n2211), .B1(n2432), .A0N(N43), .A1N(n2433), .Y(
        rdata1[13]) );
  OAI2BB2XL U790 ( .B0(n2208), .B1(n2432), .A0N(N42), .A1N(n2433), .Y(
        rdata1[14]) );
  OAI2BB2XL U791 ( .B0(n2205), .B1(n2432), .A0N(N41), .A1N(n2433), .Y(
        rdata1[15]) );
  OAI2BB2XL U792 ( .B0(n2202), .B1(n2431), .A0N(N40), .A1N(n2433), .Y(
        rdata1[16]) );
  OAI2BB2XL U793 ( .B0(n2199), .B1(n2432), .A0N(N39), .A1N(n2432), .Y(
        rdata1[17]) );
  OAI2BB2XL U794 ( .B0(n2190), .B1(n2431), .A0N(N36), .A1N(n2432), .Y(
        rdata1[20]) );
  OAI2BB2XL U795 ( .B0(n2187), .B1(n2431), .A0N(N35), .A1N(n2432), .Y(
        rdata1[21]) );
  OAI2BB2XL U796 ( .B0(n2184), .B1(n2431), .A0N(N34), .A1N(n2432), .Y(
        rdata1[22]) );
  OAI2BB2XL U797 ( .B0(n2181), .B1(n2431), .A0N(N33), .A1N(n2433), .Y(
        rdata1[23]) );
  NAND4X1 U798 ( .A(n48), .B(n49), .C(n50), .D(n51), .Y(n47) );
  XNOR2XL U799 ( .A(N18), .B(wsel[1]), .Y(n48) );
  NOR4X1 U800 ( .A(n52), .B(n2621), .C(n53), .D(n54), .Y(n51) );
  NAND4X1 U801 ( .A(n57), .B(n58), .C(n59), .D(n60), .Y(n56) );
  XNOR2XL U802 ( .A(N13), .B(wsel[1]), .Y(n57) );
  NOR4X1 U803 ( .A(n61), .B(n2621), .C(n62), .D(n63), .Y(n60) );
  MXI2X1 U804 ( .A(n1610), .B(n1611), .S0(n2090), .Y(N91) );
  MX4X1 U805 ( .A(n1677), .B(n1675), .C(n1676), .D(n1674), .S0(n2094), .S1(
        n2101), .Y(n1611) );
  MX4X1 U806 ( .A(n1681), .B(n1679), .C(n1680), .D(n1678), .S0(n2094), .S1(
        n2101), .Y(n1610) );
  MXI4X1 U807 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n2145), .S1(n2122), .Y(
        n1677) );
  MXI2X1 U808 ( .A(n1612), .B(n1613), .S0(n2090), .Y(N90) );
  MX4X1 U809 ( .A(n1689), .B(n1687), .C(n1688), .D(n1686), .S0(n2094), .S1(
        n2101), .Y(n1612) );
  MX4X1 U810 ( .A(n1685), .B(n1683), .C(n1684), .D(n1682), .S0(n2094), .S1(
        n2101), .Y(n1613) );
  MXI4X1 U811 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n2146), .S1(n2122), .Y(
        n1687) );
  MXI2X1 U812 ( .A(n1614), .B(n1615), .S0(n2090), .Y(N89) );
  MX4X1 U813 ( .A(n1697), .B(n1695), .C(n1696), .D(n1694), .S0(n2094), .S1(
        n2101), .Y(n1614) );
  MX4X1 U814 ( .A(n1693), .B(n1691), .C(n1692), .D(n1690), .S0(n2094), .S1(
        n2101), .Y(n1615) );
  MXI4X1 U815 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n2146), .S1(n2122), .Y(
        n1695) );
  MXI2X1 U816 ( .A(n1616), .B(n1617), .S0(n2090), .Y(N88) );
  MX4X1 U817 ( .A(n1705), .B(n1703), .C(n1704), .D(n1702), .S0(n2094), .S1(
        n2101), .Y(n1616) );
  MX4X1 U818 ( .A(n1701), .B(n1699), .C(n1700), .D(n1698), .S0(n2094), .S1(
        n2101), .Y(n1617) );
  MXI4X1 U819 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n2147), .S1(n2123), .Y(
        n1703) );
  MXI2X1 U820 ( .A(n1618), .B(n1619), .S0(n2090), .Y(N87) );
  MX4X1 U821 ( .A(n1713), .B(n1711), .C(n1712), .D(n1710), .S0(n2094), .S1(
        n2101), .Y(n1618) );
  MX4X1 U822 ( .A(n1709), .B(n1707), .C(n1708), .D(n1706), .S0(n2094), .S1(
        n2101), .Y(n1619) );
  MXI4X1 U823 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n2147), .S1(n2123), .Y(
        n1711) );
  MXI2X1 U824 ( .A(n1620), .B(n1621), .S0(n2090), .Y(N86) );
  MX4X1 U825 ( .A(n1717), .B(n1715), .C(n1716), .D(n1714), .S0(n2094), .S1(
        n2101), .Y(n1621) );
  MX4X1 U826 ( .A(n1721), .B(n1719), .C(n1720), .D(n1718), .S0(n2094), .S1(
        n2101), .Y(n1620) );
  MXI4X1 U827 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n2147), .S1(n2123), .Y(
        n1717) );
  MXI2X1 U828 ( .A(n1622), .B(n1623), .S0(n2090), .Y(N85) );
  MX4X1 U829 ( .A(n1729), .B(n1727), .C(n1728), .D(n1726), .S0(n2094), .S1(
        n2101), .Y(n1622) );
  MX4X1 U830 ( .A(n1725), .B(n1723), .C(n1724), .D(n1722), .S0(n2094), .S1(
        n2101), .Y(n1623) );
  MXI4X1 U831 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n2148), .S1(n2124), .Y(
        n1727) );
  MXI2X1 U832 ( .A(n1624), .B(n1625), .S0(n2090), .Y(N84) );
  MX4X1 U833 ( .A(n1733), .B(n1731), .C(n1732), .D(n1730), .S0(n2094), .S1(
        n2101), .Y(n1625) );
  MX4X1 U834 ( .A(n1737), .B(n1735), .C(n1736), .D(n1734), .S0(n2094), .S1(
        n2101), .Y(n1624) );
  MXI2X1 U835 ( .A(n1626), .B(n1627), .S0(n2091), .Y(N83) );
  MX4X1 U836 ( .A(n1741), .B(n1739), .C(n1740), .D(n1738), .S0(n2095), .S1(
        n2102), .Y(n1627) );
  MX4X1 U837 ( .A(n1745), .B(n1743), .C(n1744), .D(n1742), .S0(n2095), .S1(
        n2102), .Y(n1626) );
  MXI4X1 U838 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n2149), .S1(n2124), .Y(
        n1741) );
  MXI2X1 U839 ( .A(n1628), .B(n1629), .S0(n2091), .Y(N82) );
  MX4X1 U840 ( .A(n1749), .B(n1747), .C(n1748), .D(n1746), .S0(n2095), .S1(
        n2102), .Y(n1629) );
  MX4X1 U841 ( .A(n1753), .B(n1751), .C(n1752), .D(n1750), .S0(n2095), .S1(
        n2102), .Y(n1628) );
  MXI4X1 U842 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n2149), .S1(n2125), .Y(
        n1749) );
  MXI2X1 U843 ( .A(n1630), .B(n1631), .S0(n2091), .Y(N81) );
  MX4X1 U844 ( .A(n1757), .B(n1755), .C(n1756), .D(n1754), .S0(n2095), .S1(
        n2102), .Y(n1631) );
  MX4X1 U845 ( .A(n1761), .B(n1759), .C(n1760), .D(n1758), .S0(n2095), .S1(
        n2102), .Y(n1630) );
  MXI4X1 U846 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1757) );
  MXI2X1 U847 ( .A(n1632), .B(n1633), .S0(n2091), .Y(N80) );
  MX4X1 U848 ( .A(n1765), .B(n1763), .C(n1764), .D(n1762), .S0(n2095), .S1(
        n2102), .Y(n1633) );
  MX4X1 U849 ( .A(n1769), .B(n1767), .C(n1768), .D(n1766), .S0(n2095), .S1(
        n2102), .Y(n1632) );
  MXI4X1 U850 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1765) );
  MXI2X1 U851 ( .A(n1634), .B(n1635), .S0(n2091), .Y(N79) );
  MX4X1 U852 ( .A(n1777), .B(n1775), .C(n1776), .D(n1774), .S0(n2095), .S1(
        n2102), .Y(n1634) );
  MX4X1 U853 ( .A(n1773), .B(n1771), .C(n1772), .D(n1770), .S0(n2095), .S1(
        n2102), .Y(n1635) );
  MXI4X1 U854 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n2145), .S1(n2126), 
        .Y(n1775) );
  MXI2X1 U855 ( .A(n1636), .B(n1637), .S0(n2091), .Y(N78) );
  MX4X1 U856 ( .A(n1781), .B(n1779), .C(n1780), .D(n1778), .S0(n2095), .S1(
        n2102), .Y(n1637) );
  MX4X1 U857 ( .A(n1785), .B(n1783), .C(n1784), .D(n1782), .S0(n2095), .S1(
        n2102), .Y(n1636) );
  MXI4X1 U858 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n2145), .S1(n2126), 
        .Y(n1781) );
  MXI2X1 U859 ( .A(n1638), .B(n1639), .S0(n2091), .Y(N77) );
  MX4X1 U860 ( .A(n1789), .B(n1787), .C(n1788), .D(n1786), .S0(n2096), .S1(
        n2103), .Y(n1639) );
  MX4X1 U861 ( .A(n1793), .B(n1791), .C(n1792), .D(n1790), .S0(n2096), .S1(
        n2103), .Y(n1638) );
  MXI4X1 U862 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1789) );
  MXI2X1 U863 ( .A(n1640), .B(n1641), .S0(n2091), .Y(N76) );
  MX4X1 U864 ( .A(n1797), .B(n1795), .C(n1796), .D(n1794), .S0(n2096), .S1(
        n2103), .Y(n1641) );
  MX4X1 U865 ( .A(n1801), .B(n1799), .C(n1800), .D(n1798), .S0(n2096), .S1(
        n2103), .Y(n1640) );
  MXI2X1 U866 ( .A(n1642), .B(n1643), .S0(n2091), .Y(N75) );
  MX4X1 U867 ( .A(n1805), .B(n1803), .C(n1804), .D(n1802), .S0(n2096), .S1(
        n2103), .Y(n1643) );
  MX4X1 U868 ( .A(n1809), .B(n1807), .C(n1808), .D(n1806), .S0(n2096), .S1(
        n2103), .Y(n1642) );
  MXI4X1 U869 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1805) );
  MXI2X1 U870 ( .A(n1644), .B(n1645), .S0(n2091), .Y(N74) );
  MX4X1 U871 ( .A(n1813), .B(n1811), .C(n1812), .D(n1810), .S0(n2096), .S1(
        n2103), .Y(n1645) );
  MX4X1 U872 ( .A(n1817), .B(n1815), .C(n1816), .D(n1814), .S0(n2096), .S1(
        n2103), .Y(n1644) );
  MXI4X1 U873 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1813) );
  MXI2X1 U874 ( .A(n1646), .B(n1647), .S0(n2091), .Y(N73) );
  MX4X1 U875 ( .A(n1821), .B(n1819), .C(n1820), .D(n1818), .S0(n2096), .S1(
        n2103), .Y(n1647) );
  MX4X1 U876 ( .A(n1825), .B(n1823), .C(n1824), .D(n1822), .S0(n2096), .S1(
        n2103), .Y(n1646) );
  MXI4X1 U877 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n2142), .S1(n2117), 
        .Y(n1821) );
  MXI2X1 U879 ( .A(n1648), .B(n1649), .S0(n2091), .Y(N72) );
  MX4X1 U880 ( .A(n1829), .B(n1827), .C(n1828), .D(n1826), .S0(n2096), .S1(
        n2103), .Y(n1649) );
  MX4X1 U881 ( .A(n1833), .B(n1831), .C(n1832), .D(n1830), .S0(n2096), .S1(
        n2103), .Y(n1648) );
  MXI4X1 U882 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n2142), .S1(n2118), 
        .Y(n1829) );
  MXI2X1 U883 ( .A(n1650), .B(n1651), .S0(n2092), .Y(N71) );
  MX4X1 U884 ( .A(n1837), .B(n1835), .C(n1836), .D(n1834), .S0(n2097), .S1(
        n2104), .Y(n1651) );
  MX4X1 U885 ( .A(n1841), .B(n1839), .C(n1840), .D(n1838), .S0(n2097), .S1(
        n2104), .Y(n1650) );
  MXI2X1 U886 ( .A(n1652), .B(n1653), .S0(n2092), .Y(N70) );
  MX4X1 U887 ( .A(n1845), .B(n1843), .C(n1844), .D(n1842), .S0(n2097), .S1(
        n2104), .Y(n1653) );
  MX4X1 U888 ( .A(n1849), .B(n1847), .C(n1848), .D(n1846), .S0(n2097), .S1(
        n2104), .Y(n1652) );
  MXI4X1 U889 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1845) );
  MXI2X1 U890 ( .A(n1654), .B(n1655), .S0(n2092), .Y(N69) );
  MX4X1 U891 ( .A(n1853), .B(n1851), .C(n1852), .D(n1850), .S0(n2097), .S1(
        n2104), .Y(n1655) );
  MX4X1 U892 ( .A(n1857), .B(n1855), .C(n1856), .D(n1854), .S0(n2097), .S1(
        n2104), .Y(n1654) );
  MXI4X1 U893 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n2145), .S1(n2119), 
        .Y(n1853) );
  MXI2X1 U894 ( .A(n1656), .B(n1657), .S0(n2092), .Y(N68) );
  MX4X1 U895 ( .A(n1861), .B(n1859), .C(n1860), .D(n1858), .S0(n2097), .S1(
        n2104), .Y(n1657) );
  MX4X1 U896 ( .A(n1865), .B(n1863), .C(n1864), .D(n1862), .S0(n2097), .S1(
        n2104), .Y(n1656) );
  MXI4X1 U897 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1861) );
  MXI2X1 U898 ( .A(n1658), .B(n1659), .S0(n2092), .Y(N67) );
  MX4X1 U899 ( .A(n1869), .B(n1867), .C(n1868), .D(n1866), .S0(n2097), .S1(
        n2104), .Y(n1659) );
  MX4X1 U900 ( .A(n1873), .B(n1871), .C(n1872), .D(n1870), .S0(n2097), .S1(
        n2104), .Y(n1658) );
  MXI4X1 U901 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n2143), .S1(n2119), 
        .Y(n1869) );
  MXI2X1 U902 ( .A(n1660), .B(n1661), .S0(n2092), .Y(N66) );
  MX4X1 U903 ( .A(n1877), .B(n1875), .C(n1876), .D(n1874), .S0(n2097), .S1(
        n2104), .Y(n1661) );
  MX4X1 U904 ( .A(n1881), .B(n1879), .C(n1880), .D(n1878), .S0(n2097), .S1(
        n2104), .Y(n1660) );
  MXI4X1 U905 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n2143), .S1(n2120), 
        .Y(n1877) );
  MXI2X1 U906 ( .A(n1662), .B(n1663), .S0(n2092), .Y(N65) );
  MX4X1 U907 ( .A(n1885), .B(n1883), .C(n1884), .D(n1882), .S0(n2098), .S1(
        n2105), .Y(n1663) );
  MX4X1 U908 ( .A(n1889), .B(n1887), .C(n1888), .D(n1886), .S0(n2098), .S1(
        n2105), .Y(n1662) );
  MXI4X1 U909 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n2143), .S1(n2120), 
        .Y(n1885) );
  MXI2X1 U910 ( .A(n1664), .B(n1665), .S0(n2092), .Y(N64) );
  MX4X1 U911 ( .A(n1893), .B(n1891), .C(n1892), .D(n1890), .S0(n2098), .S1(
        n2105), .Y(n1665) );
  MX4X1 U912 ( .A(n1897), .B(n1895), .C(n1896), .D(n1894), .S0(n2098), .S1(
        n2105), .Y(n1664) );
  MXI4X1 U913 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1893) );
  MXI2X1 U914 ( .A(n1666), .B(n1667), .S0(n2092), .Y(N63) );
  MX4X1 U915 ( .A(n1901), .B(n1899), .C(n1900), .D(n1898), .S0(n2098), .S1(
        n2105), .Y(n1667) );
  MX4X1 U916 ( .A(n1905), .B(n1903), .C(n1904), .D(n1902), .S0(n2098), .S1(
        n2105), .Y(n1666) );
  MXI4X1 U917 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n2144), .S1(n2121), 
        .Y(n1901) );
  MXI2X1 U918 ( .A(n1668), .B(n1669), .S0(n2092), .Y(N62) );
  MX4X1 U919 ( .A(n1909), .B(n1907), .C(n1908), .D(n1906), .S0(n2098), .S1(
        n2105), .Y(n1669) );
  MX4X1 U920 ( .A(n1913), .B(n1911), .C(n1912), .D(n1910), .S0(n2098), .S1(
        n2105), .Y(n1668) );
  MXI4X1 U921 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1909) );
  MXI2X1 U922 ( .A(n1670), .B(n1671), .S0(n2092), .Y(N61) );
  MX4X1 U923 ( .A(n1917), .B(n1915), .C(n1916), .D(n1914), .S0(n2098), .S1(
        n2105), .Y(n1671) );
  MX4X1 U924 ( .A(n1921), .B(n1919), .C(n1920), .D(n1918), .S0(n2098), .S1(
        n2105), .Y(n1670) );
  MXI4X1 U925 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1917) );
  MXI2X1 U926 ( .A(n1672), .B(n1673), .S0(n2092), .Y(N60) );
  MX4X1 U927 ( .A(n1925), .B(n1923), .C(n1924), .D(n1922), .S0(n2098), .S1(
        n2105), .Y(n1673) );
  MX4X1 U928 ( .A(n1929), .B(n1927), .C(n1928), .D(n1926), .S0(n2098), .S1(
        n2105), .Y(n1672) );
  MXI4X1 U929 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n2145), .S1(n2121), 
        .Y(n1925) );
  MXI2X1 U930 ( .A(n17), .B(n18), .S0(n1546), .Y(N56) );
  MX4X1 U931 ( .A(n1133), .B(n1131), .C(n1132), .D(n1130), .S0(n1552), .S1(
        n1561), .Y(n18) );
  MX4X1 U932 ( .A(n1137), .B(n1135), .C(n1136), .D(n1134), .S0(n1552), .S1(
        n1561), .Y(n17) );
  MXI4X1 U933 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1599), .S1(n1578), .Y(
        n1133) );
  MXI2X1 U934 ( .A(n19), .B(n20), .S0(n1546), .Y(N55) );
  MX4X1 U935 ( .A(n1145), .B(n1143), .C(n1144), .D(n1142), .S0(n1552), .S1(
        n1561), .Y(n19) );
  MX4X1 U936 ( .A(n1141), .B(n1139), .C(n1140), .D(n1138), .S0(n1552), .S1(
        n1561), .Y(n20) );
  MXI2X1 U937 ( .A(n21), .B(n22), .S0(n1546), .Y(N54) );
  MX4X1 U938 ( .A(n1153), .B(n1151), .C(n1152), .D(n1150), .S0(n1553), .S1(
        n1561), .Y(n21) );
  MX4X1 U939 ( .A(n1149), .B(n1147), .C(n1148), .D(n1146), .S0(n1553), .S1(
        n1561), .Y(n22) );
  MXI4X1 U940 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1600), .S1(n1578), .Y(
        n1151) );
  MXI2X1 U941 ( .A(n23), .B(n24), .S0(n1546), .Y(N53) );
  MX4X1 U942 ( .A(n1161), .B(n1159), .C(n1160), .D(n1158), .S0(n1553), .S1(
        n1561), .Y(n23) );
  MX4X1 U943 ( .A(n1157), .B(n1155), .C(n1156), .D(n1154), .S0(n1553), .S1(
        n1561), .Y(n24) );
  MXI4X1 U944 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1601), .S1(n1579), .Y(
        n1159) );
  MXI2X1 U945 ( .A(n25), .B(n26), .S0(n1546), .Y(N52) );
  MX4X1 U946 ( .A(n1169), .B(n1167), .C(n1168), .D(n1166), .S0(n1553), .S1(
        n1561), .Y(n25) );
  MX4X1 U947 ( .A(n1165), .B(n1163), .C(n1164), .D(n1162), .S0(n1553), .S1(
        n1561), .Y(n26) );
  MXI4X1 U948 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1601), .S1(n1579), .Y(
        n1167) );
  MXI2X1 U949 ( .A(n27), .B(n28), .S0(n1546), .Y(N51) );
  MX4X1 U950 ( .A(n1173), .B(n1171), .C(n1172), .D(n1170), .S0(n1553), .S1(
        n1561), .Y(n28) );
  MX4X1 U951 ( .A(n1177), .B(n1175), .C(n1176), .D(n1174), .S0(n1553), .S1(
        n1561), .Y(n27) );
  MXI4X1 U952 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1601), .S1(n1579), .Y(
        n1173) );
  MXI2X1 U953 ( .A(n29), .B(n30), .S0(n1546), .Y(N50) );
  MX4X1 U954 ( .A(n1185), .B(n1183), .C(n1184), .D(n1182), .S0(n1553), .S1(
        n1561), .Y(n29) );
  MX4X1 U955 ( .A(n1181), .B(n1179), .C(n1180), .D(n1178), .S0(n1553), .S1(
        n1561), .Y(n30) );
  MXI4X1 U956 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1602), .S1(n1580), .Y(
        n1183) );
  MXI2X1 U957 ( .A(n31), .B(n32), .S0(n1546), .Y(N49) );
  MX4X1 U958 ( .A(n1189), .B(n1187), .C(n1188), .D(n1186), .S0(n1553), .S1(
        n1561), .Y(n32) );
  MX4X1 U959 ( .A(n1193), .B(n1191), .C(n1192), .D(n1190), .S0(n1553), .S1(
        n1561), .Y(n31) );
  MXI4X1 U960 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1602), .S1(n1580), .Y(
        n1189) );
  MXI2X1 U961 ( .A(n33), .B(n34), .S0(n1547), .Y(N48) );
  MX4X1 U962 ( .A(n1197), .B(n1195), .C(n1196), .D(n1194), .S0(n1554), .S1(
        n1562), .Y(n34) );
  MX4X1 U963 ( .A(n1201), .B(n1199), .C(n1200), .D(n1198), .S0(n1554), .S1(
        n1562), .Y(n33) );
  MXI4X1 U964 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1603), .S1(n1580), .Y(
        n1197) );
  MXI2X1 U965 ( .A(n35), .B(n36), .S0(n1547), .Y(N47) );
  MX4X1 U966 ( .A(n1205), .B(n1203), .C(n1204), .D(n1202), .S0(n1554), .S1(
        n1562), .Y(n36) );
  MX4X1 U967 ( .A(n1209), .B(n1207), .C(n1208), .D(n1206), .S0(n1554), .S1(
        n1562), .Y(n35) );
  MXI4X1 U968 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1603), .S1(n1581), .Y(
        n1205) );
  MXI2X1 U969 ( .A(n37), .B(n38), .S0(n1547), .Y(N46) );
  MX4X1 U970 ( .A(n1213), .B(n1211), .C(n1212), .D(n1210), .S0(n1554), .S1(
        n1562), .Y(n38) );
  MX4X1 U971 ( .A(n1217), .B(n1215), .C(n1216), .D(n1214), .S0(n1554), .S1(
        n1562), .Y(n37) );
  MXI4X1 U972 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1213) );
  MXI2X1 U973 ( .A(n39), .B(n40), .S0(n1547), .Y(N45) );
  MX4X1 U974 ( .A(n1221), .B(n1219), .C(n1220), .D(n1218), .S0(n1554), .S1(
        n1562), .Y(n40) );
  MX4X1 U975 ( .A(n1225), .B(n1223), .C(n1224), .D(n1222), .S0(n1554), .S1(
        n1562), .Y(n39) );
  MXI4X1 U976 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1221) );
  MXI2X1 U977 ( .A(n41), .B(n42), .S0(n1547), .Y(N44) );
  MX4X1 U978 ( .A(n1233), .B(n1231), .C(n1232), .D(n1230), .S0(n1554), .S1(
        n1562), .Y(n41) );
  MX4X1 U979 ( .A(n1229), .B(n1227), .C(n1228), .D(n1226), .S0(n1554), .S1(
        n1562), .Y(n42) );
  MXI4X1 U980 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1605), .S1(n1582), 
        .Y(n1231) );
  MXI2X1 U981 ( .A(n43), .B(n44), .S0(n1547), .Y(N43) );
  MX4X1 U982 ( .A(n1237), .B(n1235), .C(n1236), .D(n1234), .S0(n1554), .S1(
        n1562), .Y(n44) );
  MX4X1 U983 ( .A(n1241), .B(n1239), .C(n1240), .D(n1238), .S0(n1554), .S1(
        n1562), .Y(n43) );
  MXI4X1 U984 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1237) );
  MXI2X1 U985 ( .A(n45), .B(n46), .S0(n1547), .Y(N42) );
  MX4X1 U986 ( .A(n1245), .B(n1243), .C(n1244), .D(n1242), .S0(n1555), .S1(
        n1563), .Y(n46) );
  MX4X1 U987 ( .A(n1249), .B(n1247), .C(n1248), .D(n1246), .S0(n1555), .S1(
        n1563), .Y(n45) );
  MXI2X1 U988 ( .A(n66), .B(n73), .S0(n1547), .Y(N41) );
  MX4X1 U989 ( .A(n1253), .B(n1251), .C(n1252), .D(n1250), .S0(n1555), .S1(
        n1563), .Y(n73) );
  MX4X1 U990 ( .A(n1257), .B(n1255), .C(n1256), .D(n1254), .S0(n1555), .S1(
        n1563), .Y(n66) );
  MXI4X1 U991 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1606), .S1(n1582), 
        .Y(n1253) );
  MXI2X1 U992 ( .A(n75), .B(n82), .S0(n1547), .Y(N40) );
  MX4X1 U993 ( .A(n1261), .B(n1259), .C(n1260), .D(n1258), .S0(n1555), .S1(
        n1563), .Y(n82) );
  MX4X1 U994 ( .A(n1265), .B(n1263), .C(n1264), .D(n1262), .S0(n1555), .S1(
        n1563), .Y(n75) );
  MXI4X1 U995 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1261) );
  MXI2X1 U996 ( .A(n1100), .B(n1101), .S0(n1547), .Y(N39) );
  MX4X1 U997 ( .A(n1269), .B(n1267), .C(n1268), .D(n1266), .S0(n1555), .S1(
        n1563), .Y(n1101) );
  MX4X1 U998 ( .A(n1273), .B(n1271), .C(n1272), .D(n1270), .S0(n1555), .S1(
        n1563), .Y(n1100) );
  MXI4X1 U999 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1269) );
  MXI2X1 U1000 ( .A(n1102), .B(n1103), .S0(n1547), .Y(N38) );
  MX4X1 U1001 ( .A(n1277), .B(n1275), .C(n1276), .D(n1274), .S0(n1555), .S1(
        n1563), .Y(n1103) );
  MX4X1 U1002 ( .A(n1281), .B(n1279), .C(n1280), .D(n1278), .S0(n1555), .S1(
        n1563), .Y(n1102) );
  MXI4X1 U1003 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1599), .S1(n1573), 
        .Y(n1277) );
  MXI2X1 U1004 ( .A(n1104), .B(n1105), .S0(n1547), .Y(N37) );
  MX4X1 U1005 ( .A(n1285), .B(n1283), .C(n1284), .D(n1282), .S0(n1555), .S1(
        n1563), .Y(n1105) );
  MX4X1 U1006 ( .A(n1289), .B(n1287), .C(n1288), .D(n1286), .S0(n1555), .S1(
        n1563), .Y(n1104) );
  MXI4X1 U1007 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1599), .S1(n1574), 
        .Y(n1285) );
  MXI2X1 U1008 ( .A(n1106), .B(n1107), .S0(n1548), .Y(N36) );
  MX4X1 U1009 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1556), .S1(
        n1564), .Y(n1107) );
  MX4X1 U1010 ( .A(n1297), .B(n1295), .C(n1296), .D(n1294), .S0(n1556), .S1(
        n1564), .Y(n1106) );
  MXI4X1 U1011 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1293) );
  MXI2X1 U1012 ( .A(n1108), .B(n1109), .S0(n1548), .Y(N35) );
  MX4X1 U1013 ( .A(n1301), .B(n1299), .C(n1300), .D(n1298), .S0(n1556), .S1(
        n1564), .Y(n1109) );
  MX4X1 U1014 ( .A(n1305), .B(n1303), .C(n1304), .D(n1302), .S0(n1556), .S1(
        n1564), .Y(n1108) );
  MXI4X1 U1015 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1599), .S1(n1574), 
        .Y(n1301) );
  MXI2X1 U1016 ( .A(n1110), .B(n1111), .S0(n1548), .Y(N34) );
  MX4X1 U1017 ( .A(n1309), .B(n1307), .C(n1308), .D(n1306), .S0(n1556), .S1(
        n1564), .Y(n1111) );
  MX4X1 U1018 ( .A(n1313), .B(n1311), .C(n1312), .D(n1310), .S0(n1556), .S1(
        n1564), .Y(n1110) );
  MXI4X1 U1019 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1596), .S1(n1575), 
        .Y(n1309) );
  MXI2X1 U1020 ( .A(n1112), .B(n1113), .S0(n1548), .Y(N33) );
  MX4X1 U1021 ( .A(n1317), .B(n1315), .C(n1316), .D(n1314), .S0(n1556), .S1(
        n1564), .Y(n1113) );
  MX4X1 U1022 ( .A(n1321), .B(n1319), .C(n1320), .D(n1318), .S0(n1556), .S1(
        n1564), .Y(n1112) );
  MXI4X1 U1023 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1317) );
  MXI2X1 U1024 ( .A(n1114), .B(n1115), .S0(n1548), .Y(N32) );
  MX4X1 U1025 ( .A(n1325), .B(n1323), .C(n1324), .D(n1322), .S0(n1556), .S1(
        n1564), .Y(n1115) );
  MX4X1 U1026 ( .A(n1329), .B(n1327), .C(n1328), .D(n1326), .S0(n1556), .S1(
        n1564), .Y(n1114) );
  MXI4X1 U1027 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1597), .S1(n1575), 
        .Y(n1325) );
  MXI2X1 U1028 ( .A(n1116), .B(n1117), .S0(n1548), .Y(N31) );
  MX4X1 U1029 ( .A(n1333), .B(n1331), .C(n1332), .D(n1330), .S0(n1556), .S1(
        n1564), .Y(n1117) );
  MX4X1 U1030 ( .A(n1337), .B(n1335), .C(n1336), .D(n1334), .S0(n1556), .S1(
        n1564), .Y(n1116) );
  MXI4X1 U1031 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1597), .S1(n1576), 
        .Y(n1333) );
  MXI2X1 U1032 ( .A(n1118), .B(n1119), .S0(n1548), .Y(N30) );
  MX4X1 U1033 ( .A(n1341), .B(n1339), .C(n1340), .D(n1338), .S0(n1557), .S1(
        n1565), .Y(n1119) );
  MX4X1 U1034 ( .A(n1345), .B(n1343), .C(n1344), .D(n1342), .S0(n1557), .S1(
        n1565), .Y(n1118) );
  MXI4X1 U1035 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1597), .S1(n1576), 
        .Y(n1341) );
  MXI2X1 U1036 ( .A(n1120), .B(n1121), .S0(n1548), .Y(N29) );
  MX4X1 U1037 ( .A(n1349), .B(n1347), .C(n1348), .D(n1346), .S0(n1557), .S1(
        n1565), .Y(n1121) );
  MX4X1 U1038 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1557), .S1(
        n1565), .Y(n1120) );
  MXI4X1 U1039 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1349) );
  MXI2X1 U1040 ( .A(n1122), .B(n1123), .S0(n1548), .Y(N28) );
  MX4X1 U1041 ( .A(n1357), .B(n1355), .C(n1356), .D(n1354), .S0(n1557), .S1(
        n1565), .Y(n1123) );
  MX4X1 U1042 ( .A(n1361), .B(n1359), .C(n1360), .D(n1358), .S0(n1557), .S1(
        n1565), .Y(n1122) );
  MXI4X1 U1043 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1598), .S1(n1577), 
        .Y(n1357) );
  MXI2X1 U1044 ( .A(n1124), .B(n1125), .S0(n1548), .Y(N27) );
  MX4X1 U1045 ( .A(n1365), .B(n1363), .C(n1364), .D(n1362), .S0(n1557), .S1(
        n1565), .Y(n1125) );
  MX4X1 U1046 ( .A(n1369), .B(n1367), .C(n1368), .D(n1366), .S0(n1557), .S1(
        n1565), .Y(n1124) );
  MXI4X1 U1047 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1599), .S1(n1577), 
        .Y(n1365) );
  MXI2X1 U1048 ( .A(n1126), .B(n1127), .S0(n1548), .Y(N26) );
  MX4X1 U1049 ( .A(n1373), .B(n1371), .C(n1372), .D(n1370), .S0(n1557), .S1(
        n1565), .Y(n1127) );
  MX4X1 U1050 ( .A(n1377), .B(n1375), .C(n1376), .D(n1374), .S0(n1557), .S1(
        n1565), .Y(n1126) );
  MXI4X1 U1051 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1599), .S1(n1577), 
        .Y(n1373) );
  MXI2X1 U1052 ( .A(n1128), .B(n1129), .S0(n1548), .Y(N25) );
  MX4X1 U1053 ( .A(n1381), .B(n1379), .C(n1380), .D(n1378), .S0(n1557), .S1(
        n1565), .Y(n1129) );
  MX4X1 U1054 ( .A(n1385), .B(n1383), .C(n1384), .D(n1382), .S0(n1557), .S1(
        n1565), .Y(n1128) );
  MXI4X1 U1055 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1599), .S1(n1577), 
        .Y(n1381) );
  OAI2BB2XL U1056 ( .B0(n2181), .B1(n2421), .A0N(\register[2][23] ), .A1N(
        n2421), .Y(n163) );
  OAI2BB2XL U1057 ( .B0(n2175), .B1(n2421), .A0N(\register[2][25] ), .A1N(
        n2422), .Y(n165) );
  OAI2BB2XL U1058 ( .B0(n2172), .B1(n2421), .A0N(\register[2][26] ), .A1N(
        n2422), .Y(n166) );
  OAI2BB2XL U1059 ( .B0(n2169), .B1(n2421), .A0N(\register[2][27] ), .A1N(
        n2422), .Y(n167) );
  OAI2BB2XL U1060 ( .B0(n2166), .B1(n2421), .A0N(\register[2][28] ), .A1N(
        n2422), .Y(n168) );
  OAI2BB2XL U1061 ( .B0(n2163), .B1(n2421), .A0N(\register[2][29] ), .A1N(
        n2422), .Y(n169) );
  OAI2BB2XL U1062 ( .B0(n2160), .B1(n2421), .A0N(\register[2][30] ), .A1N(
        n2417), .Y(n170) );
  OAI2BB2XL U1063 ( .B0(n2157), .B1(n2421), .A0N(\register[2][31] ), .A1N(
        n2417), .Y(n171) );
  OAI2BB2XL U1064 ( .B0(n2181), .B1(n2414), .A0N(\register[3][23] ), .A1N(
        n2414), .Y(n195) );
  OAI2BB2XL U1065 ( .B0(n2175), .B1(n2414), .A0N(\register[3][25] ), .A1N(
        n2415), .Y(n197) );
  OAI2BB2XL U1066 ( .B0(n2172), .B1(n2414), .A0N(\register[3][26] ), .A1N(
        n2415), .Y(n198) );
  OAI2BB2XL U1067 ( .B0(n2169), .B1(n2414), .A0N(\register[3][27] ), .A1N(
        n2415), .Y(n199) );
  OAI2BB2XL U1068 ( .B0(n2166), .B1(n2414), .A0N(\register[3][28] ), .A1N(
        n2415), .Y(n200) );
  OAI2BB2XL U1069 ( .B0(n2163), .B1(n2414), .A0N(\register[3][29] ), .A1N(
        n2415), .Y(n201) );
  OAI2BB2XL U1070 ( .B0(n2160), .B1(n2414), .A0N(\register[3][30] ), .A1N(
        n2416), .Y(n202) );
  OAI2BB2XL U1071 ( .B0(n2157), .B1(n2414), .A0N(\register[3][31] ), .A1N(
        n2416), .Y(n203) );
  OAI2BB2XL U1072 ( .B0(n2180), .B1(n2374), .A0N(\register[10][23] ), .A1N(
        n2374), .Y(n419) );
  OAI2BB2XL U1073 ( .B0(n2174), .B1(n2374), .A0N(\register[10][25] ), .A1N(
        n2375), .Y(n421) );
  OAI2BB2XL U1074 ( .B0(n2171), .B1(n2374), .A0N(\register[10][26] ), .A1N(
        n2375), .Y(n422) );
  OAI2BB2XL U1075 ( .B0(n2168), .B1(n2374), .A0N(\register[10][27] ), .A1N(
        n2375), .Y(n423) );
  OAI2BB2XL U1076 ( .B0(n2165), .B1(n2374), .A0N(\register[10][28] ), .A1N(
        n2375), .Y(n424) );
  OAI2BB2XL U1077 ( .B0(n2162), .B1(n2374), .A0N(\register[10][29] ), .A1N(
        n2375), .Y(n425) );
  OAI2BB2XL U1078 ( .B0(n2159), .B1(n2374), .A0N(\register[10][30] ), .A1N(
        n2370), .Y(n426) );
  OAI2BB2XL U1079 ( .B0(n2156), .B1(n2374), .A0N(\register[10][31] ), .A1N(
        n2370), .Y(n427) );
  OAI2BB2XL U1080 ( .B0(n2180), .B1(n2368), .A0N(\register[11][23] ), .A1N(
        n2368), .Y(n451) );
  OAI2BB2XL U1081 ( .B0(n2174), .B1(n2368), .A0N(\register[11][25] ), .A1N(
        n2369), .Y(n453) );
  OAI2BB2XL U1082 ( .B0(n2171), .B1(n2368), .A0N(\register[11][26] ), .A1N(
        n2369), .Y(n454) );
  OAI2BB2XL U1083 ( .B0(n2168), .B1(n2368), .A0N(\register[11][27] ), .A1N(
        n2369), .Y(n455) );
  OAI2BB2XL U1084 ( .B0(n2165), .B1(n2368), .A0N(\register[11][28] ), .A1N(
        n2369), .Y(n456) );
  OAI2BB2XL U1085 ( .B0(n2162), .B1(n2368), .A0N(\register[11][29] ), .A1N(
        n2369), .Y(n457) );
  OAI2BB2XL U1086 ( .B0(n2159), .B1(n2368), .A0N(\register[11][30] ), .A1N(
        n2364), .Y(n458) );
  OAI2BB2XL U1087 ( .B0(n2156), .B1(n2368), .A0N(\register[11][31] ), .A1N(
        n2364), .Y(n459) );
  OAI2BB2XL U1088 ( .B0(n2180), .B1(n2330), .A0N(\register[18][23] ), .A1N(
        n2330), .Y(n675) );
  OAI2BB2XL U1089 ( .B0(n2174), .B1(n2330), .A0N(\register[18][25] ), .A1N(
        n2331), .Y(n677) );
  OAI2BB2XL U1090 ( .B0(n2171), .B1(n2330), .A0N(\register[18][26] ), .A1N(
        n2331), .Y(n678) );
  OAI2BB2XL U1091 ( .B0(n2168), .B1(n2330), .A0N(\register[18][27] ), .A1N(
        n2331), .Y(n679) );
  OAI2BB2XL U1092 ( .B0(n2165), .B1(n2330), .A0N(\register[18][28] ), .A1N(
        n2331), .Y(n680) );
  OAI2BB2XL U1093 ( .B0(n2162), .B1(n2330), .A0N(\register[18][29] ), .A1N(
        n2331), .Y(n681) );
  OAI2BB2XL U1094 ( .B0(n2159), .B1(n2330), .A0N(\register[18][30] ), .A1N(
        n2326), .Y(n682) );
  OAI2BB2XL U1095 ( .B0(n2156), .B1(n2330), .A0N(\register[18][31] ), .A1N(
        n2326), .Y(n683) );
  OAI2BB2XL U1096 ( .B0(n2180), .B1(n2324), .A0N(\register[19][23] ), .A1N(
        n2324), .Y(n707) );
  OAI2BB2XL U1097 ( .B0(n2174), .B1(n2324), .A0N(\register[19][25] ), .A1N(
        n2325), .Y(n709) );
  OAI2BB2XL U1098 ( .B0(n2171), .B1(n2324), .A0N(\register[19][26] ), .A1N(
        n2325), .Y(n710) );
  OAI2BB2XL U1099 ( .B0(n2168), .B1(n2324), .A0N(\register[19][27] ), .A1N(
        n2325), .Y(n711) );
  OAI2BB2XL U1100 ( .B0(n2165), .B1(n2324), .A0N(\register[19][28] ), .A1N(
        n2325), .Y(n712) );
  OAI2BB2XL U1101 ( .B0(n2162), .B1(n2324), .A0N(\register[19][29] ), .A1N(
        n2325), .Y(n713) );
  OAI2BB2XL U1102 ( .B0(n2159), .B1(n2324), .A0N(\register[19][30] ), .A1N(
        n2320), .Y(n714) );
  OAI2BB2XL U1103 ( .B0(n2156), .B1(n2324), .A0N(\register[19][31] ), .A1N(
        n2320), .Y(n715) );
  OAI2BB2XL U1104 ( .B0(n2179), .B1(n2282), .A0N(\register[26][23] ), .A1N(
        n2282), .Y(n931) );
  OAI2BB2XL U1105 ( .B0(n2173), .B1(n2282), .A0N(\register[26][25] ), .A1N(
        n2283), .Y(n933) );
  OAI2BB2XL U1106 ( .B0(n2170), .B1(n2282), .A0N(\register[26][26] ), .A1N(
        n2283), .Y(n934) );
  OAI2BB2XL U1107 ( .B0(n2167), .B1(n2282), .A0N(\register[26][27] ), .A1N(
        n2283), .Y(n935) );
  OAI2BB2XL U1108 ( .B0(n2164), .B1(n2282), .A0N(\register[26][28] ), .A1N(
        n2283), .Y(n936) );
  OAI2BB2XL U1109 ( .B0(n2161), .B1(n2282), .A0N(\register[26][29] ), .A1N(
        n2283), .Y(n937) );
  OAI2BB2XL U1110 ( .B0(n2158), .B1(n2282), .A0N(\register[26][30] ), .A1N(
        n2278), .Y(n938) );
  OAI2BB2XL U1111 ( .B0(n2155), .B1(n2282), .A0N(\register[26][31] ), .A1N(
        n2278), .Y(n939) );
  OAI2BB2XL U1112 ( .B0(n2179), .B1(n2276), .A0N(\register[27][23] ), .A1N(
        n2276), .Y(n963) );
  OAI2BB2XL U1113 ( .B0(n2173), .B1(n2276), .A0N(\register[27][25] ), .A1N(
        n2277), .Y(n965) );
  OAI2BB2XL U1114 ( .B0(n2170), .B1(n2276), .A0N(\register[27][26] ), .A1N(
        n2277), .Y(n966) );
  OAI2BB2XL U1115 ( .B0(n2167), .B1(n2276), .A0N(\register[27][27] ), .A1N(
        n2277), .Y(n967) );
  OAI2BB2XL U1116 ( .B0(n2164), .B1(n2276), .A0N(\register[27][28] ), .A1N(
        n2277), .Y(n968) );
  OAI2BB2XL U1117 ( .B0(n2161), .B1(n2276), .A0N(\register[27][29] ), .A1N(
        n2277), .Y(n969) );
  OAI2BB2XL U1118 ( .B0(n2158), .B1(n2276), .A0N(\register[27][30] ), .A1N(
        n2272), .Y(n970) );
  OAI2BB2XL U1119 ( .B0(n2155), .B1(n2276), .A0N(\register[27][31] ), .A1N(
        n2272), .Y(n971) );
  OAI2BB2XL U1120 ( .B0(n2181), .B1(n2427), .A0N(\register[1][23] ), .A1N(
        n2427), .Y(n131) );
  OAI2BB2XL U1121 ( .B0(n2175), .B1(n2427), .A0N(\register[1][25] ), .A1N(
        n2428), .Y(n133) );
  OAI2BB2XL U1122 ( .B0(n2172), .B1(n2427), .A0N(\register[1][26] ), .A1N(
        n2428), .Y(n134) );
  OAI2BB2XL U1123 ( .B0(n2169), .B1(n2427), .A0N(\register[1][27] ), .A1N(
        n2428), .Y(n135) );
  OAI2BB2XL U1124 ( .B0(n2166), .B1(n2427), .A0N(\register[1][28] ), .A1N(
        n2428), .Y(n136) );
  OAI2BB2XL U1125 ( .B0(n2163), .B1(n2427), .A0N(\register[1][29] ), .A1N(
        n2428), .Y(n137) );
  OAI2BB2XL U1126 ( .B0(n2160), .B1(n2427), .A0N(\register[1][30] ), .A1N(
        n2423), .Y(n138) );
  OAI2BB2XL U1127 ( .B0(n2157), .B1(n2427), .A0N(\register[1][31] ), .A1N(
        n2423), .Y(n139) );
  OAI2BB2XL U1128 ( .B0(n2180), .B1(n2380), .A0N(\register[9][23] ), .A1N(
        n2380), .Y(n387) );
  OAI2BB2XL U1129 ( .B0(n2174), .B1(n2380), .A0N(\register[9][25] ), .A1N(
        n2381), .Y(n389) );
  OAI2BB2XL U1130 ( .B0(n2171), .B1(n2380), .A0N(\register[9][26] ), .A1N(
        n2381), .Y(n390) );
  OAI2BB2XL U1131 ( .B0(n2168), .B1(n2380), .A0N(\register[9][27] ), .A1N(
        n2381), .Y(n391) );
  OAI2BB2XL U1132 ( .B0(n2165), .B1(n2380), .A0N(\register[9][28] ), .A1N(
        n2381), .Y(n392) );
  OAI2BB2XL U1133 ( .B0(n2162), .B1(n2380), .A0N(\register[9][29] ), .A1N(
        n2381), .Y(n393) );
  OAI2BB2XL U1134 ( .B0(n2159), .B1(n2380), .A0N(\register[9][30] ), .A1N(
        n2376), .Y(n394) );
  OAI2BB2XL U1135 ( .B0(n2156), .B1(n2380), .A0N(\register[9][31] ), .A1N(
        n2376), .Y(n395) );
  OAI2BB2XL U1136 ( .B0(n2180), .B1(n2335), .A0N(\register[17][23] ), .A1N(
        n2335), .Y(n643) );
  OAI2BB2XL U1137 ( .B0(n2174), .B1(n2335), .A0N(\register[17][25] ), .A1N(
        n2336), .Y(n645) );
  OAI2BB2XL U1138 ( .B0(n2171), .B1(n2335), .A0N(\register[17][26] ), .A1N(
        n2336), .Y(n646) );
  OAI2BB2XL U1139 ( .B0(n2168), .B1(n2335), .A0N(\register[17][27] ), .A1N(
        n2336), .Y(n647) );
  OAI2BB2XL U1140 ( .B0(n2165), .B1(n2335), .A0N(\register[17][28] ), .A1N(
        n2336), .Y(n648) );
  OAI2BB2XL U1141 ( .B0(n2162), .B1(n2335), .A0N(\register[17][29] ), .A1N(
        n2336), .Y(n649) );
  OAI2BB2XL U1142 ( .B0(n2159), .B1(n2335), .A0N(\register[17][30] ), .A1N(
        n2335), .Y(n650) );
  OAI2BB2XL U1143 ( .B0(n2156), .B1(n2335), .A0N(\register[17][31] ), .A1N(
        n2336), .Y(n651) );
  OAI2BB2XL U1144 ( .B0(n2179), .B1(n2288), .A0N(\register[25][23] ), .A1N(
        n2288), .Y(n899) );
  OAI2BB2XL U1145 ( .B0(n2173), .B1(n2288), .A0N(\register[25][25] ), .A1N(
        n2289), .Y(n901) );
  OAI2BB2XL U1146 ( .B0(n2170), .B1(n2288), .A0N(\register[25][26] ), .A1N(
        n2289), .Y(n902) );
  OAI2BB2XL U1147 ( .B0(n2167), .B1(n2288), .A0N(\register[25][27] ), .A1N(
        n2289), .Y(n903) );
  OAI2BB2XL U1148 ( .B0(n2164), .B1(n2288), .A0N(\register[25][28] ), .A1N(
        n2289), .Y(n904) );
  OAI2BB2XL U1149 ( .B0(n2161), .B1(n2288), .A0N(\register[25][29] ), .A1N(
        n2289), .Y(n905) );
  OAI2BB2XL U1150 ( .B0(n2158), .B1(n2288), .A0N(\register[25][30] ), .A1N(
        n2285), .Y(n906) );
  OAI2BB2XL U1151 ( .B0(n2155), .B1(n2288), .A0N(\register[25][31] ), .A1N(
        n2285), .Y(n907) );
  OAI2BB2XL U1152 ( .B0(n2180), .B1(n2362), .A0N(\register[12][23] ), .A1N(
        n2362), .Y(n483) );
  OAI2BB2XL U1153 ( .B0(n2180), .B1(n2350), .A0N(\register[14][23] ), .A1N(
        n2350), .Y(n547) );
  OAI2BB2XL U1154 ( .B0(n2179), .B1(n2318), .A0N(\register[20][23] ), .A1N(
        n2318), .Y(n739) );
  OAI2BB2XL U1155 ( .B0(n2179), .B1(n2306), .A0N(\register[22][23] ), .A1N(
        n2306), .Y(n803) );
  OAI2BB2XL U1156 ( .B0(n2179), .B1(n2270), .A0N(\register[28][23] ), .A1N(
        n2270), .Y(n995) );
  OAI2BB2XL U1157 ( .B0(n2179), .B1(n2260), .A0N(\register[30][23] ), .A1N(
        n2260), .Y(n1059) );
  OAI2BB2XL U1158 ( .B0(n2174), .B1(n2362), .A0N(\register[12][25] ), .A1N(
        n2363), .Y(n485) );
  OAI2BB2XL U1159 ( .B0(n2171), .B1(n2362), .A0N(\register[12][26] ), .A1N(
        n2363), .Y(n486) );
  OAI2BB2XL U1160 ( .B0(n2168), .B1(n2362), .A0N(\register[12][27] ), .A1N(
        n2363), .Y(n487) );
  OAI2BB2XL U1161 ( .B0(n2165), .B1(n2362), .A0N(\register[12][28] ), .A1N(
        n2363), .Y(n488) );
  OAI2BB2XL U1162 ( .B0(n2162), .B1(n2362), .A0N(\register[12][29] ), .A1N(
        n2363), .Y(n489) );
  OAI2BB2XL U1163 ( .B0(n2174), .B1(n2350), .A0N(\register[14][25] ), .A1N(
        n2351), .Y(n549) );
  OAI2BB2XL U1164 ( .B0(n2171), .B1(n2350), .A0N(\register[14][26] ), .A1N(
        n2351), .Y(n550) );
  OAI2BB2XL U1165 ( .B0(n2168), .B1(n2350), .A0N(\register[14][27] ), .A1N(
        n2351), .Y(n551) );
  OAI2BB2XL U1166 ( .B0(n2165), .B1(n2350), .A0N(\register[14][28] ), .A1N(
        n2351), .Y(n552) );
  OAI2BB2XL U1167 ( .B0(n2162), .B1(n2350), .A0N(\register[14][29] ), .A1N(
        n2351), .Y(n553) );
  OAI2BB2XL U1168 ( .B0(n2173), .B1(n2318), .A0N(\register[20][25] ), .A1N(
        n2319), .Y(n741) );
  OAI2BB2XL U1169 ( .B0(n2170), .B1(n2318), .A0N(\register[20][26] ), .A1N(
        n2319), .Y(n742) );
  OAI2BB2XL U1170 ( .B0(n2167), .B1(n2318), .A0N(\register[20][27] ), .A1N(
        n2319), .Y(n743) );
  OAI2BB2XL U1171 ( .B0(n2164), .B1(n2318), .A0N(\register[20][28] ), .A1N(
        n2319), .Y(n744) );
  OAI2BB2XL U1172 ( .B0(n2161), .B1(n2318), .A0N(\register[20][29] ), .A1N(
        n2319), .Y(n745) );
  OAI2BB2XL U1173 ( .B0(n2173), .B1(n2306), .A0N(\register[22][25] ), .A1N(
        n2307), .Y(n805) );
  OAI2BB2XL U1174 ( .B0(n2170), .B1(n2306), .A0N(\register[22][26] ), .A1N(
        n2307), .Y(n806) );
  OAI2BB2XL U1175 ( .B0(n2167), .B1(n2306), .A0N(\register[22][27] ), .A1N(
        n2307), .Y(n807) );
  OAI2BB2XL U1176 ( .B0(n2164), .B1(n2306), .A0N(\register[22][28] ), .A1N(
        n2307), .Y(n808) );
  OAI2BB2XL U1177 ( .B0(n2161), .B1(n2306), .A0N(\register[22][29] ), .A1N(
        n2307), .Y(n809) );
  OAI2BB2XL U1178 ( .B0(n2173), .B1(n2270), .A0N(\register[28][25] ), .A1N(
        n2271), .Y(n997) );
  OAI2BB2XL U1179 ( .B0(n2170), .B1(n2270), .A0N(\register[28][26] ), .A1N(
        n2271), .Y(n998) );
  OAI2BB2XL U1180 ( .B0(n2167), .B1(n2270), .A0N(\register[28][27] ), .A1N(
        n2271), .Y(n999) );
  OAI2BB2XL U1181 ( .B0(n2164), .B1(n2270), .A0N(\register[28][28] ), .A1N(
        n2271), .Y(n1000) );
  OAI2BB2XL U1182 ( .B0(n2161), .B1(n2270), .A0N(\register[28][29] ), .A1N(
        n2271), .Y(n1001) );
  OAI2BB2XL U1183 ( .B0(n2173), .B1(n2260), .A0N(\register[30][25] ), .A1N(
        n2261), .Y(n1061) );
  OAI2BB2XL U1184 ( .B0(n2170), .B1(n2260), .A0N(\register[30][26] ), .A1N(
        n2261), .Y(n1062) );
  OAI2BB2XL U1185 ( .B0(n2167), .B1(n2260), .A0N(\register[30][27] ), .A1N(
        n2261), .Y(n1063) );
  OAI2BB2XL U1186 ( .B0(n2164), .B1(n2260), .A0N(\register[30][28] ), .A1N(
        n2261), .Y(n1064) );
  OAI2BB2XL U1187 ( .B0(n2161), .B1(n2260), .A0N(\register[30][29] ), .A1N(
        n2261), .Y(n1065) );
  OAI2BB2XL U1188 ( .B0(n2181), .B1(n2407), .A0N(\register[4][23] ), .A1N(
        n2407), .Y(n227) );
  OAI2BB2XL U1189 ( .B0(n2181), .B1(n2395), .A0N(\register[6][23] ), .A1N(
        n2395), .Y(n291) );
  OAI2BB2XL U1190 ( .B0(n2175), .B1(n2407), .A0N(\register[4][25] ), .A1N(
        n2408), .Y(n229) );
  OAI2BB2XL U1191 ( .B0(n2172), .B1(n2407), .A0N(\register[4][26] ), .A1N(
        n2408), .Y(n230) );
  OAI2BB2XL U1192 ( .B0(n2169), .B1(n2407), .A0N(\register[4][27] ), .A1N(
        n2408), .Y(n231) );
  OAI2BB2XL U1193 ( .B0(n2166), .B1(n2407), .A0N(\register[4][28] ), .A1N(
        n2408), .Y(n232) );
  OAI2BB2XL U1194 ( .B0(n2163), .B1(n2407), .A0N(\register[4][29] ), .A1N(
        n2408), .Y(n233) );
  OAI2BB2XL U1195 ( .B0(n2175), .B1(n2395), .A0N(\register[6][25] ), .A1N(
        n2396), .Y(n293) );
  OAI2BB2XL U1196 ( .B0(n2172), .B1(n2395), .A0N(\register[6][26] ), .A1N(
        n2396), .Y(n294) );
  OAI2BB2XL U1197 ( .B0(n2169), .B1(n2395), .A0N(\register[6][27] ), .A1N(
        n2396), .Y(n295) );
  OAI2BB2XL U1198 ( .B0(n2166), .B1(n2395), .A0N(\register[6][28] ), .A1N(
        n2396), .Y(n296) );
  OAI2BB2XL U1199 ( .B0(n2163), .B1(n2395), .A0N(\register[6][29] ), .A1N(
        n2396), .Y(n297) );
  OAI2BB2XL U1200 ( .B0(n2159), .B1(n2362), .A0N(\register[12][30] ), .A1N(
        n2358), .Y(n490) );
  OAI2BB2XL U1201 ( .B0(n2156), .B1(n2362), .A0N(\register[12][31] ), .A1N(
        n2358), .Y(n491) );
  OAI2BB2XL U1202 ( .B0(n2159), .B1(n2350), .A0N(\register[14][30] ), .A1N(
        n2350), .Y(n554) );
  OAI2BB2XL U1203 ( .B0(n2156), .B1(n2350), .A0N(\register[14][31] ), .A1N(
        n2350), .Y(n555) );
  OAI2BB2XL U1204 ( .B0(n2158), .B1(n2318), .A0N(\register[20][30] ), .A1N(
        n2314), .Y(n746) );
  OAI2BB2XL U1205 ( .B0(n2155), .B1(n2318), .A0N(\register[20][31] ), .A1N(
        n2314), .Y(n747) );
  OAI2BB2XL U1206 ( .B0(n2158), .B1(n2306), .A0N(\register[22][30] ), .A1N(
        n2302), .Y(n810) );
  OAI2BB2XL U1207 ( .B0(n2155), .B1(n2306), .A0N(\register[22][31] ), .A1N(
        n2302), .Y(n811) );
  OAI2BB2XL U1208 ( .B0(n2158), .B1(n2270), .A0N(\register[28][30] ), .A1N(
        n2267), .Y(n1002) );
  OAI2BB2XL U1209 ( .B0(n2155), .B1(n2270), .A0N(\register[28][31] ), .A1N(
        n2267), .Y(n1003) );
  OAI2BB2XL U1210 ( .B0(n2158), .B1(n2260), .A0N(\register[30][30] ), .A1N(
        n2257), .Y(n1066) );
  OAI2BB2XL U1211 ( .B0(n2155), .B1(n2260), .A0N(\register[30][31] ), .A1N(
        n2257), .Y(n1067) );
  OAI2BB2XL U1212 ( .B0(n2160), .B1(n2407), .A0N(\register[4][30] ), .A1N(
        n2403), .Y(n234) );
  OAI2BB2XL U1213 ( .B0(n2157), .B1(n2407), .A0N(\register[4][31] ), .A1N(
        n2403), .Y(n235) );
  OAI2BB2XL U1214 ( .B0(n2160), .B1(n2395), .A0N(\register[6][30] ), .A1N(
        n2394), .Y(n298) );
  OAI2BB2XL U1215 ( .B0(n2157), .B1(n2395), .A0N(\register[6][31] ), .A1N(
        n2393), .Y(n299) );
  OAI2BB2XL U1216 ( .B0(n2180), .B1(n2386), .A0N(\register[8][23] ), .A1N(
        n2386), .Y(n355) );
  OAI2BB2XL U1217 ( .B0(n2174), .B1(n2386), .A0N(\register[8][25] ), .A1N(
        n2387), .Y(n357) );
  OAI2BB2XL U1218 ( .B0(n2171), .B1(n2386), .A0N(\register[8][26] ), .A1N(
        n2387), .Y(n358) );
  OAI2BB2XL U1219 ( .B0(n2168), .B1(n2386), .A0N(\register[8][27] ), .A1N(
        n2387), .Y(n359) );
  OAI2BB2XL U1220 ( .B0(n2165), .B1(n2386), .A0N(\register[8][28] ), .A1N(
        n2387), .Y(n360) );
  OAI2BB2XL U1221 ( .B0(n2162), .B1(n2386), .A0N(\register[8][29] ), .A1N(
        n2387), .Y(n361) );
  OAI2BB2XL U1222 ( .B0(n2159), .B1(n2386), .A0N(\register[8][30] ), .A1N(
        n2382), .Y(n362) );
  OAI2BB2XL U1223 ( .B0(n2156), .B1(n2386), .A0N(\register[8][31] ), .A1N(
        n2382), .Y(n363) );
  OAI2BB2XL U1224 ( .B0(n2180), .B1(n2340), .A0N(\register[16][23] ), .A1N(
        n2340), .Y(n611) );
  OAI2BB2XL U1225 ( .B0(n2174), .B1(n2340), .A0N(\register[16][25] ), .A1N(
        n2341), .Y(n613) );
  OAI2BB2XL U1226 ( .B0(n2171), .B1(n2340), .A0N(\register[16][26] ), .A1N(
        n2341), .Y(n614) );
  OAI2BB2XL U1227 ( .B0(n2168), .B1(n2340), .A0N(\register[16][27] ), .A1N(
        n2341), .Y(n615) );
  OAI2BB2XL U1228 ( .B0(n2165), .B1(n2340), .A0N(\register[16][28] ), .A1N(
        n2341), .Y(n616) );
  OAI2BB2XL U1229 ( .B0(n2162), .B1(n2340), .A0N(\register[16][29] ), .A1N(
        n2341), .Y(n617) );
  OAI2BB2XL U1230 ( .B0(n2159), .B1(n2340), .A0N(\register[16][30] ), .A1N(
        n2338), .Y(n618) );
  OAI2BB2XL U1231 ( .B0(n2156), .B1(n2340), .A0N(\register[16][31] ), .A1N(
        n2338), .Y(n619) );
  OAI2BB2XL U1232 ( .B0(n2179), .B1(n2294), .A0N(\register[24][23] ), .A1N(
        n2294), .Y(n867) );
  OAI2BB2XL U1233 ( .B0(n2173), .B1(n2294), .A0N(\register[24][25] ), .A1N(
        n2295), .Y(n869) );
  OAI2BB2XL U1234 ( .B0(n2170), .B1(n2294), .A0N(\register[24][26] ), .A1N(
        n2295), .Y(n870) );
  OAI2BB2XL U1235 ( .B0(n2167), .B1(n2294), .A0N(\register[24][27] ), .A1N(
        n2295), .Y(n871) );
  OAI2BB2XL U1236 ( .B0(n2164), .B1(n2294), .A0N(\register[24][28] ), .A1N(
        n2295), .Y(n872) );
  OAI2BB2XL U1237 ( .B0(n2161), .B1(n2294), .A0N(\register[24][29] ), .A1N(
        n2295), .Y(n873) );
  OAI2BB2XL U1238 ( .B0(n2158), .B1(n2294), .A0N(\register[24][30] ), .A1N(
        n2290), .Y(n874) );
  OAI2BB2XL U1239 ( .B0(n2155), .B1(n2294), .A0N(\register[24][31] ), .A1N(
        n2290), .Y(n875) );
  OAI2BB2XL U1240 ( .B0(n2180), .B1(n2356), .A0N(\register[13][23] ), .A1N(
        n2356), .Y(n515) );
  OAI2BB2XL U1241 ( .B0(n2180), .B1(n2342), .A0N(\register[15][23] ), .A1N(
        n2346), .Y(n579) );
  OAI2BB2XL U1242 ( .B0(n2179), .B1(n2312), .A0N(\register[21][23] ), .A1N(
        n2312), .Y(n771) );
  OAI2BB2XL U1243 ( .B0(n2179), .B1(n2300), .A0N(\register[23][23] ), .A1N(
        n2300), .Y(n835) );
  OAI2BB2XL U1244 ( .B0(n2179), .B1(n2264), .A0N(\register[29][23] ), .A1N(
        n2264), .Y(n1027) );
  OAI2BB2XL U1245 ( .B0(n2179), .B1(n2254), .A0N(\register[31][23] ), .A1N(
        n2254), .Y(n1091) );
  OAI2BB2XL U1246 ( .B0(n2174), .B1(n2356), .A0N(\register[13][25] ), .A1N(
        n2357), .Y(n517) );
  OAI2BB2XL U1247 ( .B0(n2171), .B1(n2356), .A0N(\register[13][26] ), .A1N(
        n2357), .Y(n518) );
  OAI2BB2XL U1248 ( .B0(n2168), .B1(n2356), .A0N(\register[13][27] ), .A1N(
        n2357), .Y(n519) );
  OAI2BB2XL U1249 ( .B0(n2165), .B1(n2356), .A0N(\register[13][28] ), .A1N(
        n2357), .Y(n520) );
  OAI2BB2XL U1250 ( .B0(n2162), .B1(n2356), .A0N(\register[13][29] ), .A1N(
        n2357), .Y(n521) );
  OAI2BB2XL U1251 ( .B0(n2174), .B1(n2342), .A0N(\register[15][25] ), .A1N(
        n2346), .Y(n581) );
  OAI2BB2XL U1252 ( .B0(n2171), .B1(n2342), .A0N(\register[15][26] ), .A1N(
        n2346), .Y(n582) );
  OAI2BB2XL U1253 ( .B0(n2168), .B1(n2342), .A0N(\register[15][27] ), .A1N(
        n2346), .Y(n583) );
  OAI2BB2XL U1254 ( .B0(n2165), .B1(n2342), .A0N(\register[15][28] ), .A1N(
        n2346), .Y(n584) );
  OAI2BB2XL U1255 ( .B0(n2162), .B1(n2343), .A0N(\register[15][29] ), .A1N(
        n2346), .Y(n585) );
  OAI2BB2XL U1256 ( .B0(n2173), .B1(n2312), .A0N(\register[21][25] ), .A1N(
        n2313), .Y(n773) );
  OAI2BB2XL U1257 ( .B0(n2170), .B1(n2312), .A0N(\register[21][26] ), .A1N(
        n2313), .Y(n774) );
  OAI2BB2XL U1258 ( .B0(n2167), .B1(n2312), .A0N(\register[21][27] ), .A1N(
        n2313), .Y(n775) );
  OAI2BB2XL U1259 ( .B0(n2164), .B1(n2312), .A0N(\register[21][28] ), .A1N(
        n2313), .Y(n776) );
  OAI2BB2XL U1260 ( .B0(n2161), .B1(n2312), .A0N(\register[21][29] ), .A1N(
        n2313), .Y(n777) );
  OAI2BB2XL U1261 ( .B0(n2173), .B1(n2300), .A0N(\register[23][25] ), .A1N(
        n2301), .Y(n837) );
  OAI2BB2XL U1262 ( .B0(n2170), .B1(n2300), .A0N(\register[23][26] ), .A1N(
        n2301), .Y(n838) );
  OAI2BB2XL U1263 ( .B0(n2167), .B1(n2300), .A0N(\register[23][27] ), .A1N(
        n2301), .Y(n839) );
  OAI2BB2XL U1264 ( .B0(n2164), .B1(n2300), .A0N(\register[23][28] ), .A1N(
        n2301), .Y(n840) );
  OAI2BB2XL U1265 ( .B0(n2161), .B1(n2300), .A0N(\register[23][29] ), .A1N(
        n2301), .Y(n841) );
  OAI2BB2XL U1266 ( .B0(n2173), .B1(n2264), .A0N(\register[29][25] ), .A1N(
        n2265), .Y(n1029) );
  OAI2BB2XL U1267 ( .B0(n2170), .B1(n2264), .A0N(\register[29][26] ), .A1N(
        n2265), .Y(n1030) );
  OAI2BB2XL U1268 ( .B0(n2167), .B1(n2264), .A0N(\register[29][27] ), .A1N(
        n2265), .Y(n1031) );
  OAI2BB2XL U1269 ( .B0(n2164), .B1(n2264), .A0N(\register[29][28] ), .A1N(
        n2265), .Y(n1032) );
  OAI2BB2XL U1270 ( .B0(n2161), .B1(n2264), .A0N(\register[29][29] ), .A1N(
        n2265), .Y(n1033) );
  OAI2BB2XL U1271 ( .B0(n2173), .B1(n2254), .A0N(\register[31][25] ), .A1N(
        n2255), .Y(n1093) );
  OAI2BB2XL U1272 ( .B0(n2170), .B1(n2254), .A0N(\register[31][26] ), .A1N(
        n2255), .Y(n1094) );
  OAI2BB2XL U1273 ( .B0(n2167), .B1(n2254), .A0N(\register[31][27] ), .A1N(
        n2255), .Y(n1095) );
  OAI2BB2XL U1274 ( .B0(n2164), .B1(n2254), .A0N(\register[31][28] ), .A1N(
        n2255), .Y(n1096) );
  OAI2BB2XL U1275 ( .B0(n2161), .B1(n2254), .A0N(\register[31][29] ), .A1N(
        n2255), .Y(n1097) );
  OAI2BB2XL U1276 ( .B0(n2181), .B1(n2401), .A0N(\register[5][23] ), .A1N(
        n2401), .Y(n259) );
  OAI2BB2XL U1277 ( .B0(n2181), .B1(n2388), .A0N(\register[7][23] ), .A1N(
        n2391), .Y(n323) );
  OAI2BB2XL U1278 ( .B0(n2175), .B1(n2401), .A0N(\register[5][25] ), .A1N(
        n2402), .Y(n261) );
  OAI2BB2XL U1279 ( .B0(n2172), .B1(n2401), .A0N(\register[5][26] ), .A1N(
        n2402), .Y(n262) );
  OAI2BB2XL U1280 ( .B0(n2169), .B1(n2401), .A0N(\register[5][27] ), .A1N(
        n2402), .Y(n263) );
  OAI2BB2XL U1281 ( .B0(n2166), .B1(n2401), .A0N(\register[5][28] ), .A1N(
        n2402), .Y(n264) );
  OAI2BB2XL U1282 ( .B0(n2163), .B1(n2401), .A0N(\register[5][29] ), .A1N(
        n2402), .Y(n265) );
  OAI2BB2XL U1283 ( .B0(n2175), .B1(n2388), .A0N(\register[7][25] ), .A1N(
        n2392), .Y(n325) );
  OAI2BB2XL U1284 ( .B0(n2172), .B1(n2388), .A0N(\register[7][26] ), .A1N(
        n2392), .Y(n326) );
  OAI2BB2XL U1285 ( .B0(n2169), .B1(n2388), .A0N(\register[7][27] ), .A1N(
        n2392), .Y(n327) );
  OAI2BB2XL U1286 ( .B0(n2166), .B1(n2388), .A0N(\register[7][28] ), .A1N(
        n2392), .Y(n328) );
  OAI2BB2XL U1287 ( .B0(n2163), .B1(n2388), .A0N(\register[7][29] ), .A1N(
        n2392), .Y(n329) );
  OAI2BB2XL U1288 ( .B0(n2159), .B1(n2356), .A0N(\register[13][30] ), .A1N(
        n2352), .Y(n522) );
  OAI2BB2XL U1289 ( .B0(n2156), .B1(n2356), .A0N(\register[13][31] ), .A1N(
        n2352), .Y(n523) );
  OAI2BB2XL U1290 ( .B0(n2159), .B1(n2343), .A0N(\register[15][30] ), .A1N(
        n2342), .Y(n586) );
  OAI2BB2XL U1291 ( .B0(n2156), .B1(n2343), .A0N(\register[15][31] ), .A1N(
        n2342), .Y(n587) );
  OAI2BB2XL U1292 ( .B0(n2158), .B1(n2312), .A0N(\register[21][30] ), .A1N(
        n2308), .Y(n778) );
  OAI2BB2XL U1293 ( .B0(n2155), .B1(n2312), .A0N(\register[21][31] ), .A1N(
        n2308), .Y(n779) );
  OAI2BB2XL U1294 ( .B0(n2158), .B1(n2300), .A0N(\register[23][30] ), .A1N(
        n2296), .Y(n842) );
  OAI2BB2XL U1295 ( .B0(n2155), .B1(n2300), .A0N(\register[23][31] ), .A1N(
        n2296), .Y(n843) );
  OAI2BB2XL U1296 ( .B0(n2158), .B1(n2264), .A0N(\register[29][30] ), .A1N(
        n2262), .Y(n1034) );
  OAI2BB2XL U1297 ( .B0(n2155), .B1(n2264), .A0N(\register[29][31] ), .A1N(
        n2262), .Y(n1035) );
  OAI2BB2XL U1298 ( .B0(n2158), .B1(n2254), .A0N(\register[31][30] ), .A1N(
        n2250), .Y(n1098) );
  OAI2BB2XL U1299 ( .B0(n2155), .B1(n2254), .A0N(\register[31][31] ), .A1N(
        n2250), .Y(n1099) );
  OAI2BB2XL U1300 ( .B0(n2160), .B1(n2401), .A0N(\register[5][30] ), .A1N(
        n2397), .Y(n266) );
  OAI2BB2XL U1301 ( .B0(n2157), .B1(n2401), .A0N(\register[5][31] ), .A1N(
        n2397), .Y(n267) );
  OAI2BB2XL U1302 ( .B0(n2160), .B1(n2388), .A0N(\register[7][30] ), .A1N(
        n2388), .Y(n330) );
  OAI2BB2XL U1303 ( .B0(n2157), .B1(n2390), .A0N(\register[7][31] ), .A1N(
        n2388), .Y(n331) );
  OAI2BB2XL U1304 ( .B0(n2248), .B1(n2373), .A0N(\register[10][0] ), .A1N(
        n2370), .Y(n396) );
  OAI2BB2XL U1305 ( .B0(n2245), .B1(n2372), .A0N(\register[10][1] ), .A1N(
        n2370), .Y(n397) );
  OAI2BB2XL U1306 ( .B0(n2242), .B1(n2372), .A0N(\register[10][2] ), .A1N(
        n2370), .Y(n398) );
  OAI2BB2XL U1307 ( .B0(n2240), .B1(n2372), .A0N(\register[10][3] ), .A1N(
        n2375), .Y(n399) );
  OAI2BB2XL U1308 ( .B0(n2237), .B1(n2372), .A0N(\register[10][4] ), .A1N(
        n2370), .Y(n400) );
  OAI2BB2XL U1309 ( .B0(n2234), .B1(n2372), .A0N(\register[10][5] ), .A1N(
        n2375), .Y(n401) );
  OAI2BB2XL U1310 ( .B0(n2231), .B1(n2372), .A0N(\register[10][6] ), .A1N(
        n2375), .Y(n402) );
  OAI2BB2XL U1311 ( .B0(n2228), .B1(n2372), .A0N(\register[10][7] ), .A1N(
        n2375), .Y(n403) );
  OAI2BB2XL U1312 ( .B0(n2225), .B1(n2372), .A0N(\register[10][8] ), .A1N(
        n2375), .Y(n404) );
  OAI2BB2XL U1313 ( .B0(n2222), .B1(n2372), .A0N(\register[10][9] ), .A1N(
        n2375), .Y(n405) );
  OAI2BB2XL U1314 ( .B0(n2219), .B1(n2372), .A0N(\register[10][10] ), .A1N(
        n2375), .Y(n406) );
  OAI2BB2XL U1315 ( .B0(n2216), .B1(n2372), .A0N(\register[10][11] ), .A1N(
        n2375), .Y(n407) );
  OAI2BB2XL U1316 ( .B0(n2213), .B1(n2372), .A0N(\register[10][12] ), .A1N(
        n2375), .Y(n408) );
  OAI2BB2XL U1317 ( .B0(n2210), .B1(n2373), .A0N(\register[10][13] ), .A1N(
        n2375), .Y(n409) );
  OAI2BB2XL U1318 ( .B0(n2207), .B1(n2373), .A0N(\register[10][14] ), .A1N(
        n2375), .Y(n410) );
  OAI2BB2XL U1319 ( .B0(n2204), .B1(n2373), .A0N(\register[10][15] ), .A1N(
        n2374), .Y(n411) );
  OAI2BB2XL U1320 ( .B0(n2201), .B1(n2373), .A0N(\register[10][16] ), .A1N(
        n2375), .Y(n412) );
  OAI2BB2XL U1321 ( .B0(n2198), .B1(n2373), .A0N(\register[10][17] ), .A1N(
        n2374), .Y(n413) );
  OAI2BB2XL U1322 ( .B0(n2195), .B1(n2373), .A0N(\register[10][18] ), .A1N(
        n2374), .Y(n414) );
  OAI2BB2XL U1323 ( .B0(n2192), .B1(n2373), .A0N(\register[10][19] ), .A1N(
        n2374), .Y(n415) );
  OAI2BB2XL U1324 ( .B0(n2189), .B1(n2373), .A0N(\register[10][20] ), .A1N(
        n2374), .Y(n416) );
  OAI2BB2XL U1325 ( .B0(n2186), .B1(n2373), .A0N(\register[10][21] ), .A1N(
        n2374), .Y(n417) );
  OAI2BB2XL U1326 ( .B0(n2183), .B1(n2373), .A0N(\register[10][22] ), .A1N(
        n2375), .Y(n418) );
  OAI2BB2XL U1327 ( .B0(n2177), .B1(n2373), .A0N(\register[10][24] ), .A1N(
        n2375), .Y(n420) );
  OAI2BB2XL U1328 ( .B0(n2248), .B1(n2367), .A0N(\register[11][0] ), .A1N(
        n2364), .Y(n428) );
  OAI2BB2XL U1329 ( .B0(n2245), .B1(n2366), .A0N(\register[11][1] ), .A1N(
        n2364), .Y(n429) );
  OAI2BB2XL U1330 ( .B0(n2242), .B1(n2366), .A0N(\register[11][2] ), .A1N(
        n2364), .Y(n430) );
  OAI2BB2XL U1331 ( .B0(n2240), .B1(n2366), .A0N(\register[11][3] ), .A1N(
        n2369), .Y(n431) );
  OAI2BB2XL U1332 ( .B0(n2237), .B1(n2366), .A0N(\register[11][4] ), .A1N(
        n2364), .Y(n432) );
  OAI2BB2XL U1333 ( .B0(n2234), .B1(n2366), .A0N(\register[11][5] ), .A1N(
        n2369), .Y(n433) );
  OAI2BB2XL U1334 ( .B0(n2231), .B1(n2366), .A0N(\register[11][6] ), .A1N(
        n2369), .Y(n434) );
  OAI2BB2XL U1335 ( .B0(n2228), .B1(n2366), .A0N(\register[11][7] ), .A1N(
        n2369), .Y(n435) );
  OAI2BB2XL U1336 ( .B0(n2225), .B1(n2366), .A0N(\register[11][8] ), .A1N(
        n2369), .Y(n436) );
  OAI2BB2XL U1337 ( .B0(n2222), .B1(n2366), .A0N(\register[11][9] ), .A1N(
        n2369), .Y(n437) );
  OAI2BB2XL U1338 ( .B0(n2219), .B1(n2366), .A0N(\register[11][10] ), .A1N(
        n2369), .Y(n438) );
  OAI2BB2XL U1339 ( .B0(n2216), .B1(n2366), .A0N(\register[11][11] ), .A1N(
        n2369), .Y(n439) );
  OAI2BB2XL U1340 ( .B0(n2213), .B1(n2366), .A0N(\register[11][12] ), .A1N(
        n2369), .Y(n440) );
  OAI2BB2XL U1341 ( .B0(n2210), .B1(n2367), .A0N(\register[11][13] ), .A1N(
        n2369), .Y(n441) );
  OAI2BB2XL U1342 ( .B0(n2207), .B1(n2367), .A0N(\register[11][14] ), .A1N(
        n2369), .Y(n442) );
  OAI2BB2XL U1343 ( .B0(n2204), .B1(n2367), .A0N(\register[11][15] ), .A1N(
        n2368), .Y(n443) );
  OAI2BB2XL U1344 ( .B0(n2201), .B1(n2367), .A0N(\register[11][16] ), .A1N(
        n2369), .Y(n444) );
  OAI2BB2XL U1345 ( .B0(n2198), .B1(n2367), .A0N(\register[11][17] ), .A1N(
        n2368), .Y(n445) );
  OAI2BB2XL U1346 ( .B0(n2195), .B1(n2367), .A0N(\register[11][18] ), .A1N(
        n2368), .Y(n446) );
  OAI2BB2XL U1347 ( .B0(n2192), .B1(n2367), .A0N(\register[11][19] ), .A1N(
        n2368), .Y(n447) );
  OAI2BB2XL U1348 ( .B0(n2189), .B1(n2367), .A0N(\register[11][20] ), .A1N(
        n2368), .Y(n448) );
  OAI2BB2XL U1349 ( .B0(n2186), .B1(n2367), .A0N(\register[11][21] ), .A1N(
        n2368), .Y(n449) );
  OAI2BB2XL U1350 ( .B0(n2183), .B1(n2367), .A0N(\register[11][22] ), .A1N(
        n2369), .Y(n450) );
  OAI2BB2XL U1351 ( .B0(n2177), .B1(n2367), .A0N(\register[11][24] ), .A1N(
        n2369), .Y(n452) );
  OAI2BB2XL U1352 ( .B0(n2248), .B1(n2329), .A0N(\register[18][0] ), .A1N(
        n2326), .Y(n652) );
  OAI2BB2XL U1353 ( .B0(n2245), .B1(n2328), .A0N(\register[18][1] ), .A1N(
        n2326), .Y(n653) );
  OAI2BB2XL U1354 ( .B0(n2242), .B1(n2328), .A0N(\register[18][2] ), .A1N(
        n2326), .Y(n654) );
  OAI2BB2XL U1355 ( .B0(n2240), .B1(n2328), .A0N(\register[18][3] ), .A1N(
        n2331), .Y(n655) );
  OAI2BB2XL U1356 ( .B0(n2237), .B1(n2328), .A0N(\register[18][4] ), .A1N(
        n2326), .Y(n656) );
  OAI2BB2XL U1357 ( .B0(n2234), .B1(n2328), .A0N(\register[18][5] ), .A1N(
        n2331), .Y(n657) );
  OAI2BB2XL U1358 ( .B0(n2231), .B1(n2328), .A0N(\register[18][6] ), .A1N(
        n2331), .Y(n658) );
  OAI2BB2XL U1359 ( .B0(n2228), .B1(n2328), .A0N(\register[18][7] ), .A1N(
        n2331), .Y(n659) );
  OAI2BB2XL U1360 ( .B0(n2225), .B1(n2328), .A0N(\register[18][8] ), .A1N(
        n2331), .Y(n660) );
  OAI2BB2XL U1361 ( .B0(n2222), .B1(n2328), .A0N(\register[18][9] ), .A1N(
        n2331), .Y(n661) );
  OAI2BB2XL U1362 ( .B0(n2219), .B1(n2328), .A0N(\register[18][10] ), .A1N(
        n2331), .Y(n662) );
  OAI2BB2XL U1363 ( .B0(n2216), .B1(n2328), .A0N(\register[18][11] ), .A1N(
        n2331), .Y(n663) );
  OAI2BB2XL U1364 ( .B0(n2213), .B1(n2328), .A0N(\register[18][12] ), .A1N(
        n2331), .Y(n664) );
  OAI2BB2XL U1365 ( .B0(n2210), .B1(n2329), .A0N(\register[18][13] ), .A1N(
        n2331), .Y(n665) );
  OAI2BB2XL U1366 ( .B0(n2207), .B1(n2329), .A0N(\register[18][14] ), .A1N(
        n2331), .Y(n666) );
  OAI2BB2XL U1367 ( .B0(n2204), .B1(n2329), .A0N(\register[18][15] ), .A1N(
        n2330), .Y(n667) );
  OAI2BB2XL U1368 ( .B0(n2201), .B1(n2329), .A0N(\register[18][16] ), .A1N(
        n2331), .Y(n668) );
  OAI2BB2XL U1369 ( .B0(n2198), .B1(n2329), .A0N(\register[18][17] ), .A1N(
        n2330), .Y(n669) );
  OAI2BB2XL U1370 ( .B0(n2195), .B1(n2329), .A0N(\register[18][18] ), .A1N(
        n2330), .Y(n670) );
  OAI2BB2XL U1371 ( .B0(n2192), .B1(n2329), .A0N(\register[18][19] ), .A1N(
        n2330), .Y(n671) );
  OAI2BB2XL U1372 ( .B0(n2189), .B1(n2329), .A0N(\register[18][20] ), .A1N(
        n2330), .Y(n672) );
  OAI2BB2XL U1373 ( .B0(n2186), .B1(n2329), .A0N(\register[18][21] ), .A1N(
        n2330), .Y(n673) );
  OAI2BB2XL U1374 ( .B0(n2183), .B1(n2329), .A0N(\register[18][22] ), .A1N(
        n2331), .Y(n674) );
  OAI2BB2XL U1375 ( .B0(n2177), .B1(n2329), .A0N(\register[18][24] ), .A1N(
        n2331), .Y(n676) );
  OAI2BB2XL U1376 ( .B0(n2248), .B1(n2323), .A0N(\register[19][0] ), .A1N(
        n2320), .Y(n684) );
  OAI2BB2XL U1377 ( .B0(n2245), .B1(n2322), .A0N(\register[19][1] ), .A1N(
        n2320), .Y(n685) );
  OAI2BB2XL U1378 ( .B0(n2242), .B1(n2322), .A0N(\register[19][2] ), .A1N(
        n2320), .Y(n686) );
  OAI2BB2XL U1379 ( .B0(n2240), .B1(n2322), .A0N(\register[19][3] ), .A1N(
        n2325), .Y(n687) );
  OAI2BB2XL U1380 ( .B0(n2237), .B1(n2322), .A0N(\register[19][4] ), .A1N(
        n2320), .Y(n688) );
  OAI2BB2XL U1381 ( .B0(n2234), .B1(n2322), .A0N(\register[19][5] ), .A1N(
        n2325), .Y(n689) );
  OAI2BB2XL U1382 ( .B0(n2231), .B1(n2322), .A0N(\register[19][6] ), .A1N(
        n2325), .Y(n690) );
  OAI2BB2XL U1383 ( .B0(n2228), .B1(n2322), .A0N(\register[19][7] ), .A1N(
        n2325), .Y(n691) );
  OAI2BB2XL U1384 ( .B0(n2225), .B1(n2322), .A0N(\register[19][8] ), .A1N(
        n2325), .Y(n692) );
  OAI2BB2XL U1385 ( .B0(n2222), .B1(n2322), .A0N(\register[19][9] ), .A1N(
        n2325), .Y(n693) );
  OAI2BB2XL U1386 ( .B0(n2219), .B1(n2322), .A0N(\register[19][10] ), .A1N(
        n2325), .Y(n694) );
  OAI2BB2XL U1387 ( .B0(n2216), .B1(n2322), .A0N(\register[19][11] ), .A1N(
        n2325), .Y(n695) );
  OAI2BB2XL U1388 ( .B0(n2213), .B1(n2322), .A0N(\register[19][12] ), .A1N(
        n2325), .Y(n696) );
  OAI2BB2XL U1389 ( .B0(n2210), .B1(n2323), .A0N(\register[19][13] ), .A1N(
        n2325), .Y(n697) );
  OAI2BB2XL U1390 ( .B0(n2207), .B1(n2323), .A0N(\register[19][14] ), .A1N(
        n2325), .Y(n698) );
  OAI2BB2XL U1391 ( .B0(n2204), .B1(n2323), .A0N(\register[19][15] ), .A1N(
        n2324), .Y(n699) );
  OAI2BB2XL U1392 ( .B0(n2201), .B1(n2323), .A0N(\register[19][16] ), .A1N(
        n2325), .Y(n700) );
  OAI2BB2XL U1393 ( .B0(n2198), .B1(n2323), .A0N(\register[19][17] ), .A1N(
        n2324), .Y(n701) );
  OAI2BB2XL U1394 ( .B0(n2195), .B1(n2323), .A0N(\register[19][18] ), .A1N(
        n2324), .Y(n702) );
  OAI2BB2XL U1395 ( .B0(n2192), .B1(n2323), .A0N(\register[19][19] ), .A1N(
        n2324), .Y(n703) );
  OAI2BB2XL U1396 ( .B0(n2189), .B1(n2323), .A0N(\register[19][20] ), .A1N(
        n2324), .Y(n704) );
  OAI2BB2XL U1397 ( .B0(n2186), .B1(n2323), .A0N(\register[19][21] ), .A1N(
        n2324), .Y(n705) );
  OAI2BB2XL U1398 ( .B0(n2183), .B1(n2323), .A0N(\register[19][22] ), .A1N(
        n2325), .Y(n706) );
  OAI2BB2XL U1399 ( .B0(n2177), .B1(n2323), .A0N(\register[19][24] ), .A1N(
        n2325), .Y(n708) );
  OAI2BB2XL U1400 ( .B0(n2247), .B1(n2281), .A0N(\register[26][0] ), .A1N(
        n2278), .Y(n908) );
  OAI2BB2XL U1401 ( .B0(n2244), .B1(n2280), .A0N(\register[26][1] ), .A1N(
        n2278), .Y(n909) );
  OAI2BB2XL U1402 ( .B0(n2241), .B1(n2280), .A0N(\register[26][2] ), .A1N(
        n2278), .Y(n910) );
  OAI2BB2XL U1403 ( .B0(n2239), .B1(n2280), .A0N(\register[26][3] ), .A1N(
        n2283), .Y(n911) );
  OAI2BB2XL U1404 ( .B0(n2236), .B1(n2280), .A0N(\register[26][4] ), .A1N(
        n2278), .Y(n912) );
  OAI2BB2XL U1405 ( .B0(n2233), .B1(n2280), .A0N(\register[26][5] ), .A1N(
        n2283), .Y(n913) );
  OAI2BB2XL U1406 ( .B0(n2230), .B1(n2280), .A0N(\register[26][6] ), .A1N(
        n2283), .Y(n914) );
  OAI2BB2XL U1407 ( .B0(n2227), .B1(n2280), .A0N(\register[26][7] ), .A1N(
        n2283), .Y(n915) );
  OAI2BB2XL U1408 ( .B0(n2224), .B1(n2280), .A0N(\register[26][8] ), .A1N(
        n2283), .Y(n916) );
  OAI2BB2XL U1409 ( .B0(n2221), .B1(n2280), .A0N(\register[26][9] ), .A1N(
        n2283), .Y(n917) );
  OAI2BB2XL U1410 ( .B0(n2218), .B1(n2280), .A0N(\register[26][10] ), .A1N(
        n2283), .Y(n918) );
  OAI2BB2XL U1411 ( .B0(n2215), .B1(n2280), .A0N(\register[26][11] ), .A1N(
        n2283), .Y(n919) );
  OAI2BB2XL U1412 ( .B0(n2212), .B1(n2280), .A0N(\register[26][12] ), .A1N(
        n2283), .Y(n920) );
  OAI2BB2XL U1413 ( .B0(n2209), .B1(n2281), .A0N(\register[26][13] ), .A1N(
        n2283), .Y(n921) );
  OAI2BB2XL U1414 ( .B0(n2206), .B1(n2281), .A0N(\register[26][14] ), .A1N(
        n2283), .Y(n922) );
  OAI2BB2XL U1415 ( .B0(n2203), .B1(n2281), .A0N(\register[26][15] ), .A1N(
        n2282), .Y(n923) );
  OAI2BB2XL U1416 ( .B0(n2200), .B1(n2281), .A0N(\register[26][16] ), .A1N(
        n2283), .Y(n924) );
  OAI2BB2XL U1417 ( .B0(n2197), .B1(n2281), .A0N(\register[26][17] ), .A1N(
        n2282), .Y(n925) );
  OAI2BB2XL U1418 ( .B0(n2194), .B1(n2281), .A0N(\register[26][18] ), .A1N(
        n2282), .Y(n926) );
  OAI2BB2XL U1419 ( .B0(n2191), .B1(n2281), .A0N(\register[26][19] ), .A1N(
        n2282), .Y(n927) );
  OAI2BB2XL U1420 ( .B0(n2188), .B1(n2281), .A0N(\register[26][20] ), .A1N(
        n2282), .Y(n928) );
  OAI2BB2XL U1421 ( .B0(n2185), .B1(n2281), .A0N(\register[26][21] ), .A1N(
        n2282), .Y(n929) );
  OAI2BB2XL U1422 ( .B0(n2182), .B1(n2281), .A0N(\register[26][22] ), .A1N(
        n2283), .Y(n930) );
  OAI2BB2XL U1423 ( .B0(n2176), .B1(n2281), .A0N(\register[26][24] ), .A1N(
        n2283), .Y(n932) );
  OAI2BB2XL U1424 ( .B0(n2247), .B1(n2275), .A0N(\register[27][0] ), .A1N(
        n2272), .Y(n940) );
  OAI2BB2XL U1425 ( .B0(n2244), .B1(n2274), .A0N(\register[27][1] ), .A1N(
        n2272), .Y(n941) );
  OAI2BB2XL U1426 ( .B0(n2241), .B1(n2274), .A0N(\register[27][2] ), .A1N(
        n2272), .Y(n942) );
  OAI2BB2XL U1427 ( .B0(n2239), .B1(n2274), .A0N(\register[27][3] ), .A1N(
        n2277), .Y(n943) );
  OAI2BB2XL U1428 ( .B0(n2236), .B1(n2274), .A0N(\register[27][4] ), .A1N(
        n2272), .Y(n944) );
  OAI2BB2XL U1429 ( .B0(n2233), .B1(n2274), .A0N(\register[27][5] ), .A1N(
        n2277), .Y(n945) );
  OAI2BB2XL U1430 ( .B0(n2230), .B1(n2274), .A0N(\register[27][6] ), .A1N(
        n2277), .Y(n946) );
  OAI2BB2XL U1431 ( .B0(n2227), .B1(n2274), .A0N(\register[27][7] ), .A1N(
        n2277), .Y(n947) );
  OAI2BB2XL U1432 ( .B0(n2224), .B1(n2274), .A0N(\register[27][8] ), .A1N(
        n2277), .Y(n948) );
  OAI2BB2XL U1433 ( .B0(n2221), .B1(n2274), .A0N(\register[27][9] ), .A1N(
        n2277), .Y(n949) );
  OAI2BB2XL U1434 ( .B0(n2218), .B1(n2274), .A0N(\register[27][10] ), .A1N(
        n2277), .Y(n950) );
  OAI2BB2XL U1435 ( .B0(n2215), .B1(n2274), .A0N(\register[27][11] ), .A1N(
        n2277), .Y(n951) );
  OAI2BB2XL U1436 ( .B0(n2212), .B1(n2274), .A0N(\register[27][12] ), .A1N(
        n2277), .Y(n952) );
  OAI2BB2XL U1437 ( .B0(n2209), .B1(n2275), .A0N(\register[27][13] ), .A1N(
        n2277), .Y(n953) );
  OAI2BB2XL U1438 ( .B0(n2206), .B1(n2275), .A0N(\register[27][14] ), .A1N(
        n2277), .Y(n954) );
  OAI2BB2XL U1439 ( .B0(n2203), .B1(n2275), .A0N(\register[27][15] ), .A1N(
        n2276), .Y(n955) );
  OAI2BB2XL U1440 ( .B0(n2200), .B1(n2275), .A0N(\register[27][16] ), .A1N(
        n2277), .Y(n956) );
  OAI2BB2XL U1441 ( .B0(n2197), .B1(n2275), .A0N(\register[27][17] ), .A1N(
        n2276), .Y(n957) );
  OAI2BB2XL U1442 ( .B0(n2194), .B1(n2275), .A0N(\register[27][18] ), .A1N(
        n2276), .Y(n958) );
  OAI2BB2XL U1443 ( .B0(n2191), .B1(n2275), .A0N(\register[27][19] ), .A1N(
        n2276), .Y(n959) );
  OAI2BB2XL U1444 ( .B0(n2188), .B1(n2275), .A0N(\register[27][20] ), .A1N(
        n2276), .Y(n960) );
  OAI2BB2XL U1445 ( .B0(n2185), .B1(n2275), .A0N(\register[27][21] ), .A1N(
        n2276), .Y(n961) );
  OAI2BB2XL U1446 ( .B0(n2182), .B1(n2275), .A0N(\register[27][22] ), .A1N(
        n2277), .Y(n962) );
  OAI2BB2XL U1447 ( .B0(n2176), .B1(n2275), .A0N(\register[27][24] ), .A1N(
        n2277), .Y(n964) );
  OAI2BB2XL U1448 ( .B0(n2248), .B1(n2379), .A0N(\register[9][0] ), .A1N(n2376), .Y(n364) );
  OAI2BB2XL U1449 ( .B0(n2245), .B1(n2378), .A0N(\register[9][1] ), .A1N(n2376), .Y(n365) );
  OAI2BB2XL U1450 ( .B0(n2242), .B1(n2378), .A0N(\register[9][2] ), .A1N(n2376), .Y(n366) );
  OAI2BB2XL U1451 ( .B0(n2240), .B1(n2378), .A0N(\register[9][3] ), .A1N(n2381), .Y(n367) );
  OAI2BB2XL U1452 ( .B0(n2237), .B1(n2378), .A0N(\register[9][4] ), .A1N(n2376), .Y(n368) );
  OAI2BB2XL U1453 ( .B0(n2234), .B1(n2378), .A0N(\register[9][5] ), .A1N(n2381), .Y(n369) );
  OAI2BB2XL U1454 ( .B0(n2231), .B1(n2378), .A0N(\register[9][6] ), .A1N(n2381), .Y(n370) );
  OAI2BB2XL U1455 ( .B0(n2228), .B1(n2378), .A0N(\register[9][7] ), .A1N(n2381), .Y(n371) );
  OAI2BB2XL U1456 ( .B0(n2225), .B1(n2378), .A0N(\register[9][8] ), .A1N(n2381), .Y(n372) );
  OAI2BB2XL U1457 ( .B0(n2222), .B1(n2378), .A0N(\register[9][9] ), .A1N(n2381), .Y(n373) );
  OAI2BB2XL U1458 ( .B0(n2219), .B1(n2378), .A0N(\register[9][10] ), .A1N(
        n2381), .Y(n374) );
  OAI2BB2XL U1459 ( .B0(n2216), .B1(n2378), .A0N(\register[9][11] ), .A1N(
        n2381), .Y(n375) );
  OAI2BB2XL U1460 ( .B0(n2213), .B1(n2378), .A0N(\register[9][12] ), .A1N(
        n2381), .Y(n376) );
  OAI2BB2XL U1461 ( .B0(n2210), .B1(n2379), .A0N(\register[9][13] ), .A1N(
        n2381), .Y(n377) );
  OAI2BB2XL U1462 ( .B0(n2207), .B1(n2379), .A0N(\register[9][14] ), .A1N(
        n2381), .Y(n378) );
  OAI2BB2XL U1463 ( .B0(n2204), .B1(n2379), .A0N(\register[9][15] ), .A1N(
        n2380), .Y(n379) );
  OAI2BB2XL U1464 ( .B0(n2201), .B1(n2379), .A0N(\register[9][16] ), .A1N(
        n2381), .Y(n380) );
  OAI2BB2XL U1465 ( .B0(n2198), .B1(n2379), .A0N(\register[9][17] ), .A1N(
        n2380), .Y(n381) );
  OAI2BB2XL U1466 ( .B0(n2195), .B1(n2379), .A0N(\register[9][18] ), .A1N(
        n2380), .Y(n382) );
  OAI2BB2XL U1467 ( .B0(n2192), .B1(n2379), .A0N(\register[9][19] ), .A1N(
        n2380), .Y(n383) );
  OAI2BB2XL U1468 ( .B0(n2189), .B1(n2379), .A0N(\register[9][20] ), .A1N(
        n2380), .Y(n384) );
  OAI2BB2XL U1469 ( .B0(n2186), .B1(n2379), .A0N(\register[9][21] ), .A1N(
        n2380), .Y(n385) );
  OAI2BB2XL U1470 ( .B0(n2183), .B1(n2379), .A0N(\register[9][22] ), .A1N(
        n2381), .Y(n386) );
  OAI2BB2XL U1471 ( .B0(n2177), .B1(n2379), .A0N(\register[9][24] ), .A1N(
        n2381), .Y(n388) );
  OAI2BB2XL U1472 ( .B0(n2248), .B1(n2334), .A0N(\register[17][0] ), .A1N(
        n2335), .Y(n620) );
  OAI2BB2XL U1473 ( .B0(n2245), .B1(n2333), .A0N(\register[17][1] ), .A1N(
        n2336), .Y(n621) );
  OAI2BB2XL U1474 ( .B0(n2242), .B1(n2333), .A0N(\register[17][2] ), .A1N(
        n2335), .Y(n622) );
  OAI2BB2XL U1475 ( .B0(n2240), .B1(n2333), .A0N(\register[17][3] ), .A1N(
        n2336), .Y(n623) );
  OAI2BB2XL U1476 ( .B0(n2237), .B1(n2333), .A0N(\register[17][4] ), .A1N(
        n2336), .Y(n624) );
  OAI2BB2XL U1477 ( .B0(n2234), .B1(n2333), .A0N(\register[17][5] ), .A1N(
        n2336), .Y(n625) );
  OAI2BB2XL U1478 ( .B0(n2231), .B1(n2333), .A0N(\register[17][6] ), .A1N(
        n2336), .Y(n626) );
  OAI2BB2XL U1479 ( .B0(n2228), .B1(n2333), .A0N(\register[17][7] ), .A1N(
        n2336), .Y(n627) );
  OAI2BB2XL U1480 ( .B0(n2225), .B1(n2333), .A0N(\register[17][8] ), .A1N(
        n2336), .Y(n628) );
  OAI2BB2XL U1481 ( .B0(n2222), .B1(n2333), .A0N(\register[17][9] ), .A1N(
        n2336), .Y(n629) );
  OAI2BB2XL U1482 ( .B0(n2219), .B1(n2333), .A0N(\register[17][10] ), .A1N(
        n2336), .Y(n630) );
  OAI2BB2XL U1483 ( .B0(n2216), .B1(n2333), .A0N(\register[17][11] ), .A1N(
        n2336), .Y(n631) );
  OAI2BB2XL U1484 ( .B0(n2213), .B1(n2333), .A0N(\register[17][12] ), .A1N(
        n2336), .Y(n632) );
  OAI2BB2XL U1485 ( .B0(n2210), .B1(n2334), .A0N(\register[17][13] ), .A1N(
        n2336), .Y(n633) );
  OAI2BB2XL U1486 ( .B0(n2207), .B1(n2334), .A0N(\register[17][14] ), .A1N(
        n2336), .Y(n634) );
  OAI2BB2XL U1487 ( .B0(n2204), .B1(n2334), .A0N(\register[17][15] ), .A1N(
        n2335), .Y(n635) );
  OAI2BB2XL U1488 ( .B0(n2201), .B1(n2334), .A0N(\register[17][16] ), .A1N(
        n2336), .Y(n636) );
  OAI2BB2XL U1489 ( .B0(n2198), .B1(n2334), .A0N(\register[17][17] ), .A1N(
        n2335), .Y(n637) );
  OAI2BB2XL U1490 ( .B0(n2195), .B1(n2334), .A0N(\register[17][18] ), .A1N(
        n2335), .Y(n638) );
  OAI2BB2XL U1491 ( .B0(n2192), .B1(n2334), .A0N(\register[17][19] ), .A1N(
        n2335), .Y(n639) );
  OAI2BB2XL U1492 ( .B0(n2189), .B1(n2334), .A0N(\register[17][20] ), .A1N(
        n2335), .Y(n640) );
  OAI2BB2XL U1493 ( .B0(n2186), .B1(n2334), .A0N(\register[17][21] ), .A1N(
        n2335), .Y(n641) );
  OAI2BB2XL U1494 ( .B0(n2183), .B1(n2334), .A0N(\register[17][22] ), .A1N(
        n2336), .Y(n642) );
  OAI2BB2XL U1495 ( .B0(n2177), .B1(n2334), .A0N(\register[17][24] ), .A1N(
        n2336), .Y(n644) );
  OAI2BB2XL U1496 ( .B0(n2247), .B1(n2287), .A0N(\register[25][0] ), .A1N(
        n2285), .Y(n876) );
  OAI2BB2XL U1497 ( .B0(n2244), .B1(n2286), .A0N(\register[25][1] ), .A1N(
        n2285), .Y(n877) );
  OAI2BB2XL U1498 ( .B0(n2241), .B1(n2286), .A0N(\register[25][2] ), .A1N(
        n2285), .Y(n878) );
  OAI2BB2XL U1499 ( .B0(n2239), .B1(n2286), .A0N(\register[25][3] ), .A1N(
        n2289), .Y(n879) );
  OAI2BB2XL U1500 ( .B0(n2236), .B1(n2286), .A0N(\register[25][4] ), .A1N(
        n2285), .Y(n880) );
  OAI2BB2XL U1501 ( .B0(n2233), .B1(n2286), .A0N(\register[25][5] ), .A1N(
        n2289), .Y(n881) );
  OAI2BB2XL U1502 ( .B0(n2230), .B1(n2286), .A0N(\register[25][6] ), .A1N(
        n2289), .Y(n882) );
  OAI2BB2XL U1503 ( .B0(n2227), .B1(n2286), .A0N(\register[25][7] ), .A1N(
        n2289), .Y(n883) );
  OAI2BB2XL U1504 ( .B0(n2224), .B1(n2286), .A0N(\register[25][8] ), .A1N(
        n2289), .Y(n884) );
  OAI2BB2XL U1505 ( .B0(n2221), .B1(n2286), .A0N(\register[25][9] ), .A1N(
        n2289), .Y(n885) );
  OAI2BB2XL U1506 ( .B0(n2218), .B1(n2286), .A0N(\register[25][10] ), .A1N(
        n2289), .Y(n886) );
  OAI2BB2XL U1507 ( .B0(n2215), .B1(n2286), .A0N(\register[25][11] ), .A1N(
        n2289), .Y(n887) );
  OAI2BB2XL U1508 ( .B0(n2212), .B1(n2286), .A0N(\register[25][12] ), .A1N(
        n2289), .Y(n888) );
  OAI2BB2XL U1509 ( .B0(n2209), .B1(n2287), .A0N(\register[25][13] ), .A1N(
        n2289), .Y(n889) );
  OAI2BB2XL U1510 ( .B0(n2206), .B1(n2287), .A0N(\register[25][14] ), .A1N(
        n2289), .Y(n890) );
  OAI2BB2XL U1511 ( .B0(n2203), .B1(n2287), .A0N(\register[25][15] ), .A1N(
        n2288), .Y(n891) );
  OAI2BB2XL U1512 ( .B0(n2200), .B1(n2287), .A0N(\register[25][16] ), .A1N(
        n2289), .Y(n892) );
  OAI2BB2XL U1513 ( .B0(n2197), .B1(n2287), .A0N(\register[25][17] ), .A1N(
        n2288), .Y(n893) );
  OAI2BB2XL U1514 ( .B0(n2194), .B1(n2287), .A0N(\register[25][18] ), .A1N(
        n2288), .Y(n894) );
  OAI2BB2XL U1515 ( .B0(n2191), .B1(n2287), .A0N(\register[25][19] ), .A1N(
        n2288), .Y(n895) );
  OAI2BB2XL U1516 ( .B0(n2188), .B1(n2287), .A0N(\register[25][20] ), .A1N(
        n2288), .Y(n896) );
  OAI2BB2XL U1517 ( .B0(n2185), .B1(n2287), .A0N(\register[25][21] ), .A1N(
        n2288), .Y(n897) );
  OAI2BB2XL U1518 ( .B0(n2182), .B1(n2287), .A0N(\register[25][22] ), .A1N(
        n2289), .Y(n898) );
  OAI2BB2XL U1519 ( .B0(n2176), .B1(n2287), .A0N(\register[25][24] ), .A1N(
        n2289), .Y(n900) );
  OAI2BB2XL U1520 ( .B0(n2204), .B1(n2361), .A0N(\register[12][15] ), .A1N(
        n2362), .Y(n475) );
  OAI2BB2XL U1521 ( .B0(n2198), .B1(n2361), .A0N(\register[12][17] ), .A1N(
        n2362), .Y(n477) );
  OAI2BB2XL U1522 ( .B0(n2195), .B1(n2361), .A0N(\register[12][18] ), .A1N(
        n2362), .Y(n478) );
  OAI2BB2XL U1523 ( .B0(n2192), .B1(n2361), .A0N(\register[12][19] ), .A1N(
        n2362), .Y(n479) );
  OAI2BB2XL U1524 ( .B0(n2189), .B1(n2361), .A0N(\register[12][20] ), .A1N(
        n2362), .Y(n480) );
  OAI2BB2XL U1525 ( .B0(n2186), .B1(n2361), .A0N(\register[12][21] ), .A1N(
        n2362), .Y(n481) );
  OAI2BB2XL U1526 ( .B0(n2204), .B1(n2349), .A0N(\register[14][15] ), .A1N(
        n2350), .Y(n539) );
  OAI2BB2XL U1527 ( .B0(n2198), .B1(n2349), .A0N(\register[14][17] ), .A1N(
        n2350), .Y(n541) );
  OAI2BB2XL U1528 ( .B0(n2195), .B1(n2349), .A0N(\register[14][18] ), .A1N(
        n2350), .Y(n542) );
  OAI2BB2XL U1529 ( .B0(n2192), .B1(n2349), .A0N(\register[14][19] ), .A1N(
        n2350), .Y(n543) );
  OAI2BB2XL U1530 ( .B0(n2189), .B1(n2349), .A0N(\register[14][20] ), .A1N(
        n2350), .Y(n544) );
  OAI2BB2XL U1531 ( .B0(n2186), .B1(n2349), .A0N(\register[14][21] ), .A1N(
        n2350), .Y(n545) );
  OAI2BB2XL U1532 ( .B0(n2203), .B1(n2317), .A0N(\register[20][15] ), .A1N(
        n2318), .Y(n731) );
  OAI2BB2XL U1533 ( .B0(n2197), .B1(n2317), .A0N(\register[20][17] ), .A1N(
        n2318), .Y(n733) );
  OAI2BB2XL U1534 ( .B0(n2194), .B1(n2317), .A0N(\register[20][18] ), .A1N(
        n2318), .Y(n734) );
  OAI2BB2XL U1535 ( .B0(n2191), .B1(n2317), .A0N(\register[20][19] ), .A1N(
        n2318), .Y(n735) );
  OAI2BB2XL U1536 ( .B0(n2188), .B1(n2317), .A0N(\register[20][20] ), .A1N(
        n2318), .Y(n736) );
  OAI2BB2XL U1537 ( .B0(n2185), .B1(n2317), .A0N(\register[20][21] ), .A1N(
        n2318), .Y(n737) );
  OAI2BB2XL U1538 ( .B0(n2203), .B1(n2305), .A0N(\register[22][15] ), .A1N(
        n2306), .Y(n795) );
  OAI2BB2XL U1539 ( .B0(n2197), .B1(n2305), .A0N(\register[22][17] ), .A1N(
        n2306), .Y(n797) );
  OAI2BB2XL U1540 ( .B0(n2194), .B1(n2305), .A0N(\register[22][18] ), .A1N(
        n2306), .Y(n798) );
  OAI2BB2XL U1541 ( .B0(n2191), .B1(n2305), .A0N(\register[22][19] ), .A1N(
        n2306), .Y(n799) );
  OAI2BB2XL U1542 ( .B0(n2188), .B1(n2305), .A0N(\register[22][20] ), .A1N(
        n2306), .Y(n800) );
  OAI2BB2XL U1543 ( .B0(n2185), .B1(n2305), .A0N(\register[22][21] ), .A1N(
        n2306), .Y(n801) );
  OAI2BB2XL U1544 ( .B0(n2203), .B1(n2269), .A0N(\register[28][15] ), .A1N(
        n2270), .Y(n987) );
  OAI2BB2XL U1545 ( .B0(n2197), .B1(n2269), .A0N(\register[28][17] ), .A1N(
        n2270), .Y(n989) );
  OAI2BB2XL U1546 ( .B0(n2194), .B1(n2269), .A0N(\register[28][18] ), .A1N(
        n2270), .Y(n990) );
  OAI2BB2XL U1547 ( .B0(n2191), .B1(n2269), .A0N(\register[28][19] ), .A1N(
        n2270), .Y(n991) );
  OAI2BB2XL U1548 ( .B0(n2188), .B1(n2269), .A0N(\register[28][20] ), .A1N(
        n2270), .Y(n992) );
  OAI2BB2XL U1549 ( .B0(n2185), .B1(n2269), .A0N(\register[28][21] ), .A1N(
        n2270), .Y(n993) );
  OAI2BB2XL U1550 ( .B0(n2203), .B1(n2259), .A0N(\register[30][15] ), .A1N(
        n2260), .Y(n1051) );
  OAI2BB2XL U1551 ( .B0(n2197), .B1(n2259), .A0N(\register[30][17] ), .A1N(
        n2260), .Y(n1053) );
  OAI2BB2XL U1552 ( .B0(n2194), .B1(n2259), .A0N(\register[30][18] ), .A1N(
        n2260), .Y(n1054) );
  OAI2BB2XL U1553 ( .B0(n2191), .B1(n2259), .A0N(\register[30][19] ), .A1N(
        n2260), .Y(n1055) );
  OAI2BB2XL U1554 ( .B0(n2188), .B1(n2259), .A0N(\register[30][20] ), .A1N(
        n2260), .Y(n1056) );
  OAI2BB2XL U1555 ( .B0(n2185), .B1(n2259), .A0N(\register[30][21] ), .A1N(
        n2260), .Y(n1057) );
  OAI2BB2XL U1556 ( .B0(n2240), .B1(n2360), .A0N(\register[12][3] ), .A1N(
        n2363), .Y(n463) );
  OAI2BB2XL U1557 ( .B0(n2234), .B1(n2360), .A0N(\register[12][5] ), .A1N(
        n2363), .Y(n465) );
  OAI2BB2XL U1558 ( .B0(n2231), .B1(n2360), .A0N(\register[12][6] ), .A1N(
        n2363), .Y(n466) );
  OAI2BB2XL U1559 ( .B0(n2228), .B1(n2360), .A0N(\register[12][7] ), .A1N(
        n2363), .Y(n467) );
  OAI2BB2XL U1560 ( .B0(n2225), .B1(n2360), .A0N(\register[12][8] ), .A1N(
        n2363), .Y(n468) );
  OAI2BB2XL U1561 ( .B0(n2222), .B1(n2360), .A0N(\register[12][9] ), .A1N(
        n2363), .Y(n469) );
  OAI2BB2XL U1562 ( .B0(n2219), .B1(n2360), .A0N(\register[12][10] ), .A1N(
        n2363), .Y(n470) );
  OAI2BB2XL U1563 ( .B0(n2216), .B1(n2360), .A0N(\register[12][11] ), .A1N(
        n2363), .Y(n471) );
  OAI2BB2XL U1564 ( .B0(n2213), .B1(n2360), .A0N(\register[12][12] ), .A1N(
        n2363), .Y(n472) );
  OAI2BB2XL U1565 ( .B0(n2210), .B1(n2361), .A0N(\register[12][13] ), .A1N(
        n2363), .Y(n473) );
  OAI2BB2XL U1566 ( .B0(n2207), .B1(n2361), .A0N(\register[12][14] ), .A1N(
        n2363), .Y(n474) );
  OAI2BB2XL U1567 ( .B0(n2201), .B1(n2361), .A0N(\register[12][16] ), .A1N(
        n2363), .Y(n476) );
  OAI2BB2XL U1568 ( .B0(n2183), .B1(n2361), .A0N(\register[12][22] ), .A1N(
        n2363), .Y(n482) );
  OAI2BB2XL U1569 ( .B0(n2177), .B1(n2361), .A0N(\register[12][24] ), .A1N(
        n2363), .Y(n484) );
  OAI2BB2XL U1570 ( .B0(n2240), .B1(n2348), .A0N(\register[14][3] ), .A1N(
        n2351), .Y(n527) );
  OAI2BB2XL U1571 ( .B0(n2234), .B1(n2348), .A0N(\register[14][5] ), .A1N(
        n2351), .Y(n529) );
  OAI2BB2XL U1572 ( .B0(n2231), .B1(n2348), .A0N(\register[14][6] ), .A1N(
        n2351), .Y(n530) );
  OAI2BB2XL U1573 ( .B0(n2228), .B1(n2348), .A0N(\register[14][7] ), .A1N(
        n2351), .Y(n531) );
  OAI2BB2XL U1574 ( .B0(n2225), .B1(n2348), .A0N(\register[14][8] ), .A1N(
        n2351), .Y(n532) );
  OAI2BB2XL U1575 ( .B0(n2222), .B1(n2348), .A0N(\register[14][9] ), .A1N(
        n2351), .Y(n533) );
  OAI2BB2XL U1576 ( .B0(n2219), .B1(n2348), .A0N(\register[14][10] ), .A1N(
        n2351), .Y(n534) );
  OAI2BB2XL U1577 ( .B0(n2216), .B1(n2348), .A0N(\register[14][11] ), .A1N(
        n2351), .Y(n535) );
  OAI2BB2XL U1578 ( .B0(n2213), .B1(n2348), .A0N(\register[14][12] ), .A1N(
        n2351), .Y(n536) );
  OAI2BB2XL U1579 ( .B0(n2210), .B1(n2349), .A0N(\register[14][13] ), .A1N(
        n2351), .Y(n537) );
  OAI2BB2XL U1580 ( .B0(n2207), .B1(n2349), .A0N(\register[14][14] ), .A1N(
        n2351), .Y(n538) );
  OAI2BB2XL U1581 ( .B0(n2201), .B1(n2349), .A0N(\register[14][16] ), .A1N(
        n2351), .Y(n540) );
  OAI2BB2XL U1582 ( .B0(n2183), .B1(n2349), .A0N(\register[14][22] ), .A1N(
        n2351), .Y(n546) );
  OAI2BB2XL U1583 ( .B0(n2177), .B1(n2349), .A0N(\register[14][24] ), .A1N(
        n2351), .Y(n548) );
  OAI2BB2XL U1584 ( .B0(n2239), .B1(n2316), .A0N(\register[20][3] ), .A1N(
        n2319), .Y(n719) );
  OAI2BB2XL U1585 ( .B0(n2233), .B1(n2316), .A0N(\register[20][5] ), .A1N(
        n2319), .Y(n721) );
  OAI2BB2XL U1586 ( .B0(n2230), .B1(n2316), .A0N(\register[20][6] ), .A1N(
        n2319), .Y(n722) );
  OAI2BB2XL U1587 ( .B0(n2227), .B1(n2316), .A0N(\register[20][7] ), .A1N(
        n2319), .Y(n723) );
  OAI2BB2XL U1588 ( .B0(n2224), .B1(n2316), .A0N(\register[20][8] ), .A1N(
        n2319), .Y(n724) );
  OAI2BB2XL U1589 ( .B0(n2221), .B1(n2316), .A0N(\register[20][9] ), .A1N(
        n2319), .Y(n725) );
  OAI2BB2XL U1590 ( .B0(n2218), .B1(n2316), .A0N(\register[20][10] ), .A1N(
        n2319), .Y(n726) );
  OAI2BB2XL U1591 ( .B0(n2215), .B1(n2316), .A0N(\register[20][11] ), .A1N(
        n2319), .Y(n727) );
  OAI2BB2XL U1592 ( .B0(n2212), .B1(n2316), .A0N(\register[20][12] ), .A1N(
        n2319), .Y(n728) );
  OAI2BB2XL U1593 ( .B0(n2209), .B1(n2317), .A0N(\register[20][13] ), .A1N(
        n2319), .Y(n729) );
  OAI2BB2XL U1594 ( .B0(n2206), .B1(n2317), .A0N(\register[20][14] ), .A1N(
        n2319), .Y(n730) );
  OAI2BB2XL U1595 ( .B0(n2200), .B1(n2317), .A0N(\register[20][16] ), .A1N(
        n2319), .Y(n732) );
  OAI2BB2XL U1596 ( .B0(n2182), .B1(n2317), .A0N(\register[20][22] ), .A1N(
        n2319), .Y(n738) );
  OAI2BB2XL U1597 ( .B0(n2176), .B1(n2317), .A0N(\register[20][24] ), .A1N(
        n2319), .Y(n740) );
  OAI2BB2XL U1598 ( .B0(n2239), .B1(n2304), .A0N(\register[22][3] ), .A1N(
        n2307), .Y(n783) );
  OAI2BB2XL U1599 ( .B0(n2233), .B1(n2304), .A0N(\register[22][5] ), .A1N(
        n2307), .Y(n785) );
  OAI2BB2XL U1600 ( .B0(n2230), .B1(n2304), .A0N(\register[22][6] ), .A1N(
        n2307), .Y(n786) );
  OAI2BB2XL U1601 ( .B0(n2227), .B1(n2304), .A0N(\register[22][7] ), .A1N(
        n2307), .Y(n787) );
  OAI2BB2XL U1602 ( .B0(n2224), .B1(n2304), .A0N(\register[22][8] ), .A1N(
        n2307), .Y(n788) );
  OAI2BB2XL U1603 ( .B0(n2221), .B1(n2304), .A0N(\register[22][9] ), .A1N(
        n2307), .Y(n789) );
  OAI2BB2XL U1604 ( .B0(n2218), .B1(n2304), .A0N(\register[22][10] ), .A1N(
        n2307), .Y(n790) );
  OAI2BB2XL U1605 ( .B0(n2215), .B1(n2304), .A0N(\register[22][11] ), .A1N(
        n2307), .Y(n791) );
  OAI2BB2XL U1606 ( .B0(n2212), .B1(n2304), .A0N(\register[22][12] ), .A1N(
        n2307), .Y(n792) );
  OAI2BB2XL U1607 ( .B0(n2209), .B1(n2305), .A0N(\register[22][13] ), .A1N(
        n2307), .Y(n793) );
  OAI2BB2XL U1608 ( .B0(n2206), .B1(n2305), .A0N(\register[22][14] ), .A1N(
        n2307), .Y(n794) );
  OAI2BB2XL U1609 ( .B0(n2200), .B1(n2305), .A0N(\register[22][16] ), .A1N(
        n2307), .Y(n796) );
  OAI2BB2XL U1610 ( .B0(n2182), .B1(n2305), .A0N(\register[22][22] ), .A1N(
        n2307), .Y(n802) );
  OAI2BB2XL U1611 ( .B0(n2176), .B1(n2305), .A0N(\register[22][24] ), .A1N(
        n2307), .Y(n804) );
  OAI2BB2XL U1612 ( .B0(n2239), .B1(n2268), .A0N(\register[28][3] ), .A1N(
        n2271), .Y(n975) );
  OAI2BB2XL U1613 ( .B0(n2233), .B1(n2268), .A0N(\register[28][5] ), .A1N(
        n2271), .Y(n977) );
  OAI2BB2XL U1614 ( .B0(n2230), .B1(n2268), .A0N(\register[28][6] ), .A1N(
        n2271), .Y(n978) );
  OAI2BB2XL U1615 ( .B0(n2227), .B1(n2268), .A0N(\register[28][7] ), .A1N(
        n2271), .Y(n979) );
  OAI2BB2XL U1616 ( .B0(n2224), .B1(n2268), .A0N(\register[28][8] ), .A1N(
        n2271), .Y(n980) );
  OAI2BB2XL U1617 ( .B0(n2221), .B1(n2268), .A0N(\register[28][9] ), .A1N(
        n2271), .Y(n981) );
  OAI2BB2XL U1618 ( .B0(n2218), .B1(n2268), .A0N(\register[28][10] ), .A1N(
        n2271), .Y(n982) );
  OAI2BB2XL U1619 ( .B0(n2215), .B1(n2268), .A0N(\register[28][11] ), .A1N(
        n2271), .Y(n983) );
  OAI2BB2XL U1620 ( .B0(n2212), .B1(n2268), .A0N(\register[28][12] ), .A1N(
        n2271), .Y(n984) );
  OAI2BB2XL U1621 ( .B0(n2209), .B1(n2269), .A0N(\register[28][13] ), .A1N(
        n2271), .Y(n985) );
  OAI2BB2XL U1622 ( .B0(n2206), .B1(n2269), .A0N(\register[28][14] ), .A1N(
        n2271), .Y(n986) );
  OAI2BB2XL U1623 ( .B0(n2200), .B1(n2269), .A0N(\register[28][16] ), .A1N(
        n2271), .Y(n988) );
  OAI2BB2XL U1624 ( .B0(n2182), .B1(n2269), .A0N(\register[28][22] ), .A1N(
        n2271), .Y(n994) );
  OAI2BB2XL U1625 ( .B0(n2176), .B1(n2269), .A0N(\register[28][24] ), .A1N(
        n2271), .Y(n996) );
  OAI2BB2XL U1626 ( .B0(n2239), .B1(n2258), .A0N(\register[30][3] ), .A1N(
        n2261), .Y(n1039) );
  OAI2BB2XL U1627 ( .B0(n2233), .B1(n2258), .A0N(\register[30][5] ), .A1N(
        n2261), .Y(n1041) );
  OAI2BB2XL U1628 ( .B0(n2230), .B1(n2258), .A0N(\register[30][6] ), .A1N(
        n2261), .Y(n1042) );
  OAI2BB2XL U1629 ( .B0(n2227), .B1(n2258), .A0N(\register[30][7] ), .A1N(
        n2261), .Y(n1043) );
  OAI2BB2XL U1630 ( .B0(n2224), .B1(n2258), .A0N(\register[30][8] ), .A1N(
        n2261), .Y(n1044) );
  OAI2BB2XL U1631 ( .B0(n2221), .B1(n2258), .A0N(\register[30][9] ), .A1N(
        n2261), .Y(n1045) );
  OAI2BB2XL U1632 ( .B0(n2218), .B1(n2258), .A0N(\register[30][10] ), .A1N(
        n2261), .Y(n1046) );
  OAI2BB2XL U1633 ( .B0(n2215), .B1(n2258), .A0N(\register[30][11] ), .A1N(
        n2261), .Y(n1047) );
  OAI2BB2XL U1634 ( .B0(n2212), .B1(n2258), .A0N(\register[30][12] ), .A1N(
        n2261), .Y(n1048) );
  OAI2BB2XL U1635 ( .B0(n2209), .B1(n2259), .A0N(\register[30][13] ), .A1N(
        n2261), .Y(n1049) );
  OAI2BB2XL U1636 ( .B0(n2206), .B1(n2259), .A0N(\register[30][14] ), .A1N(
        n2261), .Y(n1050) );
  OAI2BB2XL U1637 ( .B0(n2200), .B1(n2259), .A0N(\register[30][16] ), .A1N(
        n2261), .Y(n1052) );
  OAI2BB2XL U1638 ( .B0(n2182), .B1(n2259), .A0N(\register[30][22] ), .A1N(
        n2261), .Y(n1058) );
  OAI2BB2XL U1639 ( .B0(n2176), .B1(n2259), .A0N(\register[30][24] ), .A1N(
        n2261), .Y(n1060) );
  OAI2BB2XL U1640 ( .B0(n2248), .B1(n2361), .A0N(\register[12][0] ), .A1N(
        n2358), .Y(n460) );
  OAI2BB2XL U1641 ( .B0(n2245), .B1(n2360), .A0N(\register[12][1] ), .A1N(
        n2358), .Y(n461) );
  OAI2BB2XL U1642 ( .B0(n2242), .B1(n2360), .A0N(\register[12][2] ), .A1N(
        n2358), .Y(n462) );
  OAI2BB2XL U1643 ( .B0(n2237), .B1(n2360), .A0N(\register[12][4] ), .A1N(
        n2358), .Y(n464) );
  OAI2BB2XL U1644 ( .B0(n2248), .B1(n2349), .A0N(\register[14][0] ), .A1N(
        n2350), .Y(n524) );
  OAI2BB2XL U1645 ( .B0(n2245), .B1(n2348), .A0N(\register[14][1] ), .A1N(
        n2350), .Y(n525) );
  OAI2BB2XL U1646 ( .B0(n2242), .B1(n2348), .A0N(\register[14][2] ), .A1N(
        n2350), .Y(n526) );
  OAI2BB2XL U1647 ( .B0(n2237), .B1(n2348), .A0N(\register[14][4] ), .A1N(
        n2350), .Y(n528) );
  OAI2BB2XL U1648 ( .B0(n2247), .B1(n2317), .A0N(\register[20][0] ), .A1N(
        n2314), .Y(n716) );
  OAI2BB2XL U1649 ( .B0(n2244), .B1(n2316), .A0N(\register[20][1] ), .A1N(
        n2314), .Y(n717) );
  OAI2BB2XL U1650 ( .B0(n2241), .B1(n2316), .A0N(\register[20][2] ), .A1N(
        n2314), .Y(n718) );
  OAI2BB2XL U1651 ( .B0(n2236), .B1(n2316), .A0N(\register[20][4] ), .A1N(
        n2314), .Y(n720) );
  OAI2BB2XL U1652 ( .B0(n2247), .B1(n2305), .A0N(\register[22][0] ), .A1N(
        n2302), .Y(n780) );
  OAI2BB2XL U1653 ( .B0(n2244), .B1(n2304), .A0N(\register[22][1] ), .A1N(
        n2302), .Y(n781) );
  OAI2BB2XL U1654 ( .B0(n2241), .B1(n2304), .A0N(\register[22][2] ), .A1N(
        n2302), .Y(n782) );
  OAI2BB2XL U1655 ( .B0(n2236), .B1(n2304), .A0N(\register[22][4] ), .A1N(
        n2302), .Y(n784) );
  OAI2BB2XL U1656 ( .B0(n2247), .B1(n2269), .A0N(\register[28][0] ), .A1N(
        n2267), .Y(n972) );
  OAI2BB2XL U1657 ( .B0(n2244), .B1(n2268), .A0N(\register[28][1] ), .A1N(
        n2267), .Y(n973) );
  OAI2BB2XL U1658 ( .B0(n2241), .B1(n2268), .A0N(\register[28][2] ), .A1N(
        n2267), .Y(n974) );
  OAI2BB2XL U1659 ( .B0(n2236), .B1(n2268), .A0N(\register[28][4] ), .A1N(
        n2267), .Y(n976) );
  OAI2BB2XL U1660 ( .B0(n2247), .B1(n2259), .A0N(\register[30][0] ), .A1N(
        n2257), .Y(n1036) );
  OAI2BB2XL U1661 ( .B0(n2244), .B1(n2258), .A0N(\register[30][1] ), .A1N(
        n2257), .Y(n1037) );
  OAI2BB2XL U1662 ( .B0(n2241), .B1(n2258), .A0N(\register[30][2] ), .A1N(
        n2257), .Y(n1038) );
  OAI2BB2XL U1663 ( .B0(n2236), .B1(n2258), .A0N(\register[30][4] ), .A1N(
        n2257), .Y(n1040) );
  OAI2BB2XL U1664 ( .B0(n2248), .B1(n2385), .A0N(\register[8][0] ), .A1N(n2382), .Y(n332) );
  OAI2BB2XL U1665 ( .B0(n2245), .B1(n2384), .A0N(\register[8][1] ), .A1N(n2382), .Y(n333) );
  OAI2BB2XL U1666 ( .B0(n2242), .B1(n2384), .A0N(\register[8][2] ), .A1N(n2382), .Y(n334) );
  OAI2BB2XL U1667 ( .B0(n2240), .B1(n2384), .A0N(\register[8][3] ), .A1N(n2387), .Y(n335) );
  OAI2BB2XL U1668 ( .B0(n2237), .B1(n2384), .A0N(\register[8][4] ), .A1N(n2382), .Y(n336) );
  OAI2BB2XL U1669 ( .B0(n2234), .B1(n2384), .A0N(\register[8][5] ), .A1N(n2387), .Y(n337) );
  OAI2BB2XL U1670 ( .B0(n2231), .B1(n2384), .A0N(\register[8][6] ), .A1N(n2387), .Y(n338) );
  OAI2BB2XL U1671 ( .B0(n2228), .B1(n2384), .A0N(\register[8][7] ), .A1N(n2387), .Y(n339) );
  OAI2BB2XL U1672 ( .B0(n2225), .B1(n2384), .A0N(\register[8][8] ), .A1N(n2387), .Y(n340) );
  OAI2BB2XL U1673 ( .B0(n2222), .B1(n2384), .A0N(\register[8][9] ), .A1N(n2387), .Y(n341) );
  OAI2BB2XL U1674 ( .B0(n2219), .B1(n2384), .A0N(\register[8][10] ), .A1N(
        n2387), .Y(n342) );
  OAI2BB2XL U1675 ( .B0(n2216), .B1(n2384), .A0N(\register[8][11] ), .A1N(
        n2387), .Y(n343) );
  OAI2BB2XL U1676 ( .B0(n2213), .B1(n2384), .A0N(\register[8][12] ), .A1N(
        n2387), .Y(n344) );
  OAI2BB2XL U1677 ( .B0(n2210), .B1(n2385), .A0N(\register[8][13] ), .A1N(
        n2387), .Y(n345) );
  OAI2BB2XL U1678 ( .B0(n2207), .B1(n2385), .A0N(\register[8][14] ), .A1N(
        n2387), .Y(n346) );
  OAI2BB2XL U1679 ( .B0(n2204), .B1(n2385), .A0N(\register[8][15] ), .A1N(
        n2386), .Y(n347) );
  OAI2BB2XL U1680 ( .B0(n2201), .B1(n2385), .A0N(\register[8][16] ), .A1N(
        n2387), .Y(n348) );
  OAI2BB2XL U1681 ( .B0(n2198), .B1(n2385), .A0N(\register[8][17] ), .A1N(
        n2386), .Y(n349) );
  OAI2BB2XL U1682 ( .B0(n2195), .B1(n2385), .A0N(\register[8][18] ), .A1N(
        n2386), .Y(n350) );
  OAI2BB2XL U1683 ( .B0(n2192), .B1(n2385), .A0N(\register[8][19] ), .A1N(
        n2386), .Y(n351) );
  OAI2BB2XL U1684 ( .B0(n2189), .B1(n2385), .A0N(\register[8][20] ), .A1N(
        n2386), .Y(n352) );
  OAI2BB2XL U1685 ( .B0(n2186), .B1(n2385), .A0N(\register[8][21] ), .A1N(
        n2386), .Y(n353) );
  OAI2BB2XL U1686 ( .B0(n2183), .B1(n2385), .A0N(\register[8][22] ), .A1N(
        n2387), .Y(n354) );
  OAI2BB2XL U1687 ( .B0(n2177), .B1(n2385), .A0N(\register[8][24] ), .A1N(
        n2387), .Y(n356) );
  OAI2BB2XL U1688 ( .B0(n2248), .B1(n2338), .A0N(\register[16][0] ), .A1N(
        n2338), .Y(n588) );
  OAI2BB2XL U1689 ( .B0(n2245), .B1(n2339), .A0N(\register[16][1] ), .A1N(
        n2338), .Y(n589) );
  OAI2BB2XL U1690 ( .B0(n2242), .B1(n2339), .A0N(\register[16][2] ), .A1N(
        n2338), .Y(n590) );
  OAI2BB2XL U1691 ( .B0(n2240), .B1(n2339), .A0N(\register[16][3] ), .A1N(
        n2341), .Y(n591) );
  OAI2BB2XL U1692 ( .B0(n2237), .B1(n2339), .A0N(\register[16][4] ), .A1N(
        n2338), .Y(n592) );
  OAI2BB2XL U1693 ( .B0(n2234), .B1(n2339), .A0N(\register[16][5] ), .A1N(
        n2341), .Y(n593) );
  OAI2BB2XL U1694 ( .B0(n2231), .B1(n2339), .A0N(\register[16][6] ), .A1N(
        n2341), .Y(n594) );
  OAI2BB2XL U1695 ( .B0(n2228), .B1(n2339), .A0N(\register[16][7] ), .A1N(
        n2341), .Y(n595) );
  OAI2BB2XL U1696 ( .B0(n2225), .B1(n2339), .A0N(\register[16][8] ), .A1N(
        n2341), .Y(n596) );
  OAI2BB2XL U1697 ( .B0(n2222), .B1(n2339), .A0N(\register[16][9] ), .A1N(
        n2341), .Y(n597) );
  OAI2BB2XL U1698 ( .B0(n2219), .B1(n2339), .A0N(\register[16][10] ), .A1N(
        n2341), .Y(n598) );
  OAI2BB2XL U1699 ( .B0(n2216), .B1(n2339), .A0N(\register[16][11] ), .A1N(
        n2341), .Y(n599) );
  OAI2BB2XL U1700 ( .B0(n2213), .B1(n2339), .A0N(\register[16][12] ), .A1N(
        n2341), .Y(n600) );
  OAI2BB2XL U1701 ( .B0(n2210), .B1(n2338), .A0N(\register[16][13] ), .A1N(
        n2341), .Y(n601) );
  OAI2BB2XL U1702 ( .B0(n2207), .B1(n2338), .A0N(\register[16][14] ), .A1N(
        n2341), .Y(n602) );
  OAI2BB2XL U1703 ( .B0(n2204), .B1(n2338), .A0N(\register[16][15] ), .A1N(
        n2340), .Y(n603) );
  OAI2BB2XL U1704 ( .B0(n2201), .B1(n2338), .A0N(\register[16][16] ), .A1N(
        n2341), .Y(n604) );
  OAI2BB2XL U1705 ( .B0(n2198), .B1(n2338), .A0N(\register[16][17] ), .A1N(
        n2340), .Y(n605) );
  OAI2BB2XL U1706 ( .B0(n2195), .B1(n2339), .A0N(\register[16][18] ), .A1N(
        n2340), .Y(n606) );
  OAI2BB2XL U1707 ( .B0(n2192), .B1(n2338), .A0N(\register[16][19] ), .A1N(
        n2340), .Y(n607) );
  OAI2BB2XL U1708 ( .B0(n2189), .B1(n2339), .A0N(\register[16][20] ), .A1N(
        n2340), .Y(n608) );
  OAI2BB2XL U1709 ( .B0(n2186), .B1(n2338), .A0N(\register[16][21] ), .A1N(
        n2340), .Y(n609) );
  OAI2BB2XL U1710 ( .B0(n2183), .B1(n2339), .A0N(\register[16][22] ), .A1N(
        n2341), .Y(n610) );
  OAI2BB2XL U1711 ( .B0(n2177), .B1(n2339), .A0N(\register[16][24] ), .A1N(
        n2341), .Y(n612) );
  OAI2BB2XL U1712 ( .B0(n2247), .B1(n2293), .A0N(\register[24][0] ), .A1N(
        n2290), .Y(n844) );
  OAI2BB2XL U1713 ( .B0(n2244), .B1(n2292), .A0N(\register[24][1] ), .A1N(
        n2290), .Y(n845) );
  OAI2BB2XL U1714 ( .B0(n2241), .B1(n2292), .A0N(\register[24][2] ), .A1N(
        n2290), .Y(n846) );
  OAI2BB2XL U1715 ( .B0(n2239), .B1(n2292), .A0N(\register[24][3] ), .A1N(
        n2295), .Y(n847) );
  OAI2BB2XL U1716 ( .B0(n2236), .B1(n2292), .A0N(\register[24][4] ), .A1N(
        n2290), .Y(n848) );
  OAI2BB2XL U1717 ( .B0(n2233), .B1(n2292), .A0N(\register[24][5] ), .A1N(
        n2295), .Y(n849) );
  OAI2BB2XL U1718 ( .B0(n2230), .B1(n2292), .A0N(\register[24][6] ), .A1N(
        n2295), .Y(n850) );
  OAI2BB2XL U1719 ( .B0(n2227), .B1(n2292), .A0N(\register[24][7] ), .A1N(
        n2295), .Y(n851) );
  OAI2BB2XL U1720 ( .B0(n2224), .B1(n2292), .A0N(\register[24][8] ), .A1N(
        n2295), .Y(n852) );
  OAI2BB2XL U1721 ( .B0(n2221), .B1(n2292), .A0N(\register[24][9] ), .A1N(
        n2295), .Y(n853) );
  OAI2BB2XL U1722 ( .B0(n2218), .B1(n2292), .A0N(\register[24][10] ), .A1N(
        n2295), .Y(n854) );
  OAI2BB2XL U1723 ( .B0(n2215), .B1(n2292), .A0N(\register[24][11] ), .A1N(
        n2295), .Y(n855) );
  OAI2BB2XL U1724 ( .B0(n2212), .B1(n2292), .A0N(\register[24][12] ), .A1N(
        n2295), .Y(n856) );
  OAI2BB2XL U1725 ( .B0(n2209), .B1(n2293), .A0N(\register[24][13] ), .A1N(
        n2295), .Y(n857) );
  OAI2BB2XL U1726 ( .B0(n2206), .B1(n2293), .A0N(\register[24][14] ), .A1N(
        n2295), .Y(n858) );
  OAI2BB2XL U1727 ( .B0(n2203), .B1(n2293), .A0N(\register[24][15] ), .A1N(
        n2294), .Y(n859) );
  OAI2BB2XL U1728 ( .B0(n2200), .B1(n2293), .A0N(\register[24][16] ), .A1N(
        n2295), .Y(n860) );
  OAI2BB2XL U1729 ( .B0(n2197), .B1(n2293), .A0N(\register[24][17] ), .A1N(
        n2294), .Y(n861) );
  OAI2BB2XL U1730 ( .B0(n2194), .B1(n2293), .A0N(\register[24][18] ), .A1N(
        n2294), .Y(n862) );
  OAI2BB2XL U1731 ( .B0(n2191), .B1(n2293), .A0N(\register[24][19] ), .A1N(
        n2294), .Y(n863) );
  OAI2BB2XL U1732 ( .B0(n2188), .B1(n2293), .A0N(\register[24][20] ), .A1N(
        n2294), .Y(n864) );
  OAI2BB2XL U1733 ( .B0(n2185), .B1(n2293), .A0N(\register[24][21] ), .A1N(
        n2294), .Y(n865) );
  OAI2BB2XL U1734 ( .B0(n2182), .B1(n2293), .A0N(\register[24][22] ), .A1N(
        n2295), .Y(n866) );
  OAI2BB2XL U1735 ( .B0(n2176), .B1(n2293), .A0N(\register[24][24] ), .A1N(
        n2295), .Y(n868) );
  OAI2BB2XL U1736 ( .B0(n2204), .B1(n2355), .A0N(\register[13][15] ), .A1N(
        n2356), .Y(n507) );
  OAI2BB2XL U1737 ( .B0(n2198), .B1(n2355), .A0N(\register[13][17] ), .A1N(
        n2356), .Y(n509) );
  OAI2BB2XL U1738 ( .B0(n2195), .B1(n2355), .A0N(\register[13][18] ), .A1N(
        n2356), .Y(n510) );
  OAI2BB2XL U1739 ( .B0(n2192), .B1(n2355), .A0N(\register[13][19] ), .A1N(
        n2356), .Y(n511) );
  OAI2BB2XL U1740 ( .B0(n2189), .B1(n2355), .A0N(\register[13][20] ), .A1N(
        n2356), .Y(n512) );
  OAI2BB2XL U1741 ( .B0(n2186), .B1(n2355), .A0N(\register[13][21] ), .A1N(
        n2356), .Y(n513) );
  OAI2BB2XL U1742 ( .B0(n2204), .B1(n2345), .A0N(\register[15][15] ), .A1N(
        n2346), .Y(n571) );
  OAI2BB2XL U1743 ( .B0(n2198), .B1(n2345), .A0N(\register[15][17] ), .A1N(
        n2346), .Y(n573) );
  OAI2BB2XL U1744 ( .B0(n2195), .B1(n2345), .A0N(\register[15][18] ), .A1N(
        n2343), .Y(n574) );
  OAI2BB2XL U1745 ( .B0(n2192), .B1(n2345), .A0N(\register[15][19] ), .A1N(
        n2343), .Y(n575) );
  OAI2BB2XL U1746 ( .B0(n2189), .B1(n2345), .A0N(\register[15][20] ), .A1N(
        n2343), .Y(n576) );
  OAI2BB2XL U1747 ( .B0(n2186), .B1(n2345), .A0N(\register[15][21] ), .A1N(
        n2343), .Y(n577) );
  OAI2BB2XL U1748 ( .B0(n2203), .B1(n2311), .A0N(\register[21][15] ), .A1N(
        n2312), .Y(n763) );
  OAI2BB2XL U1749 ( .B0(n2197), .B1(n2311), .A0N(\register[21][17] ), .A1N(
        n2312), .Y(n765) );
  OAI2BB2XL U1750 ( .B0(n2194), .B1(n2311), .A0N(\register[21][18] ), .A1N(
        n2312), .Y(n766) );
  OAI2BB2XL U1751 ( .B0(n2191), .B1(n2311), .A0N(\register[21][19] ), .A1N(
        n2312), .Y(n767) );
  OAI2BB2XL U1752 ( .B0(n2188), .B1(n2311), .A0N(\register[21][20] ), .A1N(
        n2312), .Y(n768) );
  OAI2BB2XL U1753 ( .B0(n2185), .B1(n2311), .A0N(\register[21][21] ), .A1N(
        n2312), .Y(n769) );
  OAI2BB2XL U1754 ( .B0(n2203), .B1(n2299), .A0N(\register[23][15] ), .A1N(
        n2300), .Y(n827) );
  OAI2BB2XL U1755 ( .B0(n2197), .B1(n2299), .A0N(\register[23][17] ), .A1N(
        n2300), .Y(n829) );
  OAI2BB2XL U1756 ( .B0(n2194), .B1(n2299), .A0N(\register[23][18] ), .A1N(
        n2300), .Y(n830) );
  OAI2BB2XL U1757 ( .B0(n2191), .B1(n2299), .A0N(\register[23][19] ), .A1N(
        n2300), .Y(n831) );
  OAI2BB2XL U1758 ( .B0(n2188), .B1(n2299), .A0N(\register[23][20] ), .A1N(
        n2300), .Y(n832) );
  OAI2BB2XL U1759 ( .B0(n2185), .B1(n2299), .A0N(\register[23][21] ), .A1N(
        n2300), .Y(n833) );
  OAI2BB2XL U1760 ( .B0(n2203), .B1(n2263), .A0N(\register[29][15] ), .A1N(
        n2264), .Y(n1019) );
  OAI2BB2XL U1761 ( .B0(n2197), .B1(n2263), .A0N(\register[29][17] ), .A1N(
        n2264), .Y(n1021) );
  OAI2BB2XL U1762 ( .B0(n2194), .B1(n2263), .A0N(\register[29][18] ), .A1N(
        n2264), .Y(n1022) );
  OAI2BB2XL U1763 ( .B0(n2191), .B1(n2263), .A0N(\register[29][19] ), .A1N(
        n2264), .Y(n1023) );
  OAI2BB2XL U1764 ( .B0(n2188), .B1(n2263), .A0N(\register[29][20] ), .A1N(
        n2264), .Y(n1024) );
  OAI2BB2XL U1765 ( .B0(n2185), .B1(n2263), .A0N(\register[29][21] ), .A1N(
        n2264), .Y(n1025) );
  OAI2BB2XL U1766 ( .B0(n2203), .B1(n2253), .A0N(\register[31][15] ), .A1N(
        n2254), .Y(n1083) );
  OAI2BB2XL U1767 ( .B0(n2197), .B1(n2253), .A0N(\register[31][17] ), .A1N(
        n2254), .Y(n1085) );
  OAI2BB2XL U1768 ( .B0(n2194), .B1(n2253), .A0N(\register[31][18] ), .A1N(
        n2254), .Y(n1086) );
  OAI2BB2XL U1769 ( .B0(n2191), .B1(n2253), .A0N(\register[31][19] ), .A1N(
        n2254), .Y(n1087) );
  OAI2BB2XL U1770 ( .B0(n2188), .B1(n2253), .A0N(\register[31][20] ), .A1N(
        n2254), .Y(n1088) );
  OAI2BB2XL U1771 ( .B0(n2185), .B1(n2253), .A0N(\register[31][21] ), .A1N(
        n2254), .Y(n1089) );
  OAI2BB2XL U1772 ( .B0(n2240), .B1(n2354), .A0N(\register[13][3] ), .A1N(
        n2357), .Y(n495) );
  OAI2BB2XL U1773 ( .B0(n2234), .B1(n2354), .A0N(\register[13][5] ), .A1N(
        n2357), .Y(n497) );
  OAI2BB2XL U1774 ( .B0(n2231), .B1(n2354), .A0N(\register[13][6] ), .A1N(
        n2357), .Y(n498) );
  OAI2BB2XL U1775 ( .B0(n2228), .B1(n2354), .A0N(\register[13][7] ), .A1N(
        n2357), .Y(n499) );
  OAI2BB2XL U1776 ( .B0(n2225), .B1(n2354), .A0N(\register[13][8] ), .A1N(
        n2357), .Y(n500) );
  OAI2BB2XL U1777 ( .B0(n2222), .B1(n2354), .A0N(\register[13][9] ), .A1N(
        n2357), .Y(n501) );
  OAI2BB2XL U1778 ( .B0(n2219), .B1(n2354), .A0N(\register[13][10] ), .A1N(
        n2357), .Y(n502) );
  OAI2BB2XL U1779 ( .B0(n2216), .B1(n2354), .A0N(\register[13][11] ), .A1N(
        n2357), .Y(n503) );
  OAI2BB2XL U1780 ( .B0(n2213), .B1(n2354), .A0N(\register[13][12] ), .A1N(
        n2357), .Y(n504) );
  OAI2BB2XL U1781 ( .B0(n2210), .B1(n2355), .A0N(\register[13][13] ), .A1N(
        n2357), .Y(n505) );
  OAI2BB2XL U1782 ( .B0(n2207), .B1(n2355), .A0N(\register[13][14] ), .A1N(
        n2357), .Y(n506) );
  OAI2BB2XL U1783 ( .B0(n2201), .B1(n2355), .A0N(\register[13][16] ), .A1N(
        n2357), .Y(n508) );
  OAI2BB2XL U1784 ( .B0(n2183), .B1(n2355), .A0N(\register[13][22] ), .A1N(
        n2357), .Y(n514) );
  OAI2BB2XL U1785 ( .B0(n2177), .B1(n2355), .A0N(\register[13][24] ), .A1N(
        n2357), .Y(n516) );
  OAI2BB2XL U1786 ( .B0(n2240), .B1(n2344), .A0N(\register[15][3] ), .A1N(
        n2346), .Y(n559) );
  OAI2BB2XL U1787 ( .B0(n2234), .B1(n2344), .A0N(\register[15][5] ), .A1N(
        n2346), .Y(n561) );
  OAI2BB2XL U1788 ( .B0(n2231), .B1(n2344), .A0N(\register[15][6] ), .A1N(
        n2346), .Y(n562) );
  OAI2BB2XL U1789 ( .B0(n2228), .B1(n2344), .A0N(\register[15][7] ), .A1N(
        n2346), .Y(n563) );
  OAI2BB2XL U1790 ( .B0(n2225), .B1(n2344), .A0N(\register[15][8] ), .A1N(
        n2346), .Y(n564) );
  OAI2BB2XL U1791 ( .B0(n2222), .B1(n2344), .A0N(\register[15][9] ), .A1N(
        n2346), .Y(n565) );
  OAI2BB2XL U1792 ( .B0(n2219), .B1(n2344), .A0N(\register[15][10] ), .A1N(
        n2346), .Y(n566) );
  OAI2BB2XL U1793 ( .B0(n2216), .B1(n2344), .A0N(\register[15][11] ), .A1N(
        n2346), .Y(n567) );
  OAI2BB2XL U1794 ( .B0(n2213), .B1(n2344), .A0N(\register[15][12] ), .A1N(
        n2346), .Y(n568) );
  OAI2BB2XL U1795 ( .B0(n2210), .B1(n2345), .A0N(\register[15][13] ), .A1N(
        n2346), .Y(n569) );
  OAI2BB2XL U1796 ( .B0(n2207), .B1(n2345), .A0N(\register[15][14] ), .A1N(
        n2346), .Y(n570) );
  OAI2BB2XL U1797 ( .B0(n2201), .B1(n2345), .A0N(\register[15][16] ), .A1N(
        n2346), .Y(n572) );
  OAI2BB2XL U1798 ( .B0(n2183), .B1(n2345), .A0N(\register[15][22] ), .A1N(
        n2346), .Y(n578) );
  OAI2BB2XL U1799 ( .B0(n2177), .B1(n2345), .A0N(\register[15][24] ), .A1N(
        n2346), .Y(n580) );
  OAI2BB2XL U1800 ( .B0(n2239), .B1(n2310), .A0N(\register[21][3] ), .A1N(
        n2313), .Y(n751) );
  OAI2BB2XL U1801 ( .B0(n2233), .B1(n2310), .A0N(\register[21][5] ), .A1N(
        n2313), .Y(n753) );
  OAI2BB2XL U1802 ( .B0(n2230), .B1(n2310), .A0N(\register[21][6] ), .A1N(
        n2313), .Y(n754) );
  OAI2BB2XL U1803 ( .B0(n2227), .B1(n2310), .A0N(\register[21][7] ), .A1N(
        n2313), .Y(n755) );
  OAI2BB2XL U1804 ( .B0(n2224), .B1(n2310), .A0N(\register[21][8] ), .A1N(
        n2313), .Y(n756) );
  OAI2BB2XL U1805 ( .B0(n2221), .B1(n2310), .A0N(\register[21][9] ), .A1N(
        n2313), .Y(n757) );
  OAI2BB2XL U1806 ( .B0(n2218), .B1(n2310), .A0N(\register[21][10] ), .A1N(
        n2313), .Y(n758) );
  OAI2BB2XL U1807 ( .B0(n2215), .B1(n2310), .A0N(\register[21][11] ), .A1N(
        n2313), .Y(n759) );
  OAI2BB2XL U1808 ( .B0(n2212), .B1(n2310), .A0N(\register[21][12] ), .A1N(
        n2313), .Y(n760) );
  OAI2BB2XL U1809 ( .B0(n2209), .B1(n2311), .A0N(\register[21][13] ), .A1N(
        n2313), .Y(n761) );
  OAI2BB2XL U1810 ( .B0(n2206), .B1(n2311), .A0N(\register[21][14] ), .A1N(
        n2313), .Y(n762) );
  OAI2BB2XL U1811 ( .B0(n2200), .B1(n2311), .A0N(\register[21][16] ), .A1N(
        n2313), .Y(n764) );
  OAI2BB2XL U1812 ( .B0(n2182), .B1(n2311), .A0N(\register[21][22] ), .A1N(
        n2313), .Y(n770) );
  OAI2BB2XL U1813 ( .B0(n2176), .B1(n2311), .A0N(\register[21][24] ), .A1N(
        n2313), .Y(n772) );
  OAI2BB2XL U1814 ( .B0(n2239), .B1(n2298), .A0N(\register[23][3] ), .A1N(
        n2301), .Y(n815) );
  OAI2BB2XL U1815 ( .B0(n2233), .B1(n2298), .A0N(\register[23][5] ), .A1N(
        n2301), .Y(n817) );
  OAI2BB2XL U1816 ( .B0(n2230), .B1(n2298), .A0N(\register[23][6] ), .A1N(
        n2301), .Y(n818) );
  OAI2BB2XL U1817 ( .B0(n2227), .B1(n2298), .A0N(\register[23][7] ), .A1N(
        n2301), .Y(n819) );
  OAI2BB2XL U1818 ( .B0(n2224), .B1(n2298), .A0N(\register[23][8] ), .A1N(
        n2301), .Y(n820) );
  OAI2BB2XL U1819 ( .B0(n2221), .B1(n2298), .A0N(\register[23][9] ), .A1N(
        n2301), .Y(n821) );
  OAI2BB2XL U1820 ( .B0(n2218), .B1(n2298), .A0N(\register[23][10] ), .A1N(
        n2301), .Y(n822) );
  OAI2BB2XL U1821 ( .B0(n2215), .B1(n2298), .A0N(\register[23][11] ), .A1N(
        n2301), .Y(n823) );
  OAI2BB2XL U1822 ( .B0(n2212), .B1(n2298), .A0N(\register[23][12] ), .A1N(
        n2301), .Y(n824) );
  OAI2BB2XL U1823 ( .B0(n2209), .B1(n2299), .A0N(\register[23][13] ), .A1N(
        n2301), .Y(n825) );
  OAI2BB2XL U1824 ( .B0(n2206), .B1(n2299), .A0N(\register[23][14] ), .A1N(
        n2301), .Y(n826) );
  OAI2BB2XL U1825 ( .B0(n2200), .B1(n2299), .A0N(\register[23][16] ), .A1N(
        n2301), .Y(n828) );
  OAI2BB2XL U1826 ( .B0(n2182), .B1(n2299), .A0N(\register[23][22] ), .A1N(
        n2301), .Y(n834) );
  OAI2BB2XL U1827 ( .B0(n2176), .B1(n2299), .A0N(\register[23][24] ), .A1N(
        n2301), .Y(n836) );
  OAI2BB2XL U1828 ( .B0(n2239), .B1(n2262), .A0N(\register[29][3] ), .A1N(
        n2265), .Y(n1007) );
  OAI2BB2XL U1829 ( .B0(n2233), .B1(n2262), .A0N(\register[29][5] ), .A1N(
        n2265), .Y(n1009) );
  OAI2BB2XL U1830 ( .B0(n2230), .B1(n2262), .A0N(\register[29][6] ), .A1N(
        n2265), .Y(n1010) );
  OAI2BB2XL U1831 ( .B0(n2227), .B1(n2262), .A0N(\register[29][7] ), .A1N(
        n2265), .Y(n1011) );
  OAI2BB2XL U1832 ( .B0(n2224), .B1(n2262), .A0N(\register[29][8] ), .A1N(
        n2265), .Y(n1012) );
  OAI2BB2XL U1833 ( .B0(n2221), .B1(n2262), .A0N(\register[29][9] ), .A1N(
        n2265), .Y(n1013) );
  OAI2BB2XL U1834 ( .B0(n2218), .B1(n2262), .A0N(\register[29][10] ), .A1N(
        n2265), .Y(n1014) );
  OAI2BB2XL U1835 ( .B0(n2215), .B1(n2263), .A0N(\register[29][11] ), .A1N(
        n2265), .Y(n1015) );
  OAI2BB2XL U1836 ( .B0(n2212), .B1(n2262), .A0N(\register[29][12] ), .A1N(
        n2265), .Y(n1016) );
  OAI2BB2XL U1837 ( .B0(n2209), .B1(n2263), .A0N(\register[29][13] ), .A1N(
        n2265), .Y(n1017) );
  OAI2BB2XL U1838 ( .B0(n2206), .B1(n2263), .A0N(\register[29][14] ), .A1N(
        n2265), .Y(n1018) );
  OAI2BB2XL U1839 ( .B0(n2200), .B1(n2263), .A0N(\register[29][16] ), .A1N(
        n2265), .Y(n1020) );
  OAI2BB2XL U1840 ( .B0(n2182), .B1(n2263), .A0N(\register[29][22] ), .A1N(
        n2265), .Y(n1026) );
  OAI2BB2XL U1841 ( .B0(n2176), .B1(n2263), .A0N(\register[29][24] ), .A1N(
        n2265), .Y(n1028) );
  OAI2BB2XL U1842 ( .B0(n2239), .B1(n2252), .A0N(\register[31][3] ), .A1N(
        n2255), .Y(n1071) );
  OAI2BB2XL U1843 ( .B0(n2233), .B1(n2252), .A0N(\register[31][5] ), .A1N(
        n2255), .Y(n1073) );
  OAI2BB2XL U1844 ( .B0(n2230), .B1(n2252), .A0N(\register[31][6] ), .A1N(
        n2255), .Y(n1074) );
  OAI2BB2XL U1845 ( .B0(n2227), .B1(n2252), .A0N(\register[31][7] ), .A1N(
        n2255), .Y(n1075) );
  OAI2BB2XL U1846 ( .B0(n2224), .B1(n2252), .A0N(\register[31][8] ), .A1N(
        n2255), .Y(n1076) );
  OAI2BB2XL U1847 ( .B0(n2221), .B1(n2252), .A0N(\register[31][9] ), .A1N(
        n2255), .Y(n1077) );
  OAI2BB2XL U1848 ( .B0(n2218), .B1(n2252), .A0N(\register[31][10] ), .A1N(
        n2255), .Y(n1078) );
  OAI2BB2XL U1849 ( .B0(n2215), .B1(n2252), .A0N(\register[31][11] ), .A1N(
        n2255), .Y(n1079) );
  OAI2BB2XL U1850 ( .B0(n2212), .B1(n2252), .A0N(\register[31][12] ), .A1N(
        n2255), .Y(n1080) );
  OAI2BB2XL U1851 ( .B0(n2209), .B1(n2253), .A0N(\register[31][13] ), .A1N(
        n2255), .Y(n1081) );
  OAI2BB2XL U1852 ( .B0(n2206), .B1(n2253), .A0N(\register[31][14] ), .A1N(
        n2255), .Y(n1082) );
  OAI2BB2XL U1853 ( .B0(n2200), .B1(n2253), .A0N(\register[31][16] ), .A1N(
        n2255), .Y(n1084) );
  OAI2BB2XL U1854 ( .B0(n2182), .B1(n2253), .A0N(\register[31][22] ), .A1N(
        n2255), .Y(n1090) );
  OAI2BB2XL U1855 ( .B0(n2176), .B1(n2253), .A0N(\register[31][24] ), .A1N(
        n2255), .Y(n1092) );
  OAI2BB2XL U1856 ( .B0(n2248), .B1(n2355), .A0N(\register[13][0] ), .A1N(
        n2352), .Y(n492) );
  OAI2BB2XL U1857 ( .B0(n2245), .B1(n2354), .A0N(\register[13][1] ), .A1N(
        n2352), .Y(n493) );
  OAI2BB2XL U1858 ( .B0(n2242), .B1(n2354), .A0N(\register[13][2] ), .A1N(
        n2352), .Y(n494) );
  OAI2BB2XL U1859 ( .B0(n2237), .B1(n2354), .A0N(\register[13][4] ), .A1N(
        n2352), .Y(n496) );
  OAI2BB2XL U1860 ( .B0(n2248), .B1(n2345), .A0N(\register[15][0] ), .A1N(
        n2342), .Y(n556) );
  OAI2BB2XL U1861 ( .B0(n2245), .B1(n2344), .A0N(\register[15][1] ), .A1N(
        n2342), .Y(n557) );
  OAI2BB2XL U1862 ( .B0(n2242), .B1(n2344), .A0N(\register[15][2] ), .A1N(
        n2342), .Y(n558) );
  OAI2BB2XL U1863 ( .B0(n2237), .B1(n2344), .A0N(\register[15][4] ), .A1N(
        n2342), .Y(n560) );
  OAI2BB2XL U1864 ( .B0(n2247), .B1(n2311), .A0N(\register[21][0] ), .A1N(
        n2308), .Y(n748) );
  OAI2BB2XL U1865 ( .B0(n2244), .B1(n2310), .A0N(\register[21][1] ), .A1N(
        n2308), .Y(n749) );
  OAI2BB2XL U1866 ( .B0(n2241), .B1(n2310), .A0N(\register[21][2] ), .A1N(
        n2308), .Y(n750) );
  OAI2BB2XL U1867 ( .B0(n2236), .B1(n2310), .A0N(\register[21][4] ), .A1N(
        n2308), .Y(n752) );
  OAI2BB2XL U1868 ( .B0(n2247), .B1(n2299), .A0N(\register[23][0] ), .A1N(
        n2296), .Y(n812) );
  OAI2BB2XL U1869 ( .B0(n2244), .B1(n2298), .A0N(\register[23][1] ), .A1N(
        n2296), .Y(n813) );
  OAI2BB2XL U1870 ( .B0(n2241), .B1(n2298), .A0N(\register[23][2] ), .A1N(
        n2296), .Y(n814) );
  OAI2BB2XL U1871 ( .B0(n2236), .B1(n2298), .A0N(\register[23][4] ), .A1N(
        n2296), .Y(n816) );
  OAI2BB2XL U1872 ( .B0(n2247), .B1(n2263), .A0N(\register[29][0] ), .A1N(
        n2262), .Y(n1004) );
  OAI2BB2XL U1873 ( .B0(n2244), .B1(n2263), .A0N(\register[29][1] ), .A1N(
        n2262), .Y(n1005) );
  OAI2BB2XL U1874 ( .B0(n2241), .B1(n2262), .A0N(\register[29][2] ), .A1N(
        n2262), .Y(n1006) );
  OAI2BB2XL U1875 ( .B0(n2236), .B1(n2263), .A0N(\register[29][4] ), .A1N(
        n2262), .Y(n1008) );
  OAI2BB2XL U1876 ( .B0(n2247), .B1(n2253), .A0N(\register[31][0] ), .A1N(
        n2250), .Y(n1068) );
  OAI2BB2XL U1877 ( .B0(n2244), .B1(n2252), .A0N(\register[31][1] ), .A1N(
        n2250), .Y(n1069) );
  OAI2BB2XL U1878 ( .B0(n2241), .B1(n2252), .A0N(\register[31][2] ), .A1N(
        n2250), .Y(n1070) );
  OAI2BB2XL U1879 ( .B0(n2236), .B1(n2252), .A0N(\register[31][4] ), .A1N(
        n2250), .Y(n1072) );
  OAI2BB2XL U1880 ( .B0(n2249), .B1(n2420), .A0N(\register[2][0] ), .A1N(n2417), .Y(n140) );
  OAI2BB2XL U1881 ( .B0(n2246), .B1(n2419), .A0N(\register[2][1] ), .A1N(n2417), .Y(n141) );
  OAI2BB2XL U1882 ( .B0(n2243), .B1(n2419), .A0N(\register[2][2] ), .A1N(n2417), .Y(n142) );
  OAI2BB2XL U1883 ( .B0(n2239), .B1(n2419), .A0N(\register[2][3] ), .A1N(n2422), .Y(n143) );
  OAI2BB2XL U1884 ( .B0(n2238), .B1(n2419), .A0N(\register[2][4] ), .A1N(n2417), .Y(n144) );
  OAI2BB2XL U1885 ( .B0(n2235), .B1(n2419), .A0N(\register[2][5] ), .A1N(n2422), .Y(n145) );
  OAI2BB2XL U1886 ( .B0(n2232), .B1(n2419), .A0N(\register[2][6] ), .A1N(n2422), .Y(n146) );
  OAI2BB2XL U1887 ( .B0(n2229), .B1(n2419), .A0N(\register[2][7] ), .A1N(n2422), .Y(n147) );
  OAI2BB2XL U1888 ( .B0(n2226), .B1(n2419), .A0N(\register[2][8] ), .A1N(n2422), .Y(n148) );
  OAI2BB2XL U1889 ( .B0(n2223), .B1(n2419), .A0N(\register[2][9] ), .A1N(n2422), .Y(n149) );
  OAI2BB2XL U1890 ( .B0(n2220), .B1(n2419), .A0N(\register[2][10] ), .A1N(
        n2422), .Y(n150) );
  OAI2BB2XL U1891 ( .B0(n2217), .B1(n2419), .A0N(\register[2][11] ), .A1N(
        n2422), .Y(n151) );
  OAI2BB2XL U1892 ( .B0(n2214), .B1(n2419), .A0N(\register[2][12] ), .A1N(
        n2422), .Y(n152) );
  OAI2BB2XL U1893 ( .B0(n2211), .B1(n2420), .A0N(\register[2][13] ), .A1N(
        n2422), .Y(n153) );
  OAI2BB2XL U1894 ( .B0(n2208), .B1(n2420), .A0N(\register[2][14] ), .A1N(
        n2422), .Y(n154) );
  OAI2BB2XL U1895 ( .B0(n2205), .B1(n2420), .A0N(\register[2][15] ), .A1N(
        n2421), .Y(n155) );
  OAI2BB2XL U1896 ( .B0(n2202), .B1(n2420), .A0N(\register[2][16] ), .A1N(
        n2422), .Y(n156) );
  OAI2BB2XL U1897 ( .B0(n2199), .B1(n2420), .A0N(\register[2][17] ), .A1N(
        n2421), .Y(n157) );
  OAI2BB2XL U1898 ( .B0(n2196), .B1(n2420), .A0N(\register[2][18] ), .A1N(
        n2421), .Y(n158) );
  OAI2BB2XL U1899 ( .B0(n2193), .B1(n2420), .A0N(\register[2][19] ), .A1N(
        n2421), .Y(n159) );
  OAI2BB2XL U1900 ( .B0(n2190), .B1(n2420), .A0N(\register[2][20] ), .A1N(
        n2421), .Y(n160) );
  OAI2BB2XL U1901 ( .B0(n2187), .B1(n2420), .A0N(\register[2][21] ), .A1N(
        n2421), .Y(n161) );
  OAI2BB2XL U1902 ( .B0(n2184), .B1(n2420), .A0N(\register[2][22] ), .A1N(
        n2422), .Y(n162) );
  OAI2BB2XL U1903 ( .B0(n2178), .B1(n2420), .A0N(\register[2][24] ), .A1N(
        n2422), .Y(n164) );
  OAI2BB2XL U1904 ( .B0(n2249), .B1(n2413), .A0N(\register[3][0] ), .A1N(n2416), .Y(n172) );
  OAI2BB2XL U1905 ( .B0(n2246), .B1(n2412), .A0N(\register[3][1] ), .A1N(n2416), .Y(n173) );
  OAI2BB2XL U1906 ( .B0(n2243), .B1(n2412), .A0N(\register[3][2] ), .A1N(n2416), .Y(n174) );
  OAI2BB2XL U1907 ( .B0(n2239), .B1(n2412), .A0N(\register[3][3] ), .A1N(n2415), .Y(n175) );
  OAI2BB2XL U1908 ( .B0(n2238), .B1(n2412), .A0N(\register[3][4] ), .A1N(n2416), .Y(n176) );
  OAI2BB2XL U1909 ( .B0(n2235), .B1(n2412), .A0N(\register[3][5] ), .A1N(n2415), .Y(n177) );
  OAI2BB2XL U1910 ( .B0(n2232), .B1(n2412), .A0N(\register[3][6] ), .A1N(n2415), .Y(n178) );
  OAI2BB2XL U1911 ( .B0(n2229), .B1(n2412), .A0N(\register[3][7] ), .A1N(n2415), .Y(n179) );
  OAI2BB2XL U1912 ( .B0(n2226), .B1(n2412), .A0N(\register[3][8] ), .A1N(n2415), .Y(n180) );
  OAI2BB2XL U1913 ( .B0(n2223), .B1(n2412), .A0N(\register[3][9] ), .A1N(n2415), .Y(n181) );
  OAI2BB2XL U1914 ( .B0(n2220), .B1(n2412), .A0N(\register[3][10] ), .A1N(
        n2415), .Y(n182) );
  OAI2BB2XL U1915 ( .B0(n2217), .B1(n2412), .A0N(\register[3][11] ), .A1N(
        n2415), .Y(n183) );
  OAI2BB2XL U1916 ( .B0(n2214), .B1(n2412), .A0N(\register[3][12] ), .A1N(
        n2415), .Y(n184) );
  OAI2BB2XL U1917 ( .B0(n2211), .B1(n2413), .A0N(\register[3][13] ), .A1N(
        n2415), .Y(n185) );
  OAI2BB2XL U1918 ( .B0(n2208), .B1(n2413), .A0N(\register[3][14] ), .A1N(
        n2415), .Y(n186) );
  OAI2BB2XL U1919 ( .B0(n2205), .B1(n2413), .A0N(\register[3][15] ), .A1N(
        n2414), .Y(n187) );
  OAI2BB2XL U1920 ( .B0(n2202), .B1(n2413), .A0N(\register[3][16] ), .A1N(
        n2415), .Y(n188) );
  OAI2BB2XL U1921 ( .B0(n2199), .B1(n2413), .A0N(\register[3][17] ), .A1N(
        n2414), .Y(n189) );
  OAI2BB2XL U1922 ( .B0(n2196), .B1(n2413), .A0N(\register[3][18] ), .A1N(
        n2414), .Y(n190) );
  OAI2BB2XL U1923 ( .B0(n2193), .B1(n2413), .A0N(\register[3][19] ), .A1N(
        n2414), .Y(n191) );
  OAI2BB2XL U1924 ( .B0(n2190), .B1(n2413), .A0N(\register[3][20] ), .A1N(
        n2414), .Y(n192) );
  OAI2BB2XL U1925 ( .B0(n2187), .B1(n2413), .A0N(\register[3][21] ), .A1N(
        n2414), .Y(n193) );
  OAI2BB2XL U1926 ( .B0(n2184), .B1(n2413), .A0N(\register[3][22] ), .A1N(
        n2415), .Y(n194) );
  OAI2BB2XL U1927 ( .B0(n2178), .B1(n2413), .A0N(\register[3][24] ), .A1N(
        n2415), .Y(n196) );
  OAI2BB2XL U1928 ( .B0(n2249), .B1(n2426), .A0N(\register[1][0] ), .A1N(n2423), .Y(n108) );
  OAI2BB2XL U1929 ( .B0(n2246), .B1(n2425), .A0N(\register[1][1] ), .A1N(n2423), .Y(n109) );
  OAI2BB2XL U1930 ( .B0(n2243), .B1(n2425), .A0N(\register[1][2] ), .A1N(n2423), .Y(n110) );
  OAI2BB2XL U1931 ( .B0(n2239), .B1(n2425), .A0N(\register[1][3] ), .A1N(n2428), .Y(n111) );
  OAI2BB2XL U1932 ( .B0(n2238), .B1(n2425), .A0N(\register[1][4] ), .A1N(n2423), .Y(n112) );
  OAI2BB2XL U1933 ( .B0(n2235), .B1(n2425), .A0N(\register[1][5] ), .A1N(n2428), .Y(n113) );
  OAI2BB2XL U1934 ( .B0(n2232), .B1(n2425), .A0N(\register[1][6] ), .A1N(n2428), .Y(n114) );
  OAI2BB2XL U1935 ( .B0(n2229), .B1(n2425), .A0N(\register[1][7] ), .A1N(n2428), .Y(n115) );
  OAI2BB2XL U1936 ( .B0(n2226), .B1(n2425), .A0N(\register[1][8] ), .A1N(n2428), .Y(n116) );
  OAI2BB2XL U1937 ( .B0(n2223), .B1(n2425), .A0N(\register[1][9] ), .A1N(n2428), .Y(n117) );
  OAI2BB2XL U1938 ( .B0(n2220), .B1(n2425), .A0N(\register[1][10] ), .A1N(
        n2428), .Y(n118) );
  OAI2BB2XL U1939 ( .B0(n2217), .B1(n2425), .A0N(\register[1][11] ), .A1N(
        n2428), .Y(n119) );
  OAI2BB2XL U1940 ( .B0(n2214), .B1(n2425), .A0N(\register[1][12] ), .A1N(
        n2428), .Y(n120) );
  OAI2BB2XL U1941 ( .B0(n2211), .B1(n2426), .A0N(\register[1][13] ), .A1N(
        n2428), .Y(n121) );
  OAI2BB2XL U1942 ( .B0(n2208), .B1(n2426), .A0N(\register[1][14] ), .A1N(
        n2428), .Y(n122) );
  OAI2BB2XL U1943 ( .B0(n2205), .B1(n2426), .A0N(\register[1][15] ), .A1N(
        n2427), .Y(n123) );
  OAI2BB2XL U1944 ( .B0(n2202), .B1(n2426), .A0N(\register[1][16] ), .A1N(
        n2428), .Y(n124) );
  OAI2BB2XL U1945 ( .B0(n2199), .B1(n2426), .A0N(\register[1][17] ), .A1N(
        n2427), .Y(n125) );
  OAI2BB2XL U1946 ( .B0(n2196), .B1(n2426), .A0N(\register[1][18] ), .A1N(
        n2427), .Y(n126) );
  OAI2BB2XL U1947 ( .B0(n2193), .B1(n2426), .A0N(\register[1][19] ), .A1N(
        n2427), .Y(n127) );
  OAI2BB2XL U1948 ( .B0(n2190), .B1(n2426), .A0N(\register[1][20] ), .A1N(
        n2427), .Y(n128) );
  OAI2BB2XL U1949 ( .B0(n2187), .B1(n2426), .A0N(\register[1][21] ), .A1N(
        n2427), .Y(n129) );
  OAI2BB2XL U1950 ( .B0(n2184), .B1(n2426), .A0N(\register[1][22] ), .A1N(
        n2428), .Y(n130) );
  OAI2BB2XL U1951 ( .B0(n2178), .B1(n2426), .A0N(\register[1][24] ), .A1N(
        n2428), .Y(n132) );
  OAI2BB2XL U1952 ( .B0(n2205), .B1(n2406), .A0N(\register[4][15] ), .A1N(
        n2407), .Y(n219) );
  OAI2BB2XL U1953 ( .B0(n2199), .B1(n2406), .A0N(\register[4][17] ), .A1N(
        n2407), .Y(n221) );
  OAI2BB2XL U1954 ( .B0(n2196), .B1(n2406), .A0N(\register[4][18] ), .A1N(
        n2407), .Y(n222) );
  OAI2BB2XL U1955 ( .B0(n2193), .B1(n2406), .A0N(\register[4][19] ), .A1N(
        n2407), .Y(n223) );
  OAI2BB2XL U1956 ( .B0(n2190), .B1(n2406), .A0N(\register[4][20] ), .A1N(
        n2407), .Y(n224) );
  OAI2BB2XL U1957 ( .B0(n2187), .B1(n2406), .A0N(\register[4][21] ), .A1N(
        n2407), .Y(n225) );
  OAI2BB2XL U1958 ( .B0(n2205), .B1(n2394), .A0N(\register[6][15] ), .A1N(
        n2395), .Y(n283) );
  OAI2BB2XL U1959 ( .B0(n2199), .B1(n2394), .A0N(\register[6][17] ), .A1N(
        n2395), .Y(n285) );
  OAI2BB2XL U1960 ( .B0(n2196), .B1(n2394), .A0N(\register[6][18] ), .A1N(
        n2395), .Y(n286) );
  OAI2BB2XL U1961 ( .B0(n2193), .B1(n2394), .A0N(\register[6][19] ), .A1N(
        n2395), .Y(n287) );
  OAI2BB2XL U1962 ( .B0(n2190), .B1(n2394), .A0N(\register[6][20] ), .A1N(
        n2395), .Y(n288) );
  OAI2BB2XL U1963 ( .B0(n2187), .B1(n2394), .A0N(\register[6][21] ), .A1N(
        n2395), .Y(n289) );
  OAI2BB2XL U1964 ( .B0(n2239), .B1(n2405), .A0N(\register[4][3] ), .A1N(n2408), .Y(n207) );
  OAI2BB2XL U1965 ( .B0(n2235), .B1(n2405), .A0N(\register[4][5] ), .A1N(n2408), .Y(n209) );
  OAI2BB2XL U1966 ( .B0(n2232), .B1(n2405), .A0N(\register[4][6] ), .A1N(n2408), .Y(n210) );
  OAI2BB2XL U1967 ( .B0(n2229), .B1(n2405), .A0N(\register[4][7] ), .A1N(n2408), .Y(n211) );
  OAI2BB2XL U1968 ( .B0(n2226), .B1(n2405), .A0N(\register[4][8] ), .A1N(n2408), .Y(n212) );
  OAI2BB2XL U1969 ( .B0(n2223), .B1(n2405), .A0N(\register[4][9] ), .A1N(n2408), .Y(n213) );
  OAI2BB2XL U1970 ( .B0(n2220), .B1(n2405), .A0N(\register[4][10] ), .A1N(
        n2408), .Y(n214) );
  OAI2BB2XL U1971 ( .B0(n2217), .B1(n2405), .A0N(\register[4][11] ), .A1N(
        n2408), .Y(n215) );
  OAI2BB2XL U1972 ( .B0(n2214), .B1(n2405), .A0N(\register[4][12] ), .A1N(
        n2408), .Y(n216) );
  OAI2BB2XL U1973 ( .B0(n2211), .B1(n2406), .A0N(\register[4][13] ), .A1N(
        n2408), .Y(n217) );
  OAI2BB2XL U1974 ( .B0(n2208), .B1(n2406), .A0N(\register[4][14] ), .A1N(
        n2408), .Y(n218) );
  OAI2BB2XL U1975 ( .B0(n2202), .B1(n2406), .A0N(\register[4][16] ), .A1N(
        n2408), .Y(n220) );
  OAI2BB2XL U1976 ( .B0(n2184), .B1(n2406), .A0N(\register[4][22] ), .A1N(
        n2408), .Y(n226) );
  OAI2BB2XL U1977 ( .B0(n2178), .B1(n2406), .A0N(\register[4][24] ), .A1N(
        n2408), .Y(n228) );
  OAI2BB2XL U1978 ( .B0(n2239), .B1(n2393), .A0N(\register[6][3] ), .A1N(n2396), .Y(n271) );
  OAI2BB2XL U1979 ( .B0(n2235), .B1(n2393), .A0N(\register[6][5] ), .A1N(n2396), .Y(n273) );
  OAI2BB2XL U1980 ( .B0(n2232), .B1(n2393), .A0N(\register[6][6] ), .A1N(n2396), .Y(n274) );
  OAI2BB2XL U1981 ( .B0(n2229), .B1(n2393), .A0N(\register[6][7] ), .A1N(n2396), .Y(n275) );
  OAI2BB2XL U1982 ( .B0(n2226), .B1(n2393), .A0N(\register[6][8] ), .A1N(n2396), .Y(n276) );
  OAI2BB2XL U1983 ( .B0(n2223), .B1(n2393), .A0N(\register[6][9] ), .A1N(n2396), .Y(n277) );
  OAI2BB2XL U1984 ( .B0(n2220), .B1(n2393), .A0N(\register[6][10] ), .A1N(
        n2396), .Y(n278) );
  OAI2BB2XL U1985 ( .B0(n2217), .B1(n2393), .A0N(\register[6][11] ), .A1N(
        n2396), .Y(n279) );
  OAI2BB2XL U1986 ( .B0(n2214), .B1(n2393), .A0N(\register[6][12] ), .A1N(
        n2396), .Y(n280) );
  OAI2BB2XL U1987 ( .B0(n2211), .B1(n2394), .A0N(\register[6][13] ), .A1N(
        n2396), .Y(n281) );
  OAI2BB2XL U1988 ( .B0(n2208), .B1(n2394), .A0N(\register[6][14] ), .A1N(
        n2396), .Y(n282) );
  OAI2BB2XL U1989 ( .B0(n2202), .B1(n2394), .A0N(\register[6][16] ), .A1N(
        n2396), .Y(n284) );
  OAI2BB2XL U1990 ( .B0(n2184), .B1(n2394), .A0N(\register[6][22] ), .A1N(
        n2396), .Y(n290) );
  OAI2BB2XL U1991 ( .B0(n2178), .B1(n2394), .A0N(\register[6][24] ), .A1N(
        n2396), .Y(n292) );
  OAI2BB2XL U1992 ( .B0(n2249), .B1(n2406), .A0N(\register[4][0] ), .A1N(n2403), .Y(n204) );
  OAI2BB2XL U1993 ( .B0(n2246), .B1(n2405), .A0N(\register[4][1] ), .A1N(n2403), .Y(n205) );
  OAI2BB2XL U1994 ( .B0(n2243), .B1(n2405), .A0N(\register[4][2] ), .A1N(n2403), .Y(n206) );
  OAI2BB2XL U1995 ( .B0(n2238), .B1(n2405), .A0N(\register[4][4] ), .A1N(n2403), .Y(n208) );
  OAI2BB2XL U1996 ( .B0(n2249), .B1(n2394), .A0N(\register[6][0] ), .A1N(n2394), .Y(n268) );
  OAI2BB2XL U1997 ( .B0(n2246), .B1(n2393), .A0N(\register[6][1] ), .A1N(n2393), .Y(n269) );
  OAI2BB2XL U1998 ( .B0(n2243), .B1(n2393), .A0N(\register[6][2] ), .A1N(n2394), .Y(n270) );
  OAI2BB2XL U1999 ( .B0(n2238), .B1(n2393), .A0N(\register[6][4] ), .A1N(n2393), .Y(n272) );
  OAI2BB2XL U2000 ( .B0(n2205), .B1(n2400), .A0N(\register[5][15] ), .A1N(
        n2401), .Y(n251) );
  OAI2BB2XL U2001 ( .B0(n2199), .B1(n2400), .A0N(\register[5][17] ), .A1N(
        n2401), .Y(n253) );
  OAI2BB2XL U2002 ( .B0(n2196), .B1(n2400), .A0N(\register[5][18] ), .A1N(
        n2401), .Y(n254) );
  OAI2BB2XL U2003 ( .B0(n2193), .B1(n2400), .A0N(\register[5][19] ), .A1N(
        n2401), .Y(n255) );
  OAI2BB2XL U2004 ( .B0(n2190), .B1(n2400), .A0N(\register[5][20] ), .A1N(
        n2401), .Y(n256) );
  OAI2BB2XL U2005 ( .B0(n2187), .B1(n2400), .A0N(\register[5][21] ), .A1N(
        n2401), .Y(n257) );
  OAI2BB2XL U2006 ( .B0(n2205), .B1(n2391), .A0N(\register[7][15] ), .A1N(
        n2391), .Y(n315) );
  OAI2BB2XL U2007 ( .B0(n2199), .B1(n2391), .A0N(\register[7][17] ), .A1N(
        n2388), .Y(n317) );
  OAI2BB2XL U2008 ( .B0(n2196), .B1(n2391), .A0N(\register[7][18] ), .A1N(
        n2391), .Y(n318) );
  OAI2BB2XL U2009 ( .B0(n2193), .B1(n2391), .A0N(\register[7][19] ), .A1N(
        n2390), .Y(n319) );
  OAI2BB2XL U2010 ( .B0(n2190), .B1(n2391), .A0N(\register[7][20] ), .A1N(
        n2388), .Y(n320) );
  OAI2BB2XL U2011 ( .B0(n2187), .B1(n2391), .A0N(\register[7][21] ), .A1N(
        n2391), .Y(n321) );
  OAI2BB2XL U2012 ( .B0(n2239), .B1(n2399), .A0N(\register[5][3] ), .A1N(n2402), .Y(n239) );
  OAI2BB2XL U2013 ( .B0(n2235), .B1(n2399), .A0N(\register[5][5] ), .A1N(n2402), .Y(n241) );
  OAI2BB2XL U2014 ( .B0(n2232), .B1(n2399), .A0N(\register[5][6] ), .A1N(n2402), .Y(n242) );
  OAI2BB2XL U2015 ( .B0(n2229), .B1(n2399), .A0N(\register[5][7] ), .A1N(n2402), .Y(n243) );
  OAI2BB2XL U2016 ( .B0(n2226), .B1(n2399), .A0N(\register[5][8] ), .A1N(n2402), .Y(n244) );
  OAI2BB2XL U2017 ( .B0(n2223), .B1(n2399), .A0N(\register[5][9] ), .A1N(n2402), .Y(n245) );
  OAI2BB2XL U2018 ( .B0(n2220), .B1(n2399), .A0N(\register[5][10] ), .A1N(
        n2402), .Y(n246) );
  OAI2BB2XL U2019 ( .B0(n2217), .B1(n2399), .A0N(\register[5][11] ), .A1N(
        n2402), .Y(n247) );
  OAI2BB2XL U2020 ( .B0(n2214), .B1(n2399), .A0N(\register[5][12] ), .A1N(
        n2402), .Y(n248) );
  OAI2BB2XL U2021 ( .B0(n2211), .B1(n2400), .A0N(\register[5][13] ), .A1N(
        n2402), .Y(n249) );
  OAI2BB2XL U2022 ( .B0(n2208), .B1(n2400), .A0N(\register[5][14] ), .A1N(
        n2402), .Y(n250) );
  OAI2BB2XL U2023 ( .B0(n2202), .B1(n2400), .A0N(\register[5][16] ), .A1N(
        n2402), .Y(n252) );
  OAI2BB2XL U2024 ( .B0(n2184), .B1(n2400), .A0N(\register[5][22] ), .A1N(
        n2402), .Y(n258) );
  OAI2BB2XL U2025 ( .B0(n2178), .B1(n2400), .A0N(\register[5][24] ), .A1N(
        n2402), .Y(n260) );
  OAI2BB2XL U2026 ( .B0(n2239), .B1(n2390), .A0N(\register[7][3] ), .A1N(n2392), .Y(n303) );
  OAI2BB2XL U2027 ( .B0(n2235), .B1(n2390), .A0N(\register[7][5] ), .A1N(n2392), .Y(n305) );
  OAI2BB2XL U2028 ( .B0(n2232), .B1(n2390), .A0N(\register[7][6] ), .A1N(n2392), .Y(n306) );
  OAI2BB2XL U2029 ( .B0(n2229), .B1(n2390), .A0N(\register[7][7] ), .A1N(n2392), .Y(n307) );
  OAI2BB2XL U2030 ( .B0(n2226), .B1(n2390), .A0N(\register[7][8] ), .A1N(n2392), .Y(n308) );
  OAI2BB2XL U2031 ( .B0(n2223), .B1(n2390), .A0N(\register[7][9] ), .A1N(n2392), .Y(n309) );
  OAI2BB2XL U2032 ( .B0(n2220), .B1(n2390), .A0N(\register[7][10] ), .A1N(
        n2392), .Y(n310) );
  OAI2BB2XL U2033 ( .B0(n2217), .B1(n2390), .A0N(\register[7][11] ), .A1N(
        n2392), .Y(n311) );
  OAI2BB2XL U2034 ( .B0(n2214), .B1(n2390), .A0N(\register[7][12] ), .A1N(
        n2392), .Y(n312) );
  OAI2BB2XL U2035 ( .B0(n2211), .B1(n2391), .A0N(\register[7][13] ), .A1N(
        n2392), .Y(n313) );
  OAI2BB2XL U2036 ( .B0(n2208), .B1(n2391), .A0N(\register[7][14] ), .A1N(
        n2392), .Y(n314) );
  OAI2BB2XL U2037 ( .B0(n2202), .B1(n2391), .A0N(\register[7][16] ), .A1N(
        n2392), .Y(n316) );
  OAI2BB2XL U2038 ( .B0(n2184), .B1(n2391), .A0N(\register[7][22] ), .A1N(
        n2392), .Y(n322) );
  OAI2BB2XL U2039 ( .B0(n2178), .B1(n2391), .A0N(\register[7][24] ), .A1N(
        n2392), .Y(n324) );
  OAI2BB2XL U2040 ( .B0(n2249), .B1(n2400), .A0N(\register[5][0] ), .A1N(n2397), .Y(n236) );
  OAI2BB2XL U2041 ( .B0(n2246), .B1(n2399), .A0N(\register[5][1] ), .A1N(n2397), .Y(n237) );
  OAI2BB2XL U2042 ( .B0(n2243), .B1(n2399), .A0N(\register[5][2] ), .A1N(n2397), .Y(n238) );
  OAI2BB2XL U2043 ( .B0(n2238), .B1(n2399), .A0N(\register[5][4] ), .A1N(n2397), .Y(n240) );
  OAI2BB2XL U2044 ( .B0(n2249), .B1(n2391), .A0N(\register[7][0] ), .A1N(n2388), .Y(n300) );
  OAI2BB2XL U2045 ( .B0(n2246), .B1(n2390), .A0N(\register[7][1] ), .A1N(n2388), .Y(n301) );
  OAI2BB2XL U2046 ( .B0(n2243), .B1(n2390), .A0N(\register[7][2] ), .A1N(n2388), .Y(n302) );
  OAI2BB2XL U2047 ( .B0(n2238), .B1(n2390), .A0N(\register[7][4] ), .A1N(n2388), .Y(n304) );
  NOR2BX1 U2048 ( .AN(n2128), .B(\register[3][0] ), .Y(n2085) );
  NOR2BX1 U2049 ( .AN(n2128), .B(\register[3][1] ), .Y(n2080) );
  NOR2BX1 U2050 ( .AN(n2128), .B(\register[3][2] ), .Y(n2075) );
  NOR2BX1 U2051 ( .AN(n2128), .B(\register[3][3] ), .Y(n2070) );
  NOR2BX1 U2052 ( .AN(n2128), .B(\register[3][4] ), .Y(n2065) );
  NOR2BX1 U2053 ( .AN(n2127), .B(\register[3][5] ), .Y(n2060) );
  NOR2BX1 U2054 ( .AN(n2128), .B(\register[3][6] ), .Y(n2055) );
  NOR2BX1 U2055 ( .AN(n2127), .B(\register[3][8] ), .Y(n2045) );
  NOR2BX1 U2056 ( .AN(n2127), .B(\register[3][9] ), .Y(n2040) );
  NOR2BX1 U2057 ( .AN(n2127), .B(\register[3][10] ), .Y(n2035) );
  NOR2BX1 U2058 ( .AN(n2127), .B(\register[3][11] ), .Y(n2030) );
  NOR2BX1 U2059 ( .AN(n2128), .B(\register[3][12] ), .Y(n2025) );
  NOR2BX1 U2060 ( .AN(n2127), .B(\register[3][13] ), .Y(n2020) );
  NOR2BX1 U2061 ( .AN(n2127), .B(\register[3][14] ), .Y(n2015) );
  NOR2BX1 U2062 ( .AN(n2127), .B(\register[3][15] ), .Y(n2010) );
  NOR2BX1 U2063 ( .AN(n2127), .B(\register[3][16] ), .Y(n2005) );
  NOR2BX1 U2064 ( .AN(n2127), .B(\register[3][17] ), .Y(n2000) );
  NOR2BX1 U2065 ( .AN(n2127), .B(\register[3][18] ), .Y(n1995) );
  NOR2BX1 U2066 ( .AN(n2127), .B(\register[3][19] ), .Y(n1990) );
  NOR2BX1 U2067 ( .AN(n2127), .B(\register[3][21] ), .Y(n1980) );
  NOR2BX1 U2068 ( .AN(n2127), .B(\register[3][22] ), .Y(n1975) );
  NOR2BX1 U2069 ( .AN(n2127), .B(\register[3][23] ), .Y(n1970) );
  NOR2BX1 U2070 ( .AN(n2127), .B(\register[3][24] ), .Y(n1965) );
  NOR2BX1 U2071 ( .AN(n2128), .B(\register[3][25] ), .Y(n1960) );
  NOR2BX1 U2072 ( .AN(n2128), .B(\register[3][26] ), .Y(n1955) );
  NOR2BX1 U2073 ( .AN(n2128), .B(\register[3][27] ), .Y(n1950) );
  NOR2BX1 U2074 ( .AN(n2128), .B(\register[3][28] ), .Y(n1945) );
  NOR2BX1 U2075 ( .AN(n2128), .B(\register[3][29] ), .Y(n1940) );
  NOR2BX1 U2076 ( .AN(n2128), .B(\register[3][30] ), .Y(n1935) );
  NOR2BX1 U2077 ( .AN(n2128), .B(\register[3][31] ), .Y(n1930) );
  NOR2BX1 U2078 ( .AN(n1584), .B(\register[3][0] ), .Y(n1541) );
  NOR2BX1 U2079 ( .AN(n1584), .B(\register[3][2] ), .Y(n1531) );
  NOR2BX1 U2080 ( .AN(n1584), .B(\register[3][3] ), .Y(n1526) );
  NOR2BX1 U2081 ( .AN(n1584), .B(\register[3][4] ), .Y(n1521) );
  NOR2BX1 U2082 ( .AN(n1583), .B(\register[3][5] ), .Y(n1516) );
  NOR2BX1 U2083 ( .AN(n1584), .B(\register[3][6] ), .Y(n1511) );
  NOR2BX1 U2084 ( .AN(n1583), .B(\register[3][7] ), .Y(n1506) );
  NOR2BX1 U2085 ( .AN(n1583), .B(\register[3][8] ), .Y(n1501) );
  NOR2BX1 U2086 ( .AN(n1583), .B(\register[3][9] ), .Y(n1496) );
  NOR2BX1 U2087 ( .AN(n1583), .B(\register[3][10] ), .Y(n1491) );
  NOR2BX1 U2088 ( .AN(n1583), .B(\register[3][11] ), .Y(n1486) );
  NOR2BX1 U2089 ( .AN(n1584), .B(\register[3][12] ), .Y(n1481) );
  NOR2BX1 U2090 ( .AN(n1583), .B(\register[3][13] ), .Y(n1476) );
  NOR2BX1 U2091 ( .AN(n1583), .B(\register[3][15] ), .Y(n1466) );
  NOR2BX1 U2092 ( .AN(n1583), .B(\register[3][16] ), .Y(n1461) );
  NOR2BX1 U2093 ( .AN(n1583), .B(\register[3][17] ), .Y(n1456) );
  NOR2BX1 U2094 ( .AN(n1583), .B(\register[3][18] ), .Y(n1451) );
  NOR2BX1 U2095 ( .AN(n1583), .B(\register[3][19] ), .Y(n1446) );
  NOR2BX1 U2096 ( .AN(n1583), .B(\register[3][20] ), .Y(n1441) );
  NOR2BX1 U2097 ( .AN(n1583), .B(\register[3][21] ), .Y(n1436) );
  NOR2BX1 U2098 ( .AN(n1583), .B(\register[3][22] ), .Y(n1431) );
  NOR2BX1 U2099 ( .AN(n1583), .B(\register[3][23] ), .Y(n1426) );
  NOR2BX1 U2100 ( .AN(n1583), .B(\register[3][24] ), .Y(n1421) );
  NOR2BX1 U2101 ( .AN(n1584), .B(\register[3][25] ), .Y(n1416) );
  NOR2BX1 U2102 ( .AN(n1584), .B(\register[3][26] ), .Y(n1411) );
  NOR2BX1 U2103 ( .AN(n1584), .B(\register[3][27] ), .Y(n1406) );
  NOR2BX1 U2104 ( .AN(n1584), .B(\register[3][28] ), .Y(n1401) );
  NOR2BX1 U2105 ( .AN(n1584), .B(\register[3][29] ), .Y(n1396) );
  NOR2BX1 U2106 ( .AN(n1584), .B(\register[3][30] ), .Y(n1391) );
  NOR2BX1 U2107 ( .AN(n1584), .B(\register[3][31] ), .Y(n1386) );
  NOR2X1 U2108 ( .A(n1579), .B(\register[1][26] ), .Y(n1413) );
  NAND2X1 U2109 ( .A(n2084), .B(n2083), .Y(n1689) );
  NOR2X1 U2110 ( .A(n2082), .B(n2081), .Y(n2084) );
  MXI2X1 U2111 ( .A(n2555), .B(n2080), .S0(n2151), .Y(n2083) );
  NOR2X1 U2112 ( .A(n2130), .B(\register[1][1] ), .Y(n2082) );
  NAND2X1 U2113 ( .A(n1540), .B(n1539), .Y(n1145) );
  NOR2X1 U2114 ( .A(n1538), .B(n1537), .Y(n1540) );
  NOR2X1 U2115 ( .A(n1586), .B(\register[1][1] ), .Y(n1538) );
  NAND2X1 U2116 ( .A(n2079), .B(n2078), .Y(n1697) );
  NOR2X1 U2117 ( .A(n2077), .B(n2076), .Y(n2079) );
  MXI2X1 U2118 ( .A(n2556), .B(n2075), .S0(n2152), .Y(n2078) );
  NOR2X1 U2119 ( .A(n2130), .B(\register[1][2] ), .Y(n2077) );
  NAND2X1 U2120 ( .A(n2074), .B(n2073), .Y(n1705) );
  NOR2X1 U2121 ( .A(n2072), .B(n2071), .Y(n2074) );
  MXI2X1 U2122 ( .A(n2557), .B(n2070), .S0(n2152), .Y(n2073) );
  NOR2X1 U2123 ( .A(n2129), .B(\register[1][3] ), .Y(n2072) );
  NAND2X1 U2124 ( .A(n2069), .B(n2068), .Y(n1713) );
  NOR2X1 U2125 ( .A(n2067), .B(n2066), .Y(n2069) );
  MXI2X1 U2126 ( .A(n2558), .B(n2065), .S0(n2152), .Y(n2068) );
  NOR2X1 U2127 ( .A(n2128), .B(\register[1][4] ), .Y(n2067) );
  NAND2X1 U2128 ( .A(n2064), .B(n2063), .Y(n1721) );
  NOR2X1 U2129 ( .A(n2062), .B(n2061), .Y(n2064) );
  MXI2X1 U2130 ( .A(n2559), .B(n2060), .S0(n2152), .Y(n2063) );
  NOR2X1 U2131 ( .A(n2129), .B(\register[1][5] ), .Y(n2062) );
  NAND2X1 U2132 ( .A(n2059), .B(n2058), .Y(n1729) );
  NOR2X1 U2133 ( .A(n2057), .B(n2056), .Y(n2059) );
  MXI2X1 U2134 ( .A(n2560), .B(n2055), .S0(n2152), .Y(n2058) );
  NOR2X1 U2135 ( .A(n2128), .B(\register[1][6] ), .Y(n2057) );
  NAND2X1 U2136 ( .A(n2054), .B(n2053), .Y(n1737) );
  NOR2X1 U2137 ( .A(n2052), .B(n2051), .Y(n2054) );
  NOR2X1 U2138 ( .A(n2129), .B(\register[1][7] ), .Y(n2052) );
  NAND2X1 U2139 ( .A(n2049), .B(n2048), .Y(n1745) );
  NOR2X1 U2140 ( .A(n2047), .B(n2046), .Y(n2049) );
  MXI2X1 U2141 ( .A(n2562), .B(n2045), .S0(n2152), .Y(n2048) );
  NOR2X1 U2142 ( .A(n2130), .B(\register[1][8] ), .Y(n2047) );
  NAND2X1 U2143 ( .A(n2044), .B(n2043), .Y(n1753) );
  NOR2X1 U2144 ( .A(n2042), .B(n2041), .Y(n2044) );
  MXI2X1 U2145 ( .A(n2563), .B(n2040), .S0(n2152), .Y(n2043) );
  NOR2X1 U2146 ( .A(n2129), .B(\register[1][9] ), .Y(n2042) );
  NAND2X1 U2147 ( .A(n2039), .B(n2038), .Y(n1761) );
  NOR2X1 U2148 ( .A(n2037), .B(n2036), .Y(n2039) );
  MXI2X1 U2149 ( .A(n2564), .B(n2035), .S0(n2152), .Y(n2038) );
  NOR2X1 U2150 ( .A(n2129), .B(\register[1][10] ), .Y(n2037) );
  NAND2X1 U2151 ( .A(n2034), .B(n2033), .Y(n1769) );
  NOR2X1 U2152 ( .A(n2032), .B(n2031), .Y(n2034) );
  MXI2X1 U2153 ( .A(n2565), .B(n2030), .S0(n2152), .Y(n2033) );
  NOR2X1 U2154 ( .A(n2130), .B(\register[1][11] ), .Y(n2032) );
  NAND2X1 U2155 ( .A(n2029), .B(n2028), .Y(n1777) );
  NOR2X1 U2156 ( .A(n2027), .B(n2026), .Y(n2029) );
  MXI2X1 U2157 ( .A(n2566), .B(n2025), .S0(n2152), .Y(n2028) );
  NOR2X1 U2158 ( .A(n2130), .B(\register[1][12] ), .Y(n2027) );
  NAND2X1 U2159 ( .A(n2024), .B(n2023), .Y(n1785) );
  NOR2X1 U2160 ( .A(n2022), .B(n2021), .Y(n2024) );
  MXI2X1 U2161 ( .A(n2567), .B(n2020), .S0(n2152), .Y(n2023) );
  NOR2X1 U2162 ( .A(n2130), .B(\register[1][13] ), .Y(n2022) );
  NAND2X1 U2163 ( .A(n2019), .B(n2018), .Y(n1793) );
  NOR2X1 U2164 ( .A(n2017), .B(n2016), .Y(n2019) );
  MXI2X1 U2165 ( .A(n2568), .B(n2015), .S0(n2152), .Y(n2018) );
  NOR2X1 U2166 ( .A(n2130), .B(\register[1][14] ), .Y(n2017) );
  NAND2X1 U2167 ( .A(n2014), .B(n2013), .Y(n1801) );
  NOR2X1 U2168 ( .A(n2012), .B(n2011), .Y(n2014) );
  MXI2X1 U2169 ( .A(n2569), .B(n2010), .S0(n2153), .Y(n2013) );
  NOR2X1 U2170 ( .A(n2131), .B(\register[1][15] ), .Y(n2012) );
  NAND2X1 U2171 ( .A(n2009), .B(n2008), .Y(n1809) );
  NOR2X1 U2172 ( .A(n2007), .B(n2006), .Y(n2009) );
  MXI2X1 U2173 ( .A(n2570), .B(n2005), .S0(n2153), .Y(n2008) );
  NOR2X1 U2174 ( .A(n2131), .B(\register[1][16] ), .Y(n2007) );
  NAND2X1 U2175 ( .A(n2004), .B(n2003), .Y(n1817) );
  NOR2X1 U2176 ( .A(n2002), .B(n2001), .Y(n2004) );
  MXI2X1 U2177 ( .A(n2571), .B(n2000), .S0(n2153), .Y(n2003) );
  NOR2X1 U2178 ( .A(n2131), .B(\register[1][17] ), .Y(n2002) );
  NAND2X1 U2179 ( .A(n1999), .B(n1998), .Y(n1825) );
  NOR2X1 U2180 ( .A(n1997), .B(n1996), .Y(n1999) );
  MXI2X1 U2181 ( .A(n2572), .B(n1995), .S0(n2153), .Y(n1998) );
  NOR2X1 U2182 ( .A(n2131), .B(\register[1][18] ), .Y(n1997) );
  NAND2X1 U2183 ( .A(n1994), .B(n1993), .Y(n1833) );
  NOR2X1 U2184 ( .A(n1992), .B(n1991), .Y(n1994) );
  MXI2X1 U2185 ( .A(n2573), .B(n1990), .S0(n2153), .Y(n1993) );
  NOR2X1 U2186 ( .A(n2131), .B(\register[1][19] ), .Y(n1992) );
  NAND2X1 U2187 ( .A(n1989), .B(n1988), .Y(n1841) );
  NOR2X1 U2188 ( .A(n1987), .B(n1986), .Y(n1989) );
  NAND2X1 U2189 ( .A(n1984), .B(n1983), .Y(n1849) );
  NOR2X1 U2190 ( .A(n1982), .B(n1981), .Y(n1984) );
  MXI2X1 U2191 ( .A(n2575), .B(n1980), .S0(n2153), .Y(n1983) );
  NOR2X1 U2192 ( .A(n2132), .B(\register[1][21] ), .Y(n1982) );
  NAND2X1 U2193 ( .A(n1979), .B(n1978), .Y(n1857) );
  NOR2X1 U2194 ( .A(n1977), .B(n1976), .Y(n1979) );
  MXI2X1 U2195 ( .A(n2576), .B(n1975), .S0(n2153), .Y(n1978) );
  NOR2X1 U2196 ( .A(n2132), .B(\register[1][22] ), .Y(n1977) );
  NAND2X1 U2197 ( .A(n1974), .B(n1973), .Y(n1865) );
  NOR2X1 U2198 ( .A(n1972), .B(n1971), .Y(n1974) );
  MXI2X1 U2199 ( .A(n2577), .B(n1970), .S0(n2153), .Y(n1973) );
  NOR2X1 U2200 ( .A(n2132), .B(\register[1][23] ), .Y(n1972) );
  NAND2X1 U2201 ( .A(n1969), .B(n1968), .Y(n1873) );
  NOR2X1 U2202 ( .A(n1967), .B(n1966), .Y(n1969) );
  MXI2X1 U2203 ( .A(n2578), .B(n1965), .S0(n2153), .Y(n1968) );
  NOR2X1 U2204 ( .A(n2132), .B(\register[1][24] ), .Y(n1967) );
  NAND2X1 U2205 ( .A(n1959), .B(n1958), .Y(n1889) );
  NOR2X1 U2206 ( .A(n1957), .B(n1956), .Y(n1959) );
  MXI2X1 U2207 ( .A(n2580), .B(n1955), .S0(n2153), .Y(n1958) );
  NOR2X1 U2208 ( .A(n2132), .B(\register[1][26] ), .Y(n1957) );
  NAND2X1 U2209 ( .A(n1944), .B(n1943), .Y(n1913) );
  NOR2X1 U2210 ( .A(n1942), .B(n1941), .Y(n1944) );
  MXI2X1 U2211 ( .A(n2583), .B(n1940), .S0(n2153), .Y(n1943) );
  NOR2X1 U2212 ( .A(n2133), .B(\register[1][29] ), .Y(n1942) );
  NAND2X1 U2213 ( .A(n1934), .B(n1933), .Y(n1929) );
  NOR2X1 U2214 ( .A(n1932), .B(n1931), .Y(n1934) );
  MXI2X1 U2215 ( .A(n2585), .B(n1930), .S0(n2153), .Y(n1933) );
  NOR2X1 U2216 ( .A(n2133), .B(\register[1][31] ), .Y(n1932) );
  NAND2X1 U2217 ( .A(n1535), .B(n1534), .Y(n1153) );
  NOR2X1 U2218 ( .A(n1533), .B(n1532), .Y(n1535) );
  MXI2X1 U2219 ( .A(n2556), .B(n1531), .S0(n1607), .Y(n1534) );
  NOR2X1 U2220 ( .A(n1586), .B(\register[1][2] ), .Y(n1533) );
  NAND2X1 U2221 ( .A(n1530), .B(n1529), .Y(n1161) );
  NOR2X1 U2222 ( .A(n1528), .B(n1527), .Y(n1530) );
  MXI2X1 U2223 ( .A(n2557), .B(n1526), .S0(n1607), .Y(n1529) );
  NOR2X1 U2224 ( .A(n1585), .B(\register[1][3] ), .Y(n1528) );
  NAND2X1 U2225 ( .A(n1525), .B(n1524), .Y(n1169) );
  NOR2X1 U2226 ( .A(n1523), .B(n1522), .Y(n1525) );
  MXI2X1 U2227 ( .A(n2558), .B(n1521), .S0(n1607), .Y(n1524) );
  NOR2X1 U2228 ( .A(n1584), .B(\register[1][4] ), .Y(n1523) );
  NAND2X1 U2229 ( .A(n1520), .B(n1519), .Y(n1177) );
  NOR2X1 U2230 ( .A(n1518), .B(n1517), .Y(n1520) );
  MXI2X1 U2231 ( .A(n2559), .B(n1516), .S0(n1607), .Y(n1519) );
  NOR2X1 U2232 ( .A(n1585), .B(\register[1][5] ), .Y(n1518) );
  NAND2X1 U2233 ( .A(n1515), .B(n1514), .Y(n1185) );
  NOR2X1 U2234 ( .A(n1513), .B(n1512), .Y(n1515) );
  MXI2X1 U2235 ( .A(n2560), .B(n1511), .S0(n1607), .Y(n1514) );
  NOR2X1 U2236 ( .A(n1584), .B(\register[1][6] ), .Y(n1513) );
  NAND2X1 U2237 ( .A(n1510), .B(n1509), .Y(n1193) );
  NOR2X1 U2238 ( .A(n1508), .B(n1507), .Y(n1510) );
  MXI2X1 U2239 ( .A(n2561), .B(n1506), .S0(n1607), .Y(n1509) );
  NOR2X1 U2240 ( .A(n1585), .B(\register[1][7] ), .Y(n1508) );
  NAND2X1 U2241 ( .A(n1505), .B(n1504), .Y(n1201) );
  NOR2X1 U2242 ( .A(n1503), .B(n1502), .Y(n1505) );
  MXI2X1 U2243 ( .A(n2562), .B(n1501), .S0(n1607), .Y(n1504) );
  NOR2X1 U2244 ( .A(n1586), .B(\register[1][8] ), .Y(n1503) );
  NAND2X1 U2245 ( .A(n1500), .B(n1499), .Y(n1209) );
  NOR2X1 U2246 ( .A(n1498), .B(n1497), .Y(n1500) );
  MXI2X1 U2247 ( .A(n2563), .B(n1496), .S0(n1607), .Y(n1499) );
  NOR2X1 U2248 ( .A(n1585), .B(\register[1][9] ), .Y(n1498) );
  NAND2X1 U2249 ( .A(n1495), .B(n1494), .Y(n1217) );
  NOR2X1 U2250 ( .A(n1493), .B(n1492), .Y(n1495) );
  MXI2X1 U2251 ( .A(n2564), .B(n1491), .S0(n1607), .Y(n1494) );
  NOR2X1 U2252 ( .A(n1585), .B(\register[1][10] ), .Y(n1493) );
  NAND2X1 U2253 ( .A(n1490), .B(n1489), .Y(n1225) );
  NOR2X1 U2254 ( .A(n1488), .B(n1487), .Y(n1490) );
  MXI2X1 U2255 ( .A(n2565), .B(n1486), .S0(n1607), .Y(n1489) );
  NOR2X1 U2256 ( .A(n1586), .B(\register[1][11] ), .Y(n1488) );
  NAND2X1 U2257 ( .A(n1485), .B(n1484), .Y(n1233) );
  NOR2X1 U2258 ( .A(n1483), .B(n1482), .Y(n1485) );
  MXI2X1 U2259 ( .A(n2566), .B(n1481), .S0(n1607), .Y(n1484) );
  NOR2X1 U2260 ( .A(n1586), .B(\register[1][12] ), .Y(n1483) );
  NAND2X1 U2261 ( .A(n1480), .B(n1479), .Y(n1241) );
  NOR2X1 U2262 ( .A(n1478), .B(n1477), .Y(n1480) );
  MXI2X1 U2263 ( .A(n2567), .B(n1476), .S0(n1607), .Y(n1479) );
  NOR2X1 U2264 ( .A(n1586), .B(\register[1][13] ), .Y(n1478) );
  NAND2X1 U2265 ( .A(n1475), .B(n1474), .Y(n1249) );
  NOR2X1 U2266 ( .A(n1473), .B(n1472), .Y(n1475) );
  NOR2X1 U2267 ( .A(n1586), .B(\register[1][14] ), .Y(n1473) );
  NAND2X1 U2268 ( .A(n1470), .B(n1469), .Y(n1257) );
  NOR2X1 U2269 ( .A(n1468), .B(n1467), .Y(n1470) );
  MXI2X1 U2270 ( .A(n2569), .B(n1466), .S0(n1608), .Y(n1469) );
  NOR2X1 U2271 ( .A(n1587), .B(\register[1][15] ), .Y(n1468) );
  NAND2X1 U2272 ( .A(n1465), .B(n1464), .Y(n1265) );
  NOR2X1 U2273 ( .A(n1463), .B(n1462), .Y(n1465) );
  MXI2X1 U2274 ( .A(n2570), .B(n1461), .S0(n1608), .Y(n1464) );
  NOR2X1 U2275 ( .A(n1587), .B(\register[1][16] ), .Y(n1463) );
  NAND2X1 U2276 ( .A(n1460), .B(n1459), .Y(n1273) );
  NOR2X1 U2277 ( .A(n1458), .B(n1457), .Y(n1460) );
  MXI2X1 U2278 ( .A(n2571), .B(n1456), .S0(n1608), .Y(n1459) );
  NOR2X1 U2279 ( .A(n1587), .B(\register[1][17] ), .Y(n1458) );
  NAND2X1 U2280 ( .A(n1455), .B(n1454), .Y(n1281) );
  NOR2X1 U2281 ( .A(n1453), .B(n1452), .Y(n1455) );
  MXI2X1 U2282 ( .A(n2572), .B(n1451), .S0(n1608), .Y(n1454) );
  NOR2X1 U2283 ( .A(n1587), .B(\register[1][18] ), .Y(n1453) );
  NAND2X1 U2284 ( .A(n1450), .B(n1449), .Y(n1289) );
  NOR2X1 U2285 ( .A(n1448), .B(n1447), .Y(n1450) );
  MXI2X1 U2286 ( .A(n2573), .B(n1446), .S0(n1608), .Y(n1449) );
  NOR2X1 U2287 ( .A(n1587), .B(\register[1][19] ), .Y(n1448) );
  NAND2X1 U2288 ( .A(n1445), .B(n1444), .Y(n1297) );
  NOR2X1 U2289 ( .A(n1443), .B(n1442), .Y(n1445) );
  MXI2X1 U2290 ( .A(n2574), .B(n1441), .S0(n1608), .Y(n1444) );
  NOR2X1 U2291 ( .A(n1587), .B(\register[1][20] ), .Y(n1443) );
  NAND2X1 U2292 ( .A(n1440), .B(n1439), .Y(n1305) );
  NOR2X1 U2293 ( .A(n1438), .B(n1437), .Y(n1440) );
  MXI2X1 U2294 ( .A(n2575), .B(n1436), .S0(n1608), .Y(n1439) );
  NOR2X1 U2295 ( .A(n1583), .B(\register[1][21] ), .Y(n1438) );
  NAND2X1 U2296 ( .A(n1435), .B(n1434), .Y(n1313) );
  NOR2X1 U2297 ( .A(n1433), .B(n1432), .Y(n1435) );
  MXI2X1 U2298 ( .A(n2576), .B(n1431), .S0(n1608), .Y(n1434) );
  NOR2X1 U2299 ( .A(n1583), .B(\register[1][22] ), .Y(n1433) );
  NAND2X1 U2300 ( .A(n1430), .B(n1429), .Y(n1321) );
  NOR2X1 U2301 ( .A(n1428), .B(n1427), .Y(n1430) );
  MXI2X1 U2302 ( .A(n2577), .B(n1426), .S0(n1608), .Y(n1429) );
  NOR2X1 U2303 ( .A(n1583), .B(\register[1][23] ), .Y(n1428) );
  NAND2X1 U2304 ( .A(n1425), .B(n1424), .Y(n1329) );
  NOR2X1 U2305 ( .A(n1423), .B(n1422), .Y(n1425) );
  MXI2X1 U2306 ( .A(n2578), .B(n1421), .S0(n1608), .Y(n1424) );
  NOR2X1 U2307 ( .A(n1577), .B(\register[1][24] ), .Y(n1423) );
  NAND2X1 U2308 ( .A(n1415), .B(n1414), .Y(n1345) );
  NOR2X1 U2309 ( .A(n1413), .B(n1412), .Y(n1415) );
  MXI2X1 U2310 ( .A(n2580), .B(n1411), .S0(n1608), .Y(n1414) );
  NOR2X1 U2311 ( .A(n1588), .B(n1609), .Y(n1412) );
  NAND2X1 U2312 ( .A(n1400), .B(n1399), .Y(n1369) );
  NOR2X1 U2313 ( .A(n1398), .B(n1397), .Y(n1400) );
  MXI2X1 U2314 ( .A(n2583), .B(n1396), .S0(n1608), .Y(n1399) );
  NOR2X1 U2315 ( .A(n1588), .B(\register[1][29] ), .Y(n1398) );
  NAND2X1 U2316 ( .A(n1390), .B(n1389), .Y(n1385) );
  NOR2X1 U2317 ( .A(n1388), .B(n1387), .Y(n1390) );
  MXI2X1 U2318 ( .A(n2585), .B(n1386), .S0(n1608), .Y(n1389) );
  NOR2X1 U2319 ( .A(n1588), .B(\register[1][31] ), .Y(n1388) );
  NAND2X1 U2320 ( .A(n2089), .B(n2088), .Y(n1681) );
  NOR2X1 U2321 ( .A(n2087), .B(n2086), .Y(n2089) );
  MXI2X1 U2322 ( .A(n2554), .B(n2085), .S0(n2151), .Y(n2088) );
  NOR2X1 U2323 ( .A(n2133), .B(\register[1][0] ), .Y(n2087) );
  NAND2X1 U2324 ( .A(n1964), .B(n1963), .Y(n1881) );
  NOR2X1 U2325 ( .A(n1962), .B(n1961), .Y(n1964) );
  MXI2X1 U2326 ( .A(n2579), .B(n1960), .S0(n2145), .Y(n1963) );
  NOR2X1 U2327 ( .A(n2132), .B(\register[1][25] ), .Y(n1962) );
  NAND2X1 U2328 ( .A(n1954), .B(n1953), .Y(n1897) );
  NOR2X1 U2329 ( .A(n1952), .B(n1951), .Y(n1954) );
  MXI2X1 U2330 ( .A(n2581), .B(n1950), .S0(n2145), .Y(n1953) );
  NOR2X1 U2331 ( .A(n2133), .B(\register[1][27] ), .Y(n1952) );
  NAND2X1 U2332 ( .A(n1949), .B(n1948), .Y(n1905) );
  NOR2X1 U2333 ( .A(n1947), .B(n1946), .Y(n1949) );
  MXI2X1 U2334 ( .A(n2582), .B(n1945), .S0(n2145), .Y(n1948) );
  NOR2X1 U2335 ( .A(n2133), .B(\register[1][28] ), .Y(n1947) );
  NAND2X1 U2336 ( .A(n1939), .B(n1938), .Y(n1921) );
  NOR2X1 U2337 ( .A(n1937), .B(n1936), .Y(n1939) );
  MXI2X1 U2338 ( .A(n2584), .B(n1935), .S0(n2145), .Y(n1938) );
  NOR2X1 U2339 ( .A(n2133), .B(\register[1][30] ), .Y(n1937) );
  NAND2X1 U2340 ( .A(n1545), .B(n1544), .Y(n1137) );
  NOR2X1 U2341 ( .A(n1543), .B(n1542), .Y(n1545) );
  MXI2X1 U2342 ( .A(n2554), .B(n1541), .S0(n1599), .Y(n1544) );
  NOR2X1 U2343 ( .A(n1588), .B(\register[1][0] ), .Y(n1543) );
  NAND2X1 U2344 ( .A(n1420), .B(n1419), .Y(n1337) );
  NOR2X1 U2345 ( .A(n1418), .B(n1417), .Y(n1420) );
  MXI2X1 U2346 ( .A(n2579), .B(n1416), .S0(n1599), .Y(n1419) );
  NOR2X1 U2347 ( .A(n1573), .B(\register[1][25] ), .Y(n1418) );
  NAND2X1 U2348 ( .A(n1410), .B(n1409), .Y(n1353) );
  NOR2X1 U2349 ( .A(n1408), .B(n1407), .Y(n1410) );
  MXI2X1 U2350 ( .A(n2581), .B(n1406), .S0(n1599), .Y(n1409) );
  NOR2X1 U2351 ( .A(n1588), .B(\register[1][27] ), .Y(n1408) );
  NAND2X1 U2352 ( .A(n1405), .B(n1404), .Y(n1361) );
  NOR2X1 U2353 ( .A(n1403), .B(n1402), .Y(n1405) );
  MXI2X1 U2354 ( .A(n2582), .B(n1401), .S0(n1599), .Y(n1404) );
  NOR2X1 U2355 ( .A(n1588), .B(\register[1][28] ), .Y(n1403) );
  NAND2X1 U2356 ( .A(n1395), .B(n1394), .Y(n1377) );
  NOR2X1 U2357 ( .A(n1393), .B(n1392), .Y(n1395) );
  MXI2X1 U2358 ( .A(n2584), .B(n1391), .S0(n1599), .Y(n1394) );
  NOR2X1 U2359 ( .A(n1588), .B(\register[1][30] ), .Y(n1393) );
  MXI4X1 U2360 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n2145), .S1(n2122), .Y(
        n1680) );
  MXI4X1 U2361 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n2145), .S1(n2122), .Y(
        n1676) );
  MXI4X1 U2362 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n2146), .S1(n2122), .Y(
        n1684) );
  MXI4X1 U2363 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n2146), .S1(n2122), .Y(
        n1688) );
  MXI4X1 U2364 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n2146), .S1(n2122), .Y(
        n1692) );
  MXI4X1 U2365 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n2146), .S1(n2122), .Y(
        n1696) );
  MXI4X1 U2366 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n2146), .S1(n2123), .Y(
        n1700) );
  MXI4X1 U2367 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n2147), .S1(n2123), .Y(
        n1704) );
  MXI4X1 U2368 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n2147), .S1(n2123), .Y(
        n1708) );
  MXI4X1 U2369 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n2147), .S1(n2123), .Y(
        n1712) );
  MXI4X1 U2370 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n2148), .S1(n2123), .Y(
        n1720) );
  MXI4X1 U2371 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n2147), .S1(n2123), .Y(
        n1716) );
  MXI4X1 U2372 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n2148), .S1(n2124), .Y(
        n1724) );
  MXI4X1 U2373 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n2148), .S1(n2124), .Y(
        n1728) );
  MXI4X1 U2374 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n2149), .S1(n2124), .Y(
        n1744) );
  MXI4X1 U2375 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n2149), .S1(n2124), .Y(
        n1740) );
  MXI4X1 U2376 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n2150), .S1(n2125), .Y(
        n1752) );
  MXI4X1 U2377 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n2149), .S1(n2125), .Y(
        n1748) );
  MXI4X1 U2378 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n2150), .S1(n2125), .Y(
        n1760) );
  MXI4X1 U2379 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1756) );
  MXI4X1 U2380 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n2145), .S1(n2125), .Y(
        n1768) );
  MXI4X1 U2381 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1764) );
  MXI4X1 U2382 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n2152), .S1(n2126), 
        .Y(n1772) );
  MXI4X1 U2383 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n2149), .S1(n2124), .Y(
        n1776) );
  MXI4X1 U2384 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n2145), .S1(n2126), .Y(
        n1784) );
  MXI4X1 U2385 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n2151), .S1(n2126), 
        .Y(n1780) );
  MXI4X1 U2386 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n2151), .S1(n2126), .Y(
        n1792) );
  MXI4X1 U2387 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1788) );
  MXI4X1 U2388 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n2149), .S1(n2124), .Y(
        n1800) );
  MXI4X1 U2389 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n2151), .S1(n2126), 
        .Y(n1796) );
  MXI4X1 U2390 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n2141), .S1(n2117), .Y(
        n1808) );
  MXI4X1 U2391 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1804) );
  MXI4X1 U2392 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n2141), .S1(n2117), .Y(
        n1816) );
  MXI4X1 U2393 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1812) );
  MXI4X1 U2394 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n2142), .S1(n2117), .Y(
        n1824) );
  MXI4X1 U2395 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n2142), .S1(n2117), 
        .Y(n1820) );
  MXI4X1 U2396 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n2142), .S1(n2118), .Y(
        n1832) );
  MXI4X1 U2397 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n2142), .S1(n2118), 
        .Y(n1828) );
  MXI4X1 U2398 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n2145), .S1(n2118), .Y(
        n1848) );
  MXI4X1 U2399 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1844) );
  MXI4X1 U2400 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n2145), .S1(n2119), .Y(
        n1856) );
  MXI4X1 U2401 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n2145), .S1(n2119), 
        .Y(n1852) );
  MXI4X1 U2402 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n2145), .S1(n2119), .Y(
        n1864) );
  MXI4X1 U2403 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1860) );
  MXI4X1 U2404 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n2143), .S1(n2119), .Y(
        n1872) );
  MXI4X1 U2405 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n2145), .S1(n2119), 
        .Y(n1868) );
  MXI4X1 U2406 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n2143), .S1(n2120), .Y(
        n1880) );
  MXI4X1 U2407 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n2143), .S1(n2120), 
        .Y(n1876) );
  MXI4X1 U2408 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n2144), .S1(n2120), .Y(
        n1888) );
  MXI4X1 U2409 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n2143), .S1(n2120), 
        .Y(n1884) );
  MXI4X1 U2410 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n2144), .S1(n2120), .Y(
        n1896) );
  MXI4X1 U2411 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1892) );
  MXI4X1 U2412 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n2145), .S1(n2121), .Y(
        n1904) );
  MXI4X1 U2413 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n2144), .S1(n2120), 
        .Y(n1900) );
  MXI4X1 U2414 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n2145), .S1(n2121), .Y(
        n1912) );
  MXI4X1 U2415 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1908) );
  MXI4X1 U2416 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n2145), .S1(n2121), .Y(
        n1920) );
  MXI4X1 U2417 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1916) );
  MXI4X1 U2418 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n2145), .S1(n2121), 
        .Y(n1924) );
  MXI4X1 U2419 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n1599), .S1(n1578), .Y(
        n1136) );
  MXI4X1 U2420 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1599), .S1(n1578), .Y(
        n1132) );
  MXI4X1 U2421 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1600), .S1(n1578), .Y(
        n1148) );
  MXI4X1 U2422 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n1600), .S1(n1578), .Y(
        n1152) );
  MXI4X1 U2423 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1600), .S1(n1579), .Y(
        n1156) );
  MXI4X1 U2424 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n1601), .S1(n1579), .Y(
        n1160) );
  MXI4X1 U2425 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1601), .S1(n1579), .Y(
        n1164) );
  MXI4X1 U2426 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n1601), .S1(n1579), .Y(
        n1168) );
  MXI4X1 U2427 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n1602), .S1(n1579), .Y(
        n1176) );
  MXI4X1 U2428 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1601), .S1(n1579), .Y(
        n1172) );
  MXI4X1 U2429 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1602), .S1(n1580), .Y(
        n1180) );
  MXI4X1 U2430 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n1602), .S1(n1580), .Y(
        n1184) );
  MXI4X1 U2431 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1603), .S1(n1580), .Y(
        n1192) );
  MXI4X1 U2432 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1602), .S1(n1580), .Y(
        n1188) );
  MXI4X1 U2433 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1603), .S1(n1580), .Y(
        n1200) );
  MXI4X1 U2434 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1603), .S1(n1580), .Y(
        n1196) );
  MXI4X1 U2435 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1604), .S1(n1581), .Y(
        n1208) );
  MXI4X1 U2436 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1603), .S1(n1581), .Y(
        n1204) );
  MXI4X1 U2437 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1604), .S1(n1581), .Y(
        n1216) );
  MXI4X1 U2438 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1212) );
  MXI4X1 U2439 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1605), .S1(n1581), .Y(
        n1224) );
  MXI4X1 U2440 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1220) );
  MXI4X1 U2441 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1605), .S1(n1582), 
        .Y(n1228) );
  MXI4X1 U2442 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1603), .S1(n1580), .Y(
        n1232) );
  MXI4X1 U2443 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1605), .S1(n1582), .Y(
        n1240) );
  MXI4X1 U2444 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1236) );
  MXI4X1 U2445 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1603), .S1(n1580), .Y(
        n1256) );
  MXI4X1 U2446 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1606), .S1(n1582), 
        .Y(n1252) );
  MXI4X1 U2447 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1595), .S1(n1573), .Y(
        n1264) );
  MXI4X1 U2448 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1260) );
  MXI4X1 U2449 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1595), .S1(n1573), .Y(
        n1272) );
  MXI4X1 U2450 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1268) );
  MXI4X1 U2451 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1599), .S1(n1573), .Y(
        n1280) );
  MXI4X1 U2452 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1599), .S1(n1573), 
        .Y(n1276) );
  MXI4X1 U2453 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1599), .S1(n1574), .Y(
        n1288) );
  MXI4X1 U2454 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1599), .S1(n1574), 
        .Y(n1284) );
  MXI4X1 U2455 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1599), .S1(n1574), .Y(
        n1296) );
  MXI4X1 U2456 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1292) );
  MXI4X1 U2457 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1599), .S1(n1574), .Y(
        n1304) );
  MXI4X1 U2458 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1599), .S1(n1574), 
        .Y(n1300) );
  MXI4X1 U2459 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1596), .S1(n1575), .Y(
        n1312) );
  MXI4X1 U2460 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1599), .S1(n1575), 
        .Y(n1308) );
  MXI4X1 U2461 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1596), .S1(n1575), .Y(
        n1320) );
  MXI4X1 U2462 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1316) );
  MXI4X1 U2463 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1597), .S1(n1575), .Y(
        n1328) );
  MXI4X1 U2464 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1596), .S1(n1575), 
        .Y(n1324) );
  MXI4X1 U2465 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1597), .S1(n1576), .Y(
        n1336) );
  MXI4X1 U2466 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1597), .S1(n1576), 
        .Y(n1332) );
  MXI4X1 U2467 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1598), .S1(n1576), .Y(
        n1344) );
  MXI4X1 U2468 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1597), .S1(n1576), 
        .Y(n1340) );
  MXI4X1 U2469 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1598), .S1(n1576), .Y(
        n1352) );
  MXI4X1 U2470 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1348) );
  MXI4X1 U2471 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1599), .S1(n1577), .Y(
        n1360) );
  MXI4X1 U2472 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1598), .S1(n1576), 
        .Y(n1356) );
  MXI4X1 U2473 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1599), .S1(n1577), .Y(
        n1368) );
  MXI4X1 U2474 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1599), .S1(n1577), 
        .Y(n1364) );
  MXI4X1 U2475 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1599), .S1(n1577), .Y(
        n1376) );
  MXI4X1 U2476 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1599), .S1(n1577), 
        .Y(n1372) );
  MXI4X1 U2477 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1606), .S1(n1583), .Y(
        n1384) );
  MXI4X1 U2478 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1599), .S1(n1577), 
        .Y(n1380) );
  MXI4X1 U2479 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n2146), .S1(n2122), .Y(
        n1685) );
  MXI4X1 U2480 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n2146), .S1(n2122), .Y(
        n1693) );
  MXI4X1 U2481 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n2147), .S1(n2123), .Y(
        n1701) );
  MXI4X1 U2482 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n2147), .S1(n2123), .Y(
        n1709) );
  MXI4X1 U2483 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n2148), .S1(n2124), .Y(
        n1725) );
  MXI4X1 U2484 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n2145), .S1(n2126), 
        .Y(n1773) );
  MXI4X1 U2485 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1600), .S1(n1578), .Y(
        n1149) );
  MXI4X1 U2486 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1601), .S1(n1579), .Y(
        n1157) );
  MXI4X1 U2487 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1601), .S1(n1579), .Y(
        n1165) );
  MXI4X1 U2488 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1602), .S1(n1580), .Y(
        n1181) );
  MXI4X1 U2489 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1605), .S1(n1582), 
        .Y(n1229) );
  MXI4X1 U2490 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n2145), .S1(n2122), .Y(
        n1678) );
  MXI4X1 U2491 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n2145), .S1(n2122), .Y(
        n1674) );
  MXI4X1 U2492 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n2145), .S1(n2122), .Y(
        n1682) );
  MXI4X1 U2493 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n2146), .S1(n2122), .Y(
        n1686) );
  MXI4X1 U2494 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n2146), .S1(n2122), .Y(
        n1690) );
  MXI4X1 U2495 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n2146), .S1(n2122), .Y(
        n1694) );
  MXI4X1 U2496 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n2146), .S1(n2123), .Y(
        n1698) );
  MXI4X1 U2497 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n2147), .S1(n2123), .Y(
        n1702) );
  MXI4X1 U2498 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n2147), .S1(n2123), .Y(
        n1706) );
  MXI4X1 U2499 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n2147), .S1(n2123), .Y(
        n1710) );
  MXI4X1 U2500 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n2148), .S1(n2123), .Y(
        n1718) );
  MXI4X1 U2501 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n2147), .S1(n2123), .Y(
        n1714) );
  MXI4X1 U2502 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n2148), .S1(n2123), .Y(
        n1722) );
  MXI4X1 U2503 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n2148), .S1(n2124), .Y(
        n1726) );
  MXI4X1 U2504 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n2149), .S1(n2124), .Y(
        n1742) );
  MXI4X1 U2505 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n2149), .S1(n2125), .Y(
        n1750) );
  MXI4X1 U2506 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n2149), .S1(n2124), .Y(
        n1746) );
  MXI4X1 U2507 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1758) );
  MXI4X1 U2508 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1754) );
  MXI4X1 U2509 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1766) );
  MXI4X1 U2510 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1762) );
  MXI4X1 U2511 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n2136), .S1(n2125), 
        .Y(n1770) );
  MXI4X1 U2512 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n2150), .S1(n2126), 
        .Y(n1774) );
  MXI4X1 U2513 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n2145), .S1(n2126), 
        .Y(n1782) );
  MXI4X1 U2514 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n2152), .S1(n2126), 
        .Y(n1778) );
  MXI4X1 U2515 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1790) );
  MXI4X1 U2516 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1786) );
  MXI4X1 U2517 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n2151), .S1(n2126), 
        .Y(n1794) );
  MXI4X1 U2518 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1806) );
  MXI4X1 U2519 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1802) );
  MXI4X1 U2520 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1814) );
  MXI4X1 U2521 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1810) );
  MXI4X1 U2522 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n2142), .S1(n2117), 
        .Y(n1822) );
  MXI4X1 U2523 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n2141), .S1(n2117), 
        .Y(n1818) );
  MXI4X1 U2524 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n2142), .S1(n2118), 
        .Y(n1830) );
  MXI4X1 U2525 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n2142), .S1(n2117), 
        .Y(n1826) );
  MXI4X1 U2526 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1846) );
  MXI4X1 U2527 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1842) );
  MXI4X1 U2528 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n2145), .S1(n2119), 
        .Y(n1854) );
  MXI4X1 U2529 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n2145), .S1(n2118), 
        .Y(n1850) );
  MXI4X1 U2530 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1862) );
  MXI4X1 U2531 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1858) );
  MXI4X1 U2532 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n2143), .S1(n2119), 
        .Y(n1870) );
  MXI4X1 U2533 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n2145), .S1(n2119), 
        .Y(n1866) );
  MXI4X1 U2534 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n2143), .S1(n2120), 
        .Y(n1878) );
  MXI4X1 U2535 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n2143), .S1(n2119), 
        .Y(n1874) );
  MXI4X1 U2536 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n2144), .S1(n2120), 
        .Y(n1886) );
  MXI4X1 U2537 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n2143), .S1(n2120), 
        .Y(n1882) );
  MXI4X1 U2538 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1894) );
  MXI4X1 U2539 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1890) );
  MXI4X1 U2540 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n2144), .S1(n2121), 
        .Y(n1902) );
  MXI4X1 U2541 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n2144), .S1(n2120), 
        .Y(n1898) );
  MXI4X1 U2542 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1910) );
  MXI4X1 U2543 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1906) );
  MXI4X1 U2544 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1918) );
  MXI4X1 U2545 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1914) );
  MXI4X1 U2546 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n2145), .S1(n2122), 
        .Y(n1926) );
  MXI4X1 U2547 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n2145), .S1(n2121), 
        .Y(n1922) );
  MXI4X1 U2548 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1599), .S1(n1578), .Y(
        n1134) );
  MXI4X1 U2549 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1599), .S1(n1578), .Y(
        n1130) );
  MXI4X1 U2550 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1600), .S1(n1578), .Y(
        n1146) );
  MXI4X1 U2551 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1600), .S1(n1578), .Y(
        n1150) );
  MXI4X1 U2552 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1600), .S1(n1579), .Y(
        n1154) );
  MXI4X1 U2553 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1601), .S1(n1579), .Y(
        n1158) );
  MXI4X1 U2554 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1601), .S1(n1579), .Y(
        n1162) );
  MXI4X1 U2555 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1601), .S1(n1579), .Y(
        n1166) );
  MXI4X1 U2556 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1602), .S1(n1579), .Y(
        n1174) );
  MXI4X1 U2557 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1601), .S1(n1579), .Y(
        n1170) );
  MXI4X1 U2558 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1602), .S1(n1579), .Y(
        n1178) );
  MXI4X1 U2559 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1602), .S1(n1580), .Y(
        n1182) );
  MXI4X1 U2560 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1602), .S1(n1580), .Y(
        n1190) );
  MXI4X1 U2561 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1602), .S1(n1580), .Y(
        n1186) );
  MXI4X1 U2562 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1603), .S1(n1580), .Y(
        n1198) );
  MXI4X1 U2563 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1606), .S1(n1583), .Y(
        n1194) );
  MXI4X1 U2564 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1603), .S1(n1581), .Y(
        n1206) );
  MXI4X1 U2565 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1603), .S1(n1580), .Y(
        n1202) );
  MXI4X1 U2566 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1214) );
  MXI4X1 U2567 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1210) );
  MXI4X1 U2568 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1222) );
  MXI4X1 U2569 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1218) );
  MXI4X1 U2570 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1605), .S1(n1581), 
        .Y(n1226) );
  MXI4X1 U2571 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1605), .S1(n1582), 
        .Y(n1230) );
  MXI4X1 U2572 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1238) );
  MXI4X1 U2573 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1234) );
  MXI4X1 U2574 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1606), .S1(n1583), 
        .Y(n1254) );
  MXI4X1 U2575 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1606), .S1(n1582), 
        .Y(n1250) );
  MXI4X1 U2576 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1262) );
  MXI4X1 U2577 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1258) );
  MXI4X1 U2578 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1270) );
  MXI4X1 U2579 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1266) );
  MXI4X1 U2580 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1599), .S1(n1573), 
        .Y(n1278) );
  MXI4X1 U2581 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1595), .S1(n1573), 
        .Y(n1274) );
  MXI4X1 U2582 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1599), .S1(n1574), 
        .Y(n1286) );
  MXI4X1 U2583 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1599), .S1(n1573), 
        .Y(n1282) );
  MXI4X1 U2584 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1294) );
  MXI4X1 U2585 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1290) );
  MXI4X1 U2586 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1599), .S1(n1574), 
        .Y(n1302) );
  MXI4X1 U2587 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1596), .S1(n1574), 
        .Y(n1298) );
  MXI4X1 U2588 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1596), .S1(n1575), 
        .Y(n1310) );
  MXI4X1 U2589 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1604), .S1(n1574), 
        .Y(n1306) );
  MXI4X1 U2590 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1318) );
  MXI4X1 U2591 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1314) );
  MXI4X1 U2592 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1597), .S1(n1575), 
        .Y(n1326) );
  MXI4X1 U2593 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1596), .S1(n1575), 
        .Y(n1322) );
  MXI4X1 U2594 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1597), .S1(n1576), 
        .Y(n1334) );
  MXI4X1 U2595 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1597), .S1(n1575), 
        .Y(n1330) );
  MXI4X1 U2596 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1598), .S1(n1576), 
        .Y(n1342) );
  MXI4X1 U2597 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1597), .S1(n1576), 
        .Y(n1338) );
  MXI4X1 U2598 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1350) );
  MXI4X1 U2599 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1346) );
  MXI4X1 U2600 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1598), .S1(n1577), 
        .Y(n1358) );
  MXI4X1 U2601 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1598), .S1(n1576), 
        .Y(n1354) );
  MXI4X1 U2602 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1599), .S1(n1577), 
        .Y(n1366) );
  MXI4X1 U2603 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1598), .S1(n1577), 
        .Y(n1362) );
  MXI4X1 U2604 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1599), .S1(n1577), 
        .Y(n1374) );
  MXI4X1 U2605 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1597), .S1(n1577), 
        .Y(n1370) );
  MXI4X1 U2606 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1599), .S1(n1578), 
        .Y(n1382) );
  MXI4X1 U2607 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1599), .S1(n1577), 
        .Y(n1378) );
  MXI4X1 U2608 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n2145), .S1(n2122), .Y(
        n1679) );
  MXI4X1 U2609 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n2145), .S1(n2122), .Y(
        n1675) );
  MXI4X1 U2610 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n2145), .S1(n2122), .Y(
        n1683) );
  MXI4X1 U2611 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n2146), .S1(n2122), .Y(
        n1691) );
  MXI4X1 U2612 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n2146), .S1(n2123), .Y(
        n1699) );
  MXI4X1 U2613 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n2147), .S1(n2123), .Y(
        n1707) );
  MXI4X1 U2614 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n2148), .S1(n2123), .Y(
        n1719) );
  MXI4X1 U2615 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n2147), .S1(n2123), .Y(
        n1715) );
  MXI4X1 U2616 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n2148), .S1(n2124), .Y(
        n1723) );
  MXI4X1 U2617 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n2149), .S1(n2124), .Y(
        n1743) );
  MXI4X1 U2618 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n2149), .S1(n2124), .Y(
        n1739) );
  MXI4X1 U2619 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n2150), .S1(n2125), .Y(
        n1751) );
  MXI4X1 U2620 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n2149), .S1(n2125), .Y(
        n1747) );
  MXI4X1 U2621 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1759) );
  MXI4X1 U2622 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n2150), .S1(n2125), 
        .Y(n1755) );
  MXI4X1 U2623 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1767) );
  MXI4X1 U2624 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n2150), .S1(n2125), 
        .Y(n1763) );
  MXI4X1 U2625 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n2145), .S1(n2125), 
        .Y(n1771) );
  MXI4X1 U2626 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n2145), .S1(n2126), 
        .Y(n1783) );
  MXI4X1 U2627 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n2145), .S1(n2126), 
        .Y(n1779) );
  MXI4X1 U2628 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1791) );
  MXI4X1 U2629 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n2151), .S1(n2126), 
        .Y(n1787) );
  MXI4X1 U2630 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n2151), .S1(n2126), 
        .Y(n1795) );
  MXI4X1 U2631 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1807) );
  MXI4X1 U2632 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n2141), .S1(n2117), 
        .Y(n1803) );
  MXI4X1 U2633 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1815) );
  MXI4X1 U2634 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n2141), .S1(n2117), 
        .Y(n1811) );
  MXI4X1 U2635 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n2142), .S1(n2117), 
        .Y(n1823) );
  MXI4X1 U2636 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n2142), .S1(n2117), 
        .Y(n1819) );
  MXI4X1 U2637 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n2142), .S1(n2118), 
        .Y(n1831) );
  MXI4X1 U2638 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n2142), .S1(n2118), 
        .Y(n1827) );
  MXI4X1 U2639 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1847) );
  MXI4X1 U2640 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n2145), .S1(n2118), 
        .Y(n1843) );
  MXI4X1 U2641 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n2145), .S1(n2119), 
        .Y(n1855) );
  MXI4X1 U2642 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n2145), .S1(n2118), 
        .Y(n1851) );
  MXI4X1 U2643 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1863) );
  MXI4X1 U2644 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n2145), .S1(n2119), 
        .Y(n1859) );
  MXI4X1 U2645 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n2143), .S1(n2119), 
        .Y(n1871) );
  MXI4X1 U2646 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n2145), .S1(n2119), 
        .Y(n1867) );
  MXI4X1 U2647 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n2143), .S1(n2120), 
        .Y(n1879) );
  MXI4X1 U2648 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n2143), .S1(n2119), 
        .Y(n1875) );
  MXI4X1 U2649 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n2144), .S1(n2120), 
        .Y(n1887) );
  MXI4X1 U2650 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n2143), .S1(n2120), 
        .Y(n1883) );
  MXI4X1 U2651 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1895) );
  MXI4X1 U2652 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n2144), .S1(n2120), 
        .Y(n1891) );
  MXI4X1 U2653 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n2145), .S1(n2121), 
        .Y(n1903) );
  MXI4X1 U2654 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n2144), .S1(n2120), 
        .Y(n1899) );
  MXI4X1 U2655 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1911) );
  MXI4X1 U2656 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n2145), .S1(n2121), 
        .Y(n1907) );
  MXI4X1 U2657 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1919) );
  MXI4X1 U2658 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n2145), .S1(n2121), 
        .Y(n1915) );
  MXI4X1 U2659 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n2145), .S1(n2119), 
        .Y(n1927) );
  MXI4X1 U2660 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n2145), .S1(n2121), 
        .Y(n1923) );
  MXI4X1 U2661 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1599), .S1(n1578), .Y(
        n1135) );
  MXI4X1 U2662 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1599), .S1(n1578), .Y(
        n1131) );
  MXI4X1 U2663 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1600), .S1(n1578), .Y(
        n1147) );
  MXI4X1 U2664 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1600), .S1(n1579), .Y(
        n1155) );
  MXI4X1 U2665 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1601), .S1(n1579), .Y(
        n1163) );
  MXI4X1 U2666 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1602), .S1(n1579), .Y(
        n1175) );
  MXI4X1 U2667 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1601), .S1(n1579), .Y(
        n1171) );
  MXI4X1 U2668 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1602), .S1(n1580), .Y(
        n1179) );
  MXI4X1 U2669 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1603), .S1(n1580), .Y(
        n1191) );
  MXI4X1 U2670 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1602), .S1(n1580), .Y(
        n1187) );
  MXI4X1 U2671 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1603), .S1(n1580), .Y(
        n1199) );
  MXI4X1 U2672 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1603), .S1(n1580), .Y(
        n1195) );
  MXI4X1 U2673 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1604), .S1(n1581), .Y(
        n1207) );
  MXI4X1 U2674 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1603), .S1(n1581), .Y(
        n1203) );
  MXI4X1 U2675 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1215) );
  MXI4X1 U2676 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1604), .S1(n1581), 
        .Y(n1211) );
  MXI4X1 U2677 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1223) );
  MXI4X1 U2678 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1604), .S1(n1581), 
        .Y(n1219) );
  MXI4X1 U2679 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1605), .S1(n1581), 
        .Y(n1227) );
  MXI4X1 U2680 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1239) );
  MXI4X1 U2681 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1605), .S1(n1582), 
        .Y(n1235) );
  MXI4X1 U2682 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1606), .S1(n1583), 
        .Y(n1255) );
  MXI4X1 U2683 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1606), .S1(n1582), 
        .Y(n1251) );
  MXI4X1 U2684 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1263) );
  MXI4X1 U2685 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1595), .S1(n1573), 
        .Y(n1259) );
  MXI4X1 U2686 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1271) );
  MXI4X1 U2687 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1595), .S1(n1573), 
        .Y(n1267) );
  MXI4X1 U2688 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1599), .S1(n1573), 
        .Y(n1279) );
  MXI4X1 U2689 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1599), .S1(n1573), 
        .Y(n1275) );
  MXI4X1 U2690 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1599), .S1(n1574), 
        .Y(n1287) );
  MXI4X1 U2691 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1599), .S1(n1574), 
        .Y(n1283) );
  MXI4X1 U2692 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1295) );
  MXI4X1 U2693 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1599), .S1(n1574), 
        .Y(n1291) );
  MXI4X1 U2694 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1599), .S1(n1574), 
        .Y(n1303) );
  MXI4X1 U2695 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1599), .S1(n1574), 
        .Y(n1299) );
  MXI4X1 U2696 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1596), .S1(n1575), 
        .Y(n1311) );
  MXI4X1 U2697 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1599), .S1(n1574), 
        .Y(n1307) );
  MXI4X1 U2698 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1319) );
  MXI4X1 U2699 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1596), .S1(n1575), 
        .Y(n1315) );
  MXI4X1 U2700 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1597), .S1(n1575), 
        .Y(n1327) );
  MXI4X1 U2701 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1596), .S1(n1575), 
        .Y(n1323) );
  MXI4X1 U2702 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1597), .S1(n1576), 
        .Y(n1335) );
  MXI4X1 U2703 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1597), .S1(n1575), 
        .Y(n1331) );
  MXI4X1 U2704 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1598), .S1(n1576), 
        .Y(n1343) );
  MXI4X1 U2705 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1597), .S1(n1576), 
        .Y(n1339) );
  MXI4X1 U2706 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1351) );
  MXI4X1 U2707 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1598), .S1(n1576), 
        .Y(n1347) );
  MXI4X1 U2708 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1599), .S1(n1577), 
        .Y(n1359) );
  MXI4X1 U2709 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1598), .S1(n1576), 
        .Y(n1355) );
  MXI4X1 U2710 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1599), .S1(n1577), 
        .Y(n1367) );
  MXI4X1 U2711 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1599), .S1(n1577), 
        .Y(n1363) );
  MXI4X1 U2712 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1599), .S1(n1577), 
        .Y(n1375) );
  MXI4X1 U2713 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1599), .S1(n1577), 
        .Y(n1371) );
  MXI4X1 U2714 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1596), .S1(n1575), 
        .Y(n1383) );
  MXI4X1 U2715 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1599), .S1(n1577), 
        .Y(n1379) );
  XNOR2XL U2716 ( .A(n2444), .B(wsel[2]), .Y(n59) );
  XNOR2XL U2717 ( .A(n2440), .B(wsel[2]), .Y(n50) );
  XNOR2XL U2718 ( .A(n2443), .B(wsel[0]), .Y(n58) );
  XNOR2XL U2719 ( .A(n2439), .B(wsel[0]), .Y(n49) );
endmodule


module extender ( shamt_i, immed_i, ExtOp_i, ExtOut_o );
  input [4:0] shamt_i;
  input [15:0] immed_i;
  output [31:0] ExtOut_o;
  input ExtOp_i;
  wire   n2, n1, n19, n20;

  CLKINVX3 U1 ( .A(ExtOp_i), .Y(n20) );
  INVXL U2 ( .A(n1), .Y(ExtOut_o[15]) );
  OAI2BB1XL U3 ( .A0N(immed_i[13]), .A1N(n20), .B0(n19), .Y(ExtOut_o[13]) );
  OAI2BB1X4 U4 ( .A0N(immed_i[15]), .A1N(n20), .B0(n19), .Y(ExtOut_o[30]) );
  INVX3 U5 ( .A(ExtOut_o[30]), .Y(n1) );
  AO22X1 U6 ( .A0(shamt_i[0]), .A1(ExtOp_i), .B0(immed_i[0]), .B1(n20), .Y(
        ExtOut_o[0]) );
  AO22X1 U7 ( .A0(shamt_i[1]), .A1(ExtOp_i), .B0(immed_i[1]), .B1(n20), .Y(
        ExtOut_o[1]) );
  AO22X1 U8 ( .A0(shamt_i[2]), .A1(ExtOp_i), .B0(immed_i[2]), .B1(n20), .Y(
        ExtOut_o[2]) );
  AO22X1 U9 ( .A0(shamt_i[3]), .A1(ExtOp_i), .B0(immed_i[3]), .B1(n20), .Y(
        ExtOut_o[3]) );
  OAI2BB1X1 U10 ( .A0N(immed_i[4]), .A1N(n20), .B0(n19), .Y(ExtOut_o[4]) );
  OAI2BB1X1 U11 ( .A0N(immed_i[5]), .A1N(n20), .B0(n19), .Y(ExtOut_o[5]) );
  OAI2BB1X1 U12 ( .A0N(immed_i[6]), .A1N(n20), .B0(n19), .Y(ExtOut_o[6]) );
  OAI2BB1X1 U13 ( .A0N(immed_i[7]), .A1N(n20), .B0(n19), .Y(ExtOut_o[7]) );
  OAI2BB1X1 U14 ( .A0N(immed_i[8]), .A1N(n20), .B0(n19), .Y(ExtOut_o[8]) );
  OAI2BB1X1 U15 ( .A0N(immed_i[9]), .A1N(n20), .B0(n19), .Y(ExtOut_o[9]) );
  OAI2BB1X1 U16 ( .A0N(immed_i[10]), .A1N(n20), .B0(n19), .Y(ExtOut_o[10]) );
  OAI2BB1X1 U17 ( .A0N(immed_i[11]), .A1N(n20), .B0(n19), .Y(ExtOut_o[11]) );
  OAI2BB1X1 U18 ( .A0N(immed_i[12]), .A1N(n20), .B0(n19), .Y(ExtOut_o[12]) );
  OAI2BB1X1 U19 ( .A0N(immed_i[14]), .A1N(n20), .B0(n19), .Y(ExtOut_o[14]) );
  INVXL U20 ( .A(n1), .Y(ExtOut_o[16]) );
  INVXL U21 ( .A(n1), .Y(ExtOut_o[17]) );
  INVXL U22 ( .A(n1), .Y(ExtOut_o[18]) );
  INVXL U23 ( .A(n1), .Y(ExtOut_o[19]) );
  INVXL U24 ( .A(n1), .Y(ExtOut_o[20]) );
  INVXL U25 ( .A(n1), .Y(ExtOut_o[21]) );
  INVXL U26 ( .A(n1), .Y(ExtOut_o[22]) );
  INVXL U27 ( .A(n1), .Y(ExtOut_o[23]) );
  INVXL U28 ( .A(n1), .Y(ExtOut_o[24]) );
  INVXL U29 ( .A(n1), .Y(ExtOut_o[25]) );
  INVXL U30 ( .A(n1), .Y(ExtOut_o[26]) );
  INVXL U31 ( .A(n1), .Y(ExtOut_o[27]) );
  INVXL U32 ( .A(n1), .Y(ExtOut_o[28]) );
  INVXL U33 ( .A(n1), .Y(ExtOut_o[29]) );
  INVXL U34 ( .A(n1), .Y(ExtOut_o[31]) );
  CLKBUFX3 U35 ( .A(n2), .Y(n19) );
  NAND2X1 U36 ( .A(shamt_i[4]), .B(ExtOp_i), .Y(n2) );
endmodule


module MUX_5_3to1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [4:0] data0_i;
  input [4:0] data1_i;
  input [4:0] data2_i;
  input [1:0] select_i;
  output [4:0] data_o;
  wire   n6, n7, n8, n9, n10, n11, n12, n13;

  NOR2BX1 U2 ( .AN(select_i[1]), .B(select_i[0]), .Y(n8) );
  NOR2BX1 U3 ( .AN(select_i[0]), .B(select_i[1]), .Y(n9) );
  NOR2X1 U4 ( .A(select_i[0]), .B(select_i[1]), .Y(n7) );
  CLKINVX1 U5 ( .A(n13), .Y(data_o[0]) );
  AOI222XL U6 ( .A0(data0_i[0]), .A1(n7), .B0(data2_i[0]), .B1(n8), .C0(
        data1_i[0]), .C1(n9), .Y(n13) );
  CLKINVX1 U7 ( .A(n12), .Y(data_o[1]) );
  AOI222XL U8 ( .A0(data0_i[1]), .A1(n7), .B0(data2_i[1]), .B1(n8), .C0(
        data1_i[1]), .C1(n9), .Y(n12) );
  CLKINVX1 U9 ( .A(n11), .Y(data_o[2]) );
  AOI222XL U10 ( .A0(data0_i[2]), .A1(n7), .B0(data2_i[2]), .B1(n8), .C0(
        data1_i[2]), .C1(n9), .Y(n11) );
  CLKINVX1 U11 ( .A(n10), .Y(data_o[3]) );
  AOI222XL U12 ( .A0(data0_i[3]), .A1(n7), .B0(data2_i[3]), .B1(n8), .C0(
        data1_i[3]), .C1(n9), .Y(n10) );
  CLKINVX1 U13 ( .A(n6), .Y(data_o[4]) );
  AOI222XL U14 ( .A0(data0_i[4]), .A1(n7), .B0(data2_i[4]), .B1(n8), .C0(
        data1_i[4]), .C1(n9), .Y(n6) );
endmodule


module MUX_32_3to1_0 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53;

  NAND2X6 U2 ( .A(select_i[0]), .B(n18), .Y(n19) );
  INVX6 U3 ( .A(select_i[0]), .Y(n16) );
  CLKINVX16 U4 ( .A(n2), .Y(n8) );
  CLKINVX12 U5 ( .A(n3), .Y(n11) );
  AND2X6 U6 ( .A(n18), .B(n16), .Y(n1) );
  INVX20 U7 ( .A(n19), .Y(n51) );
  BUFX20 U8 ( .A(n52), .Y(n2) );
  BUFX16 U9 ( .A(n52), .Y(n3) );
  INVX6 U10 ( .A(n17), .Y(n4) );
  BUFX12 U11 ( .A(n4), .Y(n5) );
  BUFX12 U12 ( .A(n4), .Y(n6) );
  BUFX12 U13 ( .A(n4), .Y(n7) );
  INVX16 U14 ( .A(n8), .Y(n9) );
  INVX12 U15 ( .A(n8), .Y(n10) );
  INVX16 U16 ( .A(n11), .Y(n12) );
  INVX16 U17 ( .A(n11), .Y(n13) );
  INVX8 U18 ( .A(n17), .Y(n52) );
  NAND2X8 U19 ( .A(select_i[1]), .B(n16), .Y(n17) );
  BUFX20 U20 ( .A(n1), .Y(n14) );
  BUFX12 U21 ( .A(n1), .Y(n15) );
  INVX3 U22 ( .A(select_i[1]), .Y(n18) );
  AO22X4 U23 ( .A0(data2_i[2]), .A1(n12), .B0(data1_i[2]), .B1(n51), .Y(n22)
         );
  AO22X4 U24 ( .A0(data2_i[18]), .A1(n7), .B0(data1_i[18]), .B1(n51), .Y(n38)
         );
  AO22X4 U25 ( .A0(data2_i[0]), .A1(n10), .B0(data1_i[0]), .B1(n51), .Y(n20)
         );
  AO21X4 U26 ( .A0(data0_i[0]), .A1(n14), .B0(n20), .Y(data_o[0]) );
  AO22X4 U27 ( .A0(data2_i[1]), .A1(n9), .B0(data1_i[1]), .B1(n51), .Y(n21) );
  AO21X4 U28 ( .A0(data0_i[1]), .A1(n14), .B0(n21), .Y(data_o[1]) );
  AO21X4 U29 ( .A0(data0_i[2]), .A1(n14), .B0(n22), .Y(data_o[2]) );
  AO22X4 U30 ( .A0(data2_i[3]), .A1(n5), .B0(data1_i[3]), .B1(n51), .Y(n23) );
  AO21X4 U31 ( .A0(data0_i[3]), .A1(n15), .B0(n23), .Y(data_o[3]) );
  AO22X4 U32 ( .A0(data2_i[4]), .A1(n13), .B0(data1_i[4]), .B1(n51), .Y(n24)
         );
  AO21X4 U33 ( .A0(data0_i[4]), .A1(n14), .B0(n24), .Y(data_o[4]) );
  AO22X4 U34 ( .A0(data2_i[5]), .A1(n12), .B0(data1_i[5]), .B1(n51), .Y(n25)
         );
  AO21X4 U35 ( .A0(data0_i[5]), .A1(n15), .B0(n25), .Y(data_o[5]) );
  AO22X4 U36 ( .A0(data2_i[6]), .A1(n9), .B0(data1_i[6]), .B1(n51), .Y(n26) );
  AO21X4 U37 ( .A0(data0_i[6]), .A1(n15), .B0(n26), .Y(data_o[6]) );
  AO22X4 U38 ( .A0(data2_i[7]), .A1(n13), .B0(data1_i[7]), .B1(n51), .Y(n27)
         );
  AO21X4 U39 ( .A0(data0_i[7]), .A1(n14), .B0(n27), .Y(data_o[7]) );
  AO22X4 U40 ( .A0(data2_i[8]), .A1(n10), .B0(data1_i[8]), .B1(n51), .Y(n28)
         );
  AO21X4 U41 ( .A0(data0_i[8]), .A1(n14), .B0(n28), .Y(data_o[8]) );
  AO22X4 U42 ( .A0(data2_i[9]), .A1(n13), .B0(data1_i[9]), .B1(n51), .Y(n29)
         );
  AO21X4 U43 ( .A0(data0_i[9]), .A1(n14), .B0(n29), .Y(data_o[9]) );
  AO22X4 U44 ( .A0(data2_i[10]), .A1(n12), .B0(data1_i[10]), .B1(n51), .Y(n30)
         );
  AO21X4 U45 ( .A0(data0_i[10]), .A1(n14), .B0(n30), .Y(data_o[10]) );
  AO22X4 U46 ( .A0(data2_i[11]), .A1(n7), .B0(data1_i[11]), .B1(n51), .Y(n31)
         );
  AO21X4 U47 ( .A0(data0_i[11]), .A1(n15), .B0(n31), .Y(data_o[11]) );
  AO22X4 U48 ( .A0(data2_i[12]), .A1(n5), .B0(data1_i[12]), .B1(n51), .Y(n32)
         );
  AO21X4 U49 ( .A0(data0_i[12]), .A1(n14), .B0(n32), .Y(data_o[12]) );
  AO22X4 U50 ( .A0(data2_i[13]), .A1(n9), .B0(data1_i[13]), .B1(n51), .Y(n33)
         );
  AO21X4 U51 ( .A0(data0_i[13]), .A1(n14), .B0(n33), .Y(data_o[13]) );
  AO22X4 U52 ( .A0(data2_i[14]), .A1(n9), .B0(data1_i[14]), .B1(n51), .Y(n34)
         );
  AO21X4 U53 ( .A0(data0_i[14]), .A1(n14), .B0(n34), .Y(data_o[14]) );
  AO22X4 U54 ( .A0(data2_i[15]), .A1(n6), .B0(data1_i[15]), .B1(n51), .Y(n35)
         );
  AO21X4 U55 ( .A0(data0_i[15]), .A1(n14), .B0(n35), .Y(data_o[15]) );
  AO22X4 U56 ( .A0(data2_i[16]), .A1(n13), .B0(data1_i[16]), .B1(n51), .Y(n36)
         );
  AO21X4 U57 ( .A0(data0_i[16]), .A1(n14), .B0(n36), .Y(data_o[16]) );
  AO22X4 U58 ( .A0(data2_i[17]), .A1(n6), .B0(data1_i[17]), .B1(n51), .Y(n37)
         );
  AO21X4 U59 ( .A0(data0_i[17]), .A1(n14), .B0(n37), .Y(data_o[17]) );
  AO21X4 U60 ( .A0(data0_i[18]), .A1(n15), .B0(n38), .Y(data_o[18]) );
  AO22X4 U61 ( .A0(data2_i[19]), .A1(n6), .B0(data1_i[19]), .B1(n51), .Y(n39)
         );
  AO21X4 U62 ( .A0(data0_i[19]), .A1(n15), .B0(n39), .Y(data_o[19]) );
  AO22X4 U63 ( .A0(data2_i[20]), .A1(n5), .B0(data1_i[20]), .B1(n51), .Y(n40)
         );
  AO21X4 U64 ( .A0(data0_i[20]), .A1(n14), .B0(n40), .Y(data_o[20]) );
  AO22X4 U65 ( .A0(data2_i[21]), .A1(n6), .B0(data1_i[21]), .B1(n51), .Y(n41)
         );
  AO21X4 U66 ( .A0(data0_i[21]), .A1(n14), .B0(n41), .Y(data_o[21]) );
  AO22X4 U67 ( .A0(data2_i[22]), .A1(n5), .B0(data1_i[22]), .B1(n51), .Y(n42)
         );
  AO21X4 U68 ( .A0(data0_i[22]), .A1(n15), .B0(n42), .Y(data_o[22]) );
  AO22X4 U69 ( .A0(data2_i[23]), .A1(n7), .B0(data1_i[23]), .B1(n51), .Y(n43)
         );
  AO21X4 U70 ( .A0(data0_i[23]), .A1(n14), .B0(n43), .Y(data_o[23]) );
  AO22X4 U71 ( .A0(data2_i[24]), .A1(n7), .B0(data1_i[24]), .B1(n51), .Y(n44)
         );
  AO21X4 U72 ( .A0(data0_i[24]), .A1(n15), .B0(n44), .Y(data_o[24]) );
  AO22X4 U73 ( .A0(data2_i[25]), .A1(n5), .B0(data1_i[25]), .B1(n51), .Y(n45)
         );
  AO21X4 U74 ( .A0(data0_i[25]), .A1(n15), .B0(n45), .Y(data_o[25]) );
  AO22X4 U75 ( .A0(data2_i[26]), .A1(n12), .B0(data1_i[26]), .B1(n51), .Y(n46)
         );
  AO21X4 U76 ( .A0(data0_i[26]), .A1(n14), .B0(n46), .Y(data_o[26]) );
  AO22X4 U77 ( .A0(data2_i[27]), .A1(n6), .B0(data1_i[27]), .B1(n51), .Y(n47)
         );
  AO21X4 U78 ( .A0(data0_i[27]), .A1(n14), .B0(n47), .Y(data_o[27]) );
  AO22X4 U79 ( .A0(data2_i[28]), .A1(n7), .B0(data1_i[28]), .B1(n51), .Y(n48)
         );
  AO21X4 U80 ( .A0(data0_i[28]), .A1(n15), .B0(n48), .Y(data_o[28]) );
  AO22X4 U81 ( .A0(data2_i[29]), .A1(n9), .B0(data1_i[29]), .B1(n51), .Y(n49)
         );
  AO21X4 U82 ( .A0(data0_i[29]), .A1(n15), .B0(n49), .Y(data_o[29]) );
  AO22X4 U83 ( .A0(data2_i[30]), .A1(n10), .B0(data1_i[30]), .B1(n51), .Y(n50)
         );
  AO21X4 U84 ( .A0(data0_i[30]), .A1(n14), .B0(n50), .Y(data_o[30]) );
  AO22X4 U85 ( .A0(data2_i[31]), .A1(n10), .B0(data1_i[31]), .B1(n51), .Y(n53)
         );
  AO21X4 U86 ( .A0(data0_i[31]), .A1(n14), .B0(n53), .Y(data_o[31]) );
endmodule


module MUX_32_3to1_2 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n59, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58;

  BUFX8 U2 ( .A(n35), .Y(n42) );
  AOI22X2 U3 ( .A0(data0_i[3]), .A1(n27), .B0(data1_i[3]), .B1(n20), .Y(n33)
         );
  OAI2BB1X4 U4 ( .A0N(data2_i[16]), .A1N(n42), .B0(n1), .Y(data_o[16]) );
  AOI22X2 U5 ( .A0(data0_i[16]), .A1(n26), .B0(data1_i[16]), .B1(n20), .Y(n1)
         );
  INVX20 U6 ( .A(n25), .Y(n27) );
  INVX20 U7 ( .A(n25), .Y(n28) );
  CLKINVX16 U8 ( .A(n40), .Y(n25) );
  INVX16 U9 ( .A(n38), .Y(n18) );
  INVX16 U10 ( .A(n29), .Y(data_o[31]) );
  INVX2 U11 ( .A(data2_i[4]), .Y(n13) );
  CLKINVX6 U12 ( .A(data2_i[31]), .Y(n30) );
  CLKINVX6 U13 ( .A(data2_i[13]), .Y(n17) );
  BUFX20 U14 ( .A(n35), .Y(n41) );
  OAI21X4 U15 ( .A0(n31), .A1(n13), .B0(n9), .Y(data_o[4]) );
  AOI22X4 U16 ( .A0(data0_i[28]), .A1(n28), .B0(data1_i[28]), .B1(n20), .Y(n12) );
  OAI2BB1X4 U17 ( .A0N(data2_i[29]), .A1N(n42), .B0(n3), .Y(data_o[29]) );
  AOI22X2 U18 ( .A0(n27), .A1(data0_i[29]), .B0(data1_i[29]), .B1(n20), .Y(n3)
         );
  AOI22X2 U19 ( .A0(data0_i[4]), .A1(n27), .B0(data1_i[4]), .B1(n20), .Y(n9)
         );
  INVX20 U20 ( .A(n25), .Y(n26) );
  OAI2BB1X4 U21 ( .A0N(data2_i[17]), .A1N(n42), .B0(n4), .Y(data_o[17]) );
  AOI22X2 U22 ( .A0(data0_i[17]), .A1(n27), .B0(data1_i[17]), .B1(n20), .Y(n4)
         );
  CLKINVX12 U23 ( .A(n18), .Y(n19) );
  OAI2BB1X4 U24 ( .A0N(data2_i[25]), .A1N(n42), .B0(n5), .Y(data_o[25]) );
  AOI22X2 U25 ( .A0(data0_i[25]), .A1(n27), .B0(data1_i[25]), .B1(n20), .Y(n5)
         );
  AOI22X2 U26 ( .A0(n19), .A1(data1_i[0]), .B0(data0_i[0]), .B1(n26), .Y(n15)
         );
  OAI2BB1X4 U27 ( .A0N(data2_i[2]), .A1N(n41), .B0(n10), .Y(n6) );
  INVX16 U28 ( .A(n41), .Y(n31) );
  AOI22X4 U29 ( .A0(data0_i[27]), .A1(n28), .B0(data1_i[27]), .B1(n19), .Y(n11) );
  INVX8 U30 ( .A(n6), .Y(n23) );
  CLKINVX12 U31 ( .A(n44), .Y(n39) );
  OA21X4 U32 ( .A0(n30), .A1(n31), .B0(n7), .Y(n29) );
  AOI22X4 U33 ( .A0(data0_i[31]), .A1(n27), .B0(data1_i[31]), .B1(n20), .Y(n7)
         );
  AOI22X4 U34 ( .A0(n27), .A1(data0_i[7]), .B0(data1_i[7]), .B1(n19), .Y(n32)
         );
  AOI22X4 U35 ( .A0(data0_i[24]), .A1(n28), .B0(data1_i[24]), .B1(n20), .Y(n22) );
  INVX4 U36 ( .A(n16), .Y(data_o[13]) );
  INVX20 U37 ( .A(n23), .Y(data_o[2]) );
  AO21X4 U38 ( .A0(data2_i[12]), .A1(n41), .B0(n49), .Y(data_o[12]) );
  OAI2BB1X4 U39 ( .A0N(data2_i[6]), .A1N(n41), .B0(n8), .Y(data_o[6]) );
  AOI22X2 U40 ( .A0(n28), .A1(data0_i[6]), .B0(data1_i[6]), .B1(n19), .Y(n8)
         );
  AND2X4 U41 ( .A(n43), .B(n39), .Y(n35) );
  CLKAND2X12 U42 ( .A(n43), .B(n44), .Y(n40) );
  AOI22X4 U43 ( .A0(data0_i[2]), .A1(n28), .B0(data1_i[2]), .B1(n20), .Y(n10)
         );
  AOI22X4 U44 ( .A0(data0_i[21]), .A1(n28), .B0(data1_i[21]), .B1(n20), .Y(n37) );
  OAI2BB1X4 U45 ( .A0N(data2_i[27]), .A1N(n41), .B0(n11), .Y(n59) );
  OAI2BB1X4 U46 ( .A0N(data2_i[28]), .A1N(n41), .B0(n12), .Y(data_o[28]) );
  OAI2BB1X4 U47 ( .A0N(data2_i[26]), .A1N(n42), .B0(n14), .Y(data_o[26]) );
  AOI22X2 U48 ( .A0(data0_i[26]), .A1(n28), .B0(data1_i[26]), .B1(n20), .Y(n14) );
  OAI2BB1X4 U49 ( .A0N(data2_i[0]), .A1N(n41), .B0(n15), .Y(data_o[0]) );
  CLKINVX20 U50 ( .A(n18), .Y(n20) );
  AO21X4 U51 ( .A0(data2_i[9]), .A1(n41), .B0(n47), .Y(data_o[9]) );
  INVX4 U52 ( .A(select_i[0]), .Y(n43) );
  AOI2BB1X4 U53 ( .A0N(n17), .A1N(n31), .B0(n50), .Y(n16) );
  NOR2X6 U54 ( .A(n43), .B(n39), .Y(n38) );
  OAI2BB1X4 U55 ( .A0N(data2_i[11]), .A1N(n41), .B0(n21), .Y(data_o[11]) );
  AOI22X2 U56 ( .A0(data0_i[11]), .A1(n28), .B0(data1_i[11]), .B1(n19), .Y(n21) );
  OAI2BB1X4 U57 ( .A0N(data2_i[24]), .A1N(n41), .B0(n22), .Y(data_o[24]) );
  OAI2BB1X4 U58 ( .A0N(data2_i[5]), .A1N(n41), .B0(n24), .Y(data_o[5]) );
  AOI22X2 U59 ( .A0(data0_i[5]), .A1(n27), .B0(data1_i[5]), .B1(n19), .Y(n24)
         );
  AO21X4 U60 ( .A0(data2_i[23]), .A1(n42), .B0(n57), .Y(data_o[23]) );
  OAI2BB1X4 U61 ( .A0N(data2_i[21]), .A1N(n41), .B0(n37), .Y(data_o[21]) );
  OAI2BB1X4 U62 ( .A0N(data2_i[7]), .A1N(n41), .B0(n32), .Y(data_o[7]) );
  OAI2BB1X4 U63 ( .A0N(data2_i[3]), .A1N(n41), .B0(n33), .Y(data_o[3]) );
  AO21X4 U64 ( .A0(data2_i[8]), .A1(n41), .B0(n46), .Y(data_o[8]) );
  BUFX20 U65 ( .A(n59), .Y(data_o[27]) );
  INVX8 U66 ( .A(select_i[1]), .Y(n44) );
  AO21X4 U67 ( .A0(data2_i[1]), .A1(n42), .B0(n45), .Y(data_o[1]) );
  AO21X4 U68 ( .A0(data2_i[20]), .A1(n42), .B0(n55), .Y(data_o[20]) );
  AO21X4 U69 ( .A0(data2_i[18]), .A1(n42), .B0(n53), .Y(data_o[18]) );
  AO22X4 U70 ( .A0(data0_i[1]), .A1(n26), .B0(data1_i[1]), .B1(n20), .Y(n45)
         );
  AO22X4 U71 ( .A0(data0_i[8]), .A1(n26), .B0(data1_i[8]), .B1(n20), .Y(n46)
         );
  AO22X4 U72 ( .A0(data0_i[9]), .A1(n26), .B0(data1_i[9]), .B1(n20), .Y(n47)
         );
  AO22X4 U73 ( .A0(data0_i[10]), .A1(n26), .B0(data1_i[10]), .B1(n20), .Y(n48)
         );
  AO21X4 U74 ( .A0(data2_i[10]), .A1(n41), .B0(n48), .Y(data_o[10]) );
  AO22X4 U75 ( .A0(data0_i[12]), .A1(n27), .B0(data1_i[12]), .B1(n19), .Y(n49)
         );
  AO22X4 U76 ( .A0(data0_i[13]), .A1(n26), .B0(data1_i[13]), .B1(n19), .Y(n50)
         );
  AO22X4 U77 ( .A0(n28), .A1(data0_i[14]), .B0(n19), .B1(data1_i[14]), .Y(n51)
         );
  AO21X4 U78 ( .A0(n42), .A1(data2_i[14]), .B0(n51), .Y(data_o[14]) );
  AO22X4 U79 ( .A0(data0_i[15]), .A1(n26), .B0(data1_i[15]), .B1(n19), .Y(n52)
         );
  AO21X4 U80 ( .A0(data2_i[15]), .A1(n42), .B0(n52), .Y(data_o[15]) );
  AO22X4 U81 ( .A0(data0_i[18]), .A1(n28), .B0(data1_i[18]), .B1(n19), .Y(n53)
         );
  AO22X4 U82 ( .A0(data0_i[19]), .A1(n26), .B0(n19), .B1(data1_i[19]), .Y(n54)
         );
  AO21X4 U83 ( .A0(data2_i[19]), .A1(n42), .B0(n54), .Y(data_o[19]) );
  AO22X4 U84 ( .A0(data0_i[20]), .A1(n26), .B0(data1_i[20]), .B1(n20), .Y(n55)
         );
  AO22X4 U85 ( .A0(data0_i[22]), .A1(n26), .B0(data1_i[22]), .B1(n20), .Y(n56)
         );
  AO21X4 U86 ( .A0(data2_i[22]), .A1(n42), .B0(n56), .Y(data_o[22]) );
  AO22X4 U87 ( .A0(data0_i[23]), .A1(n26), .B0(data1_i[23]), .B1(n19), .Y(n57)
         );
  AO22X4 U88 ( .A0(n27), .A1(data0_i[30]), .B0(data1_i[30]), .B1(n20), .Y(n58)
         );
  AO21X4 U89 ( .A0(data2_i[30]), .A1(n42), .B0(n58), .Y(data_o[30]) );
endmodule


module MUX_32_3to1_1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  AOI22X4 U2 ( .A0(data2_i[28]), .A1(n14), .B0(data1_i[28]), .B1(n2), .Y(n9)
         );
  BUFX16 U3 ( .A(n48), .Y(n14) );
  BUFX20 U4 ( .A(n5), .Y(n17) );
  INVX20 U5 ( .A(n11), .Y(n1) );
  INVX16 U6 ( .A(n1), .Y(n2) );
  INVX16 U7 ( .A(n1), .Y(n3) );
  INVX12 U8 ( .A(n1), .Y(n4) );
  INVX2 U9 ( .A(select_i[1]), .Y(n20) );
  AND2X8 U10 ( .A(n18), .B(n20), .Y(n5) );
  AOI22X4 U11 ( .A0(data2_i[6]), .A1(n13), .B0(data1_i[6]), .B1(n3), .Y(n6) );
  NAND2X6 U12 ( .A(n18), .B(select_i[1]), .Y(n19) );
  INVX12 U13 ( .A(select_i[0]), .Y(n18) );
  INVX12 U14 ( .A(n19), .Y(n48) );
  AOI22X4 U15 ( .A0(data2_i[10]), .A1(n13), .B0(data1_i[10]), .B1(n3), .Y(n8)
         );
  NOR2X8 U16 ( .A(n18), .B(select_i[1]), .Y(n11) );
  OAI2BB1X4 U17 ( .A0N(data0_i[6]), .A1N(n5), .B0(n6), .Y(data_o[6]) );
  AOI22X2 U18 ( .A0(data2_i[2]), .A1(n14), .B0(data1_i[2]), .B1(n4), .Y(n10)
         );
  OAI2BB1X4 U19 ( .A0N(data0_i[31]), .A1N(n17), .B0(n7), .Y(data_o[31]) );
  AOI22X2 U20 ( .A0(data2_i[31]), .A1(n15), .B0(data1_i[31]), .B1(n4), .Y(n7)
         );
  OR2X8 U21 ( .A(n24), .B(n12), .Y(data_o[4]) );
  AO22X4 U22 ( .A0(data2_i[8]), .A1(n13), .B0(data1_i[8]), .B1(n2), .Y(n27) );
  AO22X4 U23 ( .A0(data2_i[5]), .A1(n13), .B0(data1_i[5]), .B1(n3), .Y(n25) );
  OAI2BB1X4 U24 ( .A0N(data0_i[10]), .A1N(n16), .B0(n8), .Y(data_o[10]) );
  AO22X4 U25 ( .A0(data2_i[30]), .A1(n13), .B0(data1_i[30]), .B1(n2), .Y(n47)
         );
  AO22X4 U26 ( .A0(data2_i[9]), .A1(n15), .B0(data1_i[9]), .B1(n4), .Y(n28) );
  AO22X4 U27 ( .A0(data2_i[29]), .A1(n13), .B0(data1_i[29]), .B1(n3), .Y(n46)
         );
  OAI2BB1X4 U28 ( .A0N(data0_i[28]), .A1N(n17), .B0(n9), .Y(data_o[28]) );
  OAI2BB1X4 U29 ( .A0N(data0_i[2]), .A1N(n16), .B0(n10), .Y(data_o[2]) );
  AO22X4 U30 ( .A0(data2_i[7]), .A1(n14), .B0(data1_i[7]), .B1(n3), .Y(n26) );
  AO22X4 U31 ( .A0(data2_i[1]), .A1(n15), .B0(data1_i[1]), .B1(n2), .Y(n22) );
  AO22X2 U32 ( .A0(data2_i[4]), .A1(n15), .B0(data1_i[4]), .B1(n2), .Y(n24) );
  AO22X4 U33 ( .A0(data2_i[11]), .A1(n13), .B0(data1_i[11]), .B1(n2), .Y(n29)
         );
  AND2X1 U34 ( .A(data0_i[4]), .B(n16), .Y(n12) );
  BUFX20 U35 ( .A(n5), .Y(n16) );
  AO22X4 U36 ( .A0(data2_i[16]), .A1(n14), .B0(data1_i[16]), .B1(n4), .Y(n34)
         );
  AO22X4 U37 ( .A0(data2_i[17]), .A1(n13), .B0(data1_i[17]), .B1(n4), .Y(n35)
         );
  AO22X4 U38 ( .A0(data2_i[20]), .A1(n14), .B0(data1_i[20]), .B1(n4), .Y(n38)
         );
  AO22X4 U39 ( .A0(data2_i[15]), .A1(n15), .B0(data1_i[15]), .B1(n4), .Y(n33)
         );
  AO22X4 U40 ( .A0(data2_i[23]), .A1(n15), .B0(data1_i[23]), .B1(n4), .Y(n41)
         );
  AO22X4 U41 ( .A0(data2_i[0]), .A1(n13), .B0(data1_i[0]), .B1(n2), .Y(n21) );
  AO21X4 U42 ( .A0(data0_i[0]), .A1(n16), .B0(n21), .Y(data_o[0]) );
  AO22X4 U43 ( .A0(data2_i[21]), .A1(n14), .B0(data1_i[21]), .B1(n3), .Y(n39)
         );
  AO22X4 U44 ( .A0(data2_i[19]), .A1(n14), .B0(data1_i[19]), .B1(n3), .Y(n37)
         );
  AO22X4 U45 ( .A0(data2_i[13]), .A1(n15), .B0(data1_i[13]), .B1(n2), .Y(n31)
         );
  AO22X4 U46 ( .A0(data2_i[18]), .A1(n15), .B0(data1_i[18]), .B1(n2), .Y(n36)
         );
  AO22X4 U47 ( .A0(data2_i[26]), .A1(n13), .B0(data1_i[26]), .B1(n3), .Y(n44)
         );
  AO22X4 U48 ( .A0(data2_i[24]), .A1(n15), .B0(data1_i[24]), .B1(n3), .Y(n42)
         );
  BUFX20 U49 ( .A(n48), .Y(n15) );
  BUFX20 U50 ( .A(n48), .Y(n13) );
  AO21X4 U51 ( .A0(data0_i[1]), .A1(n16), .B0(n22), .Y(data_o[1]) );
  AO22X4 U52 ( .A0(data2_i[3]), .A1(n13), .B0(data1_i[3]), .B1(n4), .Y(n23) );
  AO21X4 U53 ( .A0(data0_i[3]), .A1(n16), .B0(n23), .Y(data_o[3]) );
  AO21X4 U54 ( .A0(data0_i[5]), .A1(n16), .B0(n25), .Y(data_o[5]) );
  AO21X4 U55 ( .A0(data0_i[7]), .A1(n16), .B0(n26), .Y(data_o[7]) );
  AO21X4 U56 ( .A0(data0_i[8]), .A1(n16), .B0(n27), .Y(data_o[8]) );
  AO21X4 U57 ( .A0(data0_i[9]), .A1(n16), .B0(n28), .Y(data_o[9]) );
  AO21X4 U58 ( .A0(data0_i[11]), .A1(n16), .B0(n29), .Y(data_o[11]) );
  AO22X4 U59 ( .A0(data2_i[12]), .A1(n15), .B0(data1_i[12]), .B1(n4), .Y(n30)
         );
  AO21X4 U60 ( .A0(data0_i[12]), .A1(n16), .B0(n30), .Y(data_o[12]) );
  AO21X4 U61 ( .A0(data0_i[13]), .A1(n17), .B0(n31), .Y(data_o[13]) );
  AO22X4 U62 ( .A0(data2_i[14]), .A1(n15), .B0(data1_i[14]), .B1(n2), .Y(n32)
         );
  AO21X4 U63 ( .A0(data0_i[14]), .A1(n17), .B0(n32), .Y(data_o[14]) );
  AO21X4 U64 ( .A0(data0_i[15]), .A1(n17), .B0(n33), .Y(data_o[15]) );
  AO21X4 U65 ( .A0(data0_i[16]), .A1(n17), .B0(n34), .Y(data_o[16]) );
  AO21X4 U66 ( .A0(data0_i[17]), .A1(n17), .B0(n35), .Y(data_o[17]) );
  AO21X4 U67 ( .A0(data0_i[18]), .A1(n17), .B0(n36), .Y(data_o[18]) );
  AO21X4 U68 ( .A0(data0_i[19]), .A1(n17), .B0(n37), .Y(data_o[19]) );
  AO21X4 U69 ( .A0(data0_i[20]), .A1(n17), .B0(n38), .Y(data_o[20]) );
  AO21X4 U70 ( .A0(data0_i[21]), .A1(n17), .B0(n39), .Y(data_o[21]) );
  AO22X4 U71 ( .A0(data2_i[22]), .A1(n15), .B0(data1_i[22]), .B1(n2), .Y(n40)
         );
  AO21X4 U72 ( .A0(data0_i[22]), .A1(n17), .B0(n40), .Y(data_o[22]) );
  AO21X4 U73 ( .A0(data0_i[23]), .A1(n17), .B0(n41), .Y(data_o[23]) );
  AO21X4 U74 ( .A0(data0_i[24]), .A1(n17), .B0(n42), .Y(data_o[24]) );
  AO22X4 U75 ( .A0(data2_i[25]), .A1(n15), .B0(data1_i[25]), .B1(n3), .Y(n43)
         );
  AO21X4 U76 ( .A0(data0_i[25]), .A1(n17), .B0(n43), .Y(data_o[25]) );
  AO21X4 U77 ( .A0(data0_i[26]), .A1(n17), .B0(n44), .Y(data_o[26]) );
  AO22X4 U78 ( .A0(data2_i[27]), .A1(n13), .B0(data1_i[27]), .B1(n3), .Y(n45)
         );
  AO21X4 U79 ( .A0(data0_i[27]), .A1(n17), .B0(n45), .Y(data_o[27]) );
  AO21X4 U80 ( .A0(data0_i[29]), .A1(n17), .B0(n46), .Y(data_o[29]) );
  AO21X4 U81 ( .A0(data0_i[30]), .A1(n17), .B0(n47), .Y(data_o[30]) );
endmodule


module forwarding ( Rs_regD, Rt_regD, RegWrite_regE, wsel_regE, RegWrite_regM, 
        wsel_regM, FU_Asel, FU_Bsel );
  input [4:0] Rs_regD;
  input [4:0] Rt_regD;
  input [4:0] wsel_regE;
  input [4:0] wsel_regM;
  output [1:0] FU_Asel;
  output [1:0] FU_Bsel;
  input RegWrite_regE, RegWrite_regM;
  wire   n55, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;

  NOR2X8 U2 ( .A(n15), .B(n16), .Y(n20) );
  NAND2X4 U3 ( .A(n45), .B(n43), .Y(n50) );
  INVX8 U4 ( .A(wsel_regE[1]), .Y(n35) );
  INVX6 U5 ( .A(wsel_regE[4]), .Y(n36) );
  INVX8 U6 ( .A(wsel_regM[1]), .Y(n45) );
  XNOR2X2 U7 ( .A(wsel_regM[1]), .B(Rs_regD[1]), .Y(n48) );
  INVX12 U8 ( .A(wsel_regE[0]), .Y(n32) );
  NOR2X6 U9 ( .A(n24), .B(n23), .Y(n55) );
  NAND2X4 U10 ( .A(n28), .B(n29), .Y(n30) );
  INVX12 U11 ( .A(wsel_regM[0]), .Y(n46) );
  INVX12 U12 ( .A(wsel_regM[2]), .Y(n43) );
  XNOR2X4 U13 ( .A(Rt_regD[4]), .B(wsel_regM[4]), .Y(n26) );
  INVX12 U14 ( .A(wsel_regM[4]), .Y(n39) );
  NOR2X6 U15 ( .A(n24), .B(n23), .Y(FU_Bsel[1]) );
  CLKAND2X4 U16 ( .A(n8), .B(n53), .Y(FU_Asel[1]) );
  NAND2X8 U17 ( .A(n33), .B(RegWrite_regE), .Y(n3) );
  NAND4X4 U18 ( .A(n6), .B(RegWrite_regM), .C(n27), .D(n26), .Y(n31) );
  INVX12 U19 ( .A(wsel_regM[3]), .Y(n44) );
  INVX12 U20 ( .A(wsel_regE[3]), .Y(n17) );
  XNOR2X4 U21 ( .A(wsel_regM[0]), .B(Rs_regD[0]), .Y(n47) );
  XNOR2X4 U22 ( .A(wsel_regE[2]), .B(Rs_regD[2]), .Y(n11) );
  INVX12 U23 ( .A(wsel_regE[2]), .Y(n34) );
  NOR2X6 U24 ( .A(wsel_regE[0]), .B(wsel_regE[3]), .Y(n37) );
  CLKAND2X12 U25 ( .A(RegWrite_regM), .B(n40), .Y(n12) );
  NOR2X8 U26 ( .A(n14), .B(n13), .Y(n21) );
  XOR2X4 U27 ( .A(wsel_regE[4]), .B(Rt_regD[4]), .Y(n13) );
  OR3X8 U28 ( .A(wsel_regM[4]), .B(wsel_regM[3]), .C(n5), .Y(n27) );
  NAND3X6 U29 ( .A(n45), .B(n46), .C(n43), .Y(n5) );
  NAND4X4 U30 ( .A(n37), .B(n36), .C(n34), .D(n35), .Y(n38) );
  NOR2X4 U31 ( .A(wsel_regE[2]), .B(wsel_regE[1]), .Y(n18) );
  NAND3X6 U32 ( .A(n46), .B(n44), .C(n39), .Y(n49) );
  NOR3X8 U33 ( .A(n2), .B(n3), .C(n1), .Y(n8) );
  XNOR2X4 U34 ( .A(n32), .B(Rs_regD[0]), .Y(n1) );
  XNOR2X4 U35 ( .A(n35), .B(Rs_regD[1]), .Y(n2) );
  XNOR2X4 U36 ( .A(n34), .B(Rt_regD[2]), .Y(n14) );
  XNOR2X2 U37 ( .A(n46), .B(Rt_regD[0]), .Y(n4) );
  NAND3X6 U38 ( .A(n19), .B(n20), .C(n21), .Y(n24) );
  NAND2X8 U39 ( .A(n22), .B(RegWrite_regE), .Y(n23) );
  XOR2X4 U40 ( .A(n32), .B(Rt_regD[0]), .Y(n22) );
  XNOR2X4 U41 ( .A(wsel_regE[4]), .B(Rs_regD[4]), .Y(n33) );
  CLKINVX2 U42 ( .A(Rt_regD[3]), .Y(n25) );
  XOR2X4 U43 ( .A(n25), .B(wsel_regM[3]), .Y(n6) );
  XOR2X4 U44 ( .A(n17), .B(Rs_regD[3]), .Y(n10) );
  XNOR2X2 U45 ( .A(wsel_regM[2]), .B(Rt_regD[2]), .Y(n29) );
  XNOR2X4 U46 ( .A(wsel_regM[1]), .B(Rt_regD[1]), .Y(n28) );
  XNOR2X4 U47 ( .A(wsel_regM[2]), .B(Rs_regD[2]), .Y(n40) );
  NAND4X2 U48 ( .A(n18), .B(n32), .C(n17), .D(n36), .Y(n19) );
  AND2X8 U49 ( .A(n41), .B(n42), .Y(n9) );
  AND3X8 U50 ( .A(n38), .B(n10), .C(n11), .Y(n53) );
  XOR2X4 U51 ( .A(n39), .B(Rs_regD[4]), .Y(n41) );
  XOR2X4 U52 ( .A(n44), .B(Rs_regD[3]), .Y(n42) );
  NAND2X6 U53 ( .A(n9), .B(n12), .Y(n52) );
  XOR2X4 U54 ( .A(Rt_regD[1]), .B(wsel_regE[1]), .Y(n15) );
  NOR4X8 U55 ( .A(n55), .B(n31), .C(n4), .D(n30), .Y(FU_Bsel[0]) );
  XOR2X4 U56 ( .A(wsel_regE[3]), .B(Rt_regD[3]), .Y(n16) );
  OAI211X2 U57 ( .A0(n49), .A1(n50), .B0(n47), .C0(n48), .Y(n51) );
  AOI211X2 U58 ( .A0(n53), .A1(n8), .B0(n52), .C0(n51), .Y(FU_Asel[0]) );
endmodule


module hazard_detection ( Branch_EX, equal, branchpred_his, JumpReg_regD, 
        MemRead_regD, Rt_regD, Rs, Rt, ICACHE_stall, DCACHE_stall, 
        stall_lw_use, stallcache, flush, pred_cond );
  input [4:0] Rt_regD;
  input [4:0] Rs;
  input [4:0] Rt;
  input Branch_EX, equal, branchpred_his, JumpReg_regD, MemRead_regD,
         ICACHE_stall, DCACHE_stall;
  output stall_lw_use, stallcache, flush, pred_cond;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;

  INVXL U2 ( .A(pred_cond), .Y(n1) );
  INVX12 U3 ( .A(n19), .Y(pred_cond) );
  INVX4 U4 ( .A(Rt_regD[2]), .Y(n7) );
  CLKINVX8 U5 ( .A(n2), .Y(stall_lw_use) );
  OR2X8 U6 ( .A(n20), .B(JumpReg_regD), .Y(n2) );
  XOR2XL U7 ( .A(Rt[1]), .B(Rt_regD[1]), .Y(n13) );
  XOR2XL U8 ( .A(Rt[4]), .B(Rt_regD[4]), .Y(n12) );
  XOR2XL U9 ( .A(Rs[1]), .B(Rt_regD[1]), .Y(n16) );
  XOR2XL U10 ( .A(Rs[4]), .B(Rt_regD[4]), .Y(n15) );
  XOR2X1 U11 ( .A(n8), .B(Rt[3]), .Y(n9) );
  XOR2X1 U12 ( .A(n7), .B(Rt[2]), .Y(n10) );
  XOR2XL U13 ( .A(Rt[0]), .B(Rt_regD[0]), .Y(n11) );
  XOR2X1 U14 ( .A(n8), .B(Rs[3]), .Y(n4) );
  XOR2X1 U15 ( .A(n7), .B(Rs[2]), .Y(n5) );
  XOR2XL U16 ( .A(Rs[0]), .B(Rt_regD[0]), .Y(n6) );
  INVXL U17 ( .A(Rt_regD[3]), .Y(n8) );
  OR2X8 U18 ( .A(ICACHE_stall), .B(DCACHE_stall), .Y(stallcache) );
  NAND3BXL U19 ( .AN(JumpReg_regD), .B(n1), .C(n20), .Y(flush) );
  NAND2X8 U20 ( .A(n3), .B(Branch_EX), .Y(n19) );
  XOR2X4 U21 ( .A(equal), .B(branchpred_his), .Y(n3) );
  NAND3BX2 U22 ( .AN(n6), .B(n5), .C(n4), .Y(n17) );
  NAND3BX2 U23 ( .AN(n11), .B(n10), .C(n9), .Y(n14) );
  OAI33X2 U24 ( .A0(n17), .A1(n16), .A2(n15), .B0(n14), .B1(n13), .B2(n12), 
        .Y(n18) );
  NAND2X2 U25 ( .A(MemRead_regD), .B(n18), .Y(n20) );
endmodule


module branch_prediction ( clk, rst_n, branch, equal, predict, branchpred_his
 );
  input clk, rst_n, branch, equal;
  output predict, branchpred_his;

  assign predict = 1'b0;
  assign branchpred_his = 1'b0;

endmodule


module precontrolDec ( instruction_next, Jump_IF, Branch_IF );
  input [31:0] instruction_next;
  output Jump_IF, Branch_IF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  AND4X6 U1 ( .A(n8), .B(n7), .C(n6), .D(instruction_next[27]), .Y(Jump_IF) );
  INVX4 U2 ( .A(instruction_next[31]), .Y(n6) );
  NOR2X8 U3 ( .A(instruction_next[28]), .B(instruction_next[29]), .Y(n8) );
  INVX6 U4 ( .A(instruction_next[30]), .Y(n7) );
  INVXL U5 ( .A(instruction_next[28]), .Y(n1) );
  CLKINVX1 U6 ( .A(n1), .Y(n2) );
  NAND4XL U7 ( .A(n3), .B(n7), .C(n2), .D(n6), .Y(n4) );
  NOR3BXL U8 ( .AN(n5), .B(n4), .C(instruction_next[26]), .Y(Branch_IF) );
  INVXL U9 ( .A(instruction_next[29]), .Y(n3) );
  INVXL U10 ( .A(instruction_next[27]), .Y(n5) );
endmodule


module nextPCcalculator_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n8, n9, n11, n12, n14, n16, n17, n19, n21, n22, n23, n24,
         n26, n27, n28, n30, n33, n34, n36, n37, n38, n39, n40, n42, n43, n44,
         n46, n47, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n69, n70, n73, n74, n76, n77, n78, n79, n80,
         n81, n84, n86, n88, n89, n90, n91, n92, n93, n94, n95, n97, n99, n100,
         n101, n104, n105, n106, n107, n108, n109, n114, n115, n116, n117,
         n118, n120, n121, n122, n124, n125, n126, n130, n131, n132, n133,
         n134, n136, n138, n139, n140, n141, n142, n143, n144, n145, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n164, n166, n169, n171, n172, n174, n177, n178, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n191, n192, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n206, n207,
         n208, n209, n210, n211, n212, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n358, n359;
  assign n23 = A[30];
  assign n27 = A[29];
  assign n39 = A[27];
  assign n43 = A[26];
  assign n55 = A[24];
  assign n65 = A[22];
  assign n77 = A[20];

  AOI21X4 U86 ( .A0(n156), .A1(n88), .B0(n89), .Y(n1) );
  OAI21X4 U88 ( .A0(n125), .A1(n90), .B0(n91), .Y(n89) );
  AOI21X4 U90 ( .A0(n109), .A1(n92), .B0(n93), .Y(n91) );
  NOR2X8 U107 ( .A(B[16]), .B(A[16]), .Y(n101) );
  OAI21X4 U118 ( .A0(n114), .A1(n122), .B0(n115), .Y(n109) );
  AOI21X4 U140 ( .A0(n145), .A1(n130), .B0(n131), .Y(n125) );
  OAI21X4 U179 ( .A0(n185), .A1(n157), .B0(n158), .Y(n156) );
  NOR2X8 U182 ( .A(n166), .B(n161), .Y(n159) );
  NOR2X8 U186 ( .A(B[9]), .B(A[9]), .Y(n161) );
  OAI21X4 U205 ( .A0(n177), .A1(n183), .B0(n178), .Y(n172) );
  AOI21X4 U220 ( .A0(n186), .A1(n194), .B0(n187), .Y(n185) );
  OAI21X4 U222 ( .A0(n192), .A1(n188), .B0(n189), .Y(n187) );
  NOR2X8 U225 ( .A(B[5]), .B(A[5]), .Y(n188) );
  NOR2X8 U231 ( .A(B[4]), .B(A[4]), .Y(n191) );
  OAI21X4 U235 ( .A0(n195), .A1(n198), .B0(n196), .Y(n194) );
  OR2X6 U248 ( .A(n359), .B(n46), .Y(n333) );
  CLKBUFX2 U249 ( .A(n166), .Y(n315) );
  AOI21X2 U250 ( .A0(n329), .A1(n202), .B0(n120), .Y(n118) );
  AOI21X2 U251 ( .A0(n329), .A1(n108), .B0(n109), .Y(n107) );
  CLKBUFX8 U252 ( .A(n329), .Y(n316) );
  XOR2X2 U253 ( .A(n184), .B(n324), .Y(SUM[6]) );
  XOR2X1 U254 ( .A(n9), .B(n155), .Y(SUM[10]) );
  OR2X6 U255 ( .A(n359), .B(n42), .Y(n335) );
  OR2X6 U256 ( .A(n359), .B(n30), .Y(n334) );
  OR2X6 U257 ( .A(n359), .B(n36), .Y(n336) );
  OR2X6 U258 ( .A(n359), .B(n86), .Y(n354) );
  OR2X6 U259 ( .A(n359), .B(n54), .Y(n347) );
  OR2X6 U260 ( .A(n359), .B(n76), .Y(n348) );
  INVX3 U261 ( .A(n172), .Y(n174) );
  INVX2 U262 ( .A(n185), .Y(n184) );
  NAND2X1 U263 ( .A(n126), .B(n108), .Y(n106) );
  NOR2X4 U264 ( .A(n153), .B(n150), .Y(n144) );
  NOR2X6 U265 ( .A(B[10]), .B(A[10]), .Y(n153) );
  BUFX6 U266 ( .A(n198), .Y(n349) );
  XOR2X4 U267 ( .A(n331), .B(n317), .Y(SUM[4]) );
  NAND2X2 U268 ( .A(n212), .B(n192), .Y(n317) );
  NOR2X1 U269 ( .A(B[2]), .B(A[2]), .Y(n197) );
  XOR2X4 U270 ( .A(n319), .B(n318), .Y(SUM[7]) );
  CLKINVX20 U271 ( .A(n12), .Y(n318) );
  AO21X4 U272 ( .A0(n184), .A1(n210), .B0(n181), .Y(n319) );
  XNOR2X4 U273 ( .A(n320), .B(n11), .Y(SUM[8]) );
  AO21X4 U274 ( .A0(n184), .A1(n171), .B0(n343), .Y(n320) );
  OAI2BB1X4 U275 ( .A0N(n164), .A1N(n184), .B0(n321), .Y(n351) );
  OA21X4 U276 ( .A0(n174), .A1(n315), .B0(n169), .Y(n321) );
  XNOR2X4 U277 ( .A(n57), .B(n322), .Y(SUM[24]) );
  CLKINVX20 U278 ( .A(n340), .Y(n322) );
  XOR2X4 U279 ( .A(n323), .B(n14), .Y(SUM[5]) );
  OA21X4 U280 ( .A0(n331), .A1(n191), .B0(n192), .Y(n323) );
  CLKAND2X8 U281 ( .A(n210), .B(n183), .Y(n324) );
  OR2X4 U282 ( .A(B[11]), .B(A[11]), .Y(n325) );
  AOI2BB1X4 U283 ( .A0N(n155), .A1N(n97), .B0(n326), .Y(n339) );
  AO21X4 U284 ( .A0(n329), .A1(n99), .B0(n100), .Y(n326) );
  INVXL U285 ( .A(n166), .Y(n208) );
  NOR2X8 U286 ( .A(B[17]), .B(A[17]), .Y(n94) );
  NAND2X6 U287 ( .A(B[14]), .B(A[14]), .Y(n122) );
  NOR2X4 U288 ( .A(B[14]), .B(A[14]), .Y(n121) );
  NOR2X6 U289 ( .A(n101), .B(n94), .Y(n92) );
  OR2X6 U290 ( .A(n359), .B(n26), .Y(n338) );
  NAND2X8 U291 ( .A(B[10]), .B(A[10]), .Y(n154) );
  NOR2X6 U292 ( .A(B[12]), .B(A[12]), .Y(n139) );
  NOR2X6 U293 ( .A(B[6]), .B(A[6]), .Y(n182) );
  NOR2X4 U294 ( .A(n191), .B(n188), .Y(n186) );
  CLKAND2X3 U295 ( .A(n144), .B(n204), .Y(n353) );
  CLKAND2X3 U296 ( .A(n203), .B(n133), .Y(n332) );
  CLKAND2X3 U297 ( .A(n200), .B(n104), .Y(n350) );
  INVX1 U298 ( .A(n56), .Y(n340) );
  CLKINVX1 U299 ( .A(n24), .Y(n337) );
  AND2X2 U300 ( .A(n207), .B(n162), .Y(n352) );
  BUFX4 U301 ( .A(A[1]), .Y(SUM[1]) );
  BUFX4 U302 ( .A(A[0]), .Y(SUM[0]) );
  NOR2BX4 U303 ( .AN(n21), .B(n359), .Y(n19) );
  NOR2X2 U304 ( .A(n22), .B(n30), .Y(n21) );
  OA21X1 U305 ( .A0(n198), .A1(n195), .B0(n196), .Y(n331) );
  NOR2X6 U306 ( .A(n139), .B(n132), .Y(n130) );
  NAND2X6 U307 ( .A(n159), .B(n171), .Y(n157) );
  OA21X4 U308 ( .A0(n114), .A1(n122), .B0(n115), .Y(n327) );
  NOR2X8 U309 ( .A(B[15]), .B(A[15]), .Y(n114) );
  NOR2X8 U310 ( .A(B[17]), .B(A[17]), .Y(n328) );
  NAND2X6 U311 ( .A(A[6]), .B(B[6]), .Y(n183) );
  NOR2X8 U312 ( .A(B[7]), .B(A[7]), .Y(n177) );
  AOI21X1 U313 ( .A0(n204), .A1(n145), .B0(n138), .Y(n136) );
  AO21X4 U314 ( .A0(n145), .A1(n130), .B0(n131), .Y(n329) );
  NAND2X6 U315 ( .A(n344), .B(n133), .Y(n131) );
  OR2XL U316 ( .A(B[3]), .B(A[3]), .Y(n330) );
  XOR2X4 U317 ( .A(n134), .B(n332), .Y(SUM[13]) );
  INVX3 U318 ( .A(n17), .Y(SUM[2]) );
  NAND2BX2 U319 ( .AN(n197), .B(n349), .Y(n17) );
  XOR2X4 U320 ( .A(n333), .B(n44), .Y(SUM[26]) );
  NOR2X4 U321 ( .A(n359), .B(n64), .Y(n63) );
  XOR2X4 U322 ( .A(n334), .B(n28), .Y(SUM[29]) );
  XOR2X4 U323 ( .A(n335), .B(n40), .Y(SUM[27]) );
  XOR2X4 U324 ( .A(n336), .B(n34), .Y(SUM[28]) );
  XOR2X1 U325 ( .A(n16), .B(n349), .Y(SUM[3]) );
  XNOR2X4 U326 ( .A(n338), .B(n337), .Y(SUM[30]) );
  XOR2X2 U327 ( .A(n86), .B(n359), .Y(SUM[18]) );
  XOR2X4 U328 ( .A(n339), .B(n2), .Y(SUM[17]) );
  AOI2BB1X4 U329 ( .A0N(n155), .A1N(n124), .B0(n316), .Y(n346) );
  OAI21X4 U330 ( .A0(n117), .A1(n155), .B0(n118), .Y(n116) );
  XOR2X4 U331 ( .A(n19), .B(A[31]), .Y(SUM[31]) );
  INVXL U332 ( .A(n191), .Y(n212) );
  NAND2X1 U333 ( .A(n330), .B(n196), .Y(n16) );
  XOR2X4 U334 ( .A(n346), .B(n341), .Y(SUM[14]) );
  NAND2X2 U335 ( .A(n202), .B(n122), .Y(n341) );
  INVX4 U336 ( .A(n200), .Y(n342) );
  INVX2 U337 ( .A(n101), .Y(n200) );
  NOR2X8 U338 ( .A(n86), .B(n84), .Y(n81) );
  INVX4 U339 ( .A(A[18]), .Y(n86) );
  NAND2X8 U340 ( .A(n81), .B(n73), .Y(n70) );
  INVX3 U341 ( .A(n174), .Y(n343) );
  NAND2X4 U342 ( .A(B[9]), .B(A[9]), .Y(n162) );
  OR2X6 U343 ( .A(n132), .B(n140), .Y(n344) );
  NAND2X2 U344 ( .A(B[13]), .B(A[13]), .Y(n133) );
  CLKBUFX2 U345 ( .A(n154), .Y(n345) );
  NOR2X4 U346 ( .A(n70), .B(n359), .Y(n67) );
  NOR2X4 U347 ( .A(n80), .B(n359), .Y(n79) );
  XOR2X4 U348 ( .A(n347), .B(n52), .Y(SUM[25]) );
  XOR2X4 U349 ( .A(n348), .B(n74), .Y(SUM[21]) );
  NOR2X4 U350 ( .A(n58), .B(n359), .Y(n57) );
  INVX6 U351 ( .A(A[25]), .Y(n52) );
  XOR2X4 U352 ( .A(n63), .B(A[23]), .Y(SUM[23]) );
  INVX6 U353 ( .A(A[23]), .Y(n62) );
  INVX6 U354 ( .A(A[21]), .Y(n74) );
  OAI21X4 U355 ( .A0(n106), .A1(n155), .B0(n107), .Y(n105) );
  NAND2X1 U356 ( .A(n208), .B(n169), .Y(n11) );
  INVX8 U357 ( .A(n156), .Y(n155) );
  OAI21X4 U358 ( .A0(n327), .A1(n342), .B0(n104), .Y(n100) );
  NOR2X6 U359 ( .A(n182), .B(n177), .Y(n171) );
  NAND2X6 U360 ( .A(B[2]), .B(A[2]), .Y(n198) );
  INVX2 U361 ( .A(n132), .Y(n203) );
  XOR2X4 U362 ( .A(n105), .B(n350), .Y(SUM[16]) );
  OR2X8 U363 ( .A(n150), .B(n154), .Y(n355) );
  XOR2X4 U364 ( .A(n351), .B(n352), .Y(SUM[9]) );
  NOR2X6 U365 ( .A(n34), .B(n38), .Y(n33) );
  NAND2X4 U366 ( .A(n39), .B(n43), .Y(n38) );
  INVX6 U367 ( .A(n121), .Y(n202) );
  NAND2X6 U368 ( .A(n61), .B(n51), .Y(n50) );
  NOR2X8 U369 ( .A(n66), .B(n62), .Y(n61) );
  NOR2X4 U370 ( .A(n56), .B(n52), .Y(n51) );
  NOR2X8 U371 ( .A(B[13]), .B(A[13]), .Y(n132) );
  OAI2BB1X1 U372 ( .A0N(n353), .A1N(n156), .B0(n136), .Y(n134) );
  NOR2BX1 U373 ( .AN(n171), .B(n166), .Y(n164) );
  NAND2X1 U374 ( .A(n47), .B(n37), .Y(n36) );
  XNOR2X4 U375 ( .A(n67), .B(n66), .Y(SUM[22]) );
  OAI21X4 U376 ( .A0(n142), .A1(n155), .B0(n143), .Y(n141) );
  XNOR2X4 U377 ( .A(n152), .B(n8), .Y(SUM[11]) );
  OAI21X4 U378 ( .A0(n153), .A1(n155), .B0(n345), .Y(n152) );
  NAND2X2 U379 ( .A(n126), .B(n202), .Y(n117) );
  NAND2X4 U380 ( .A(n99), .B(n126), .Y(n97) );
  CLKINVX8 U381 ( .A(n124), .Y(n126) );
  INVX3 U382 ( .A(n153), .Y(n206) );
  INVX8 U383 ( .A(n77), .Y(n78) );
  NOR2X6 U384 ( .A(n78), .B(n74), .Y(n73) );
  XOR2X4 U385 ( .A(n354), .B(n84), .Y(SUM[19]) );
  INVX4 U386 ( .A(A[19]), .Y(n84) );
  NOR2X8 U387 ( .A(B[8]), .B(A[8]), .Y(n166) );
  NAND2X2 U388 ( .A(n209), .B(n178), .Y(n12) );
  NAND2X4 U389 ( .A(B[8]), .B(A[8]), .Y(n169) );
  NOR2X8 U390 ( .A(n70), .B(n50), .Y(n47) );
  NOR2X4 U391 ( .A(n70), .B(n60), .Y(n59) );
  CLKINVX2 U392 ( .A(n70), .Y(n69) );
  NAND2X8 U393 ( .A(B[12]), .B(A[12]), .Y(n140) );
  INVX1 U394 ( .A(n47), .Y(n46) );
  AOI21X4 U395 ( .A0(n172), .A1(n159), .B0(n160), .Y(n158) );
  NAND2X8 U396 ( .A(n355), .B(n151), .Y(n145) );
  NAND2X4 U397 ( .A(A[11]), .B(B[11]), .Y(n151) );
  OAI21X4 U398 ( .A0(n328), .A1(n104), .B0(n95), .Y(n93) );
  NAND2X4 U399 ( .A(B[17]), .B(A[17]), .Y(n95) );
  NAND2X1 U400 ( .A(n47), .B(n43), .Y(n42) );
  XNOR2X4 U401 ( .A(n79), .B(n78), .Y(SUM[20]) );
  NAND2X4 U402 ( .A(B[15]), .B(A[15]), .Y(n115) );
  XOR2X4 U403 ( .A(n141), .B(n358), .Y(SUM[12]) );
  INVX2 U404 ( .A(n59), .Y(n58) );
  NAND2X1 U405 ( .A(n59), .B(n55), .Y(n54) );
  XNOR2X4 U406 ( .A(n116), .B(n4), .Y(SUM[15]) );
  INVX6 U407 ( .A(n182), .Y(n210) );
  INVX4 U408 ( .A(n65), .Y(n66) );
  NAND2BX4 U409 ( .AN(n30), .B(n27), .Y(n26) );
  NOR2X8 U410 ( .A(B[11]), .B(A[11]), .Y(n150) );
  CLKINVX6 U411 ( .A(n139), .Y(n204) );
  NAND2X4 U412 ( .A(n47), .B(n33), .Y(n30) );
  INVXL U413 ( .A(n145), .Y(n143) );
  NAND2X4 U414 ( .A(B[3]), .B(A[3]), .Y(n196) );
  NAND2X8 U415 ( .A(n144), .B(n130), .Y(n124) );
  NAND2XL U416 ( .A(n206), .B(n154), .Y(n9) );
  NOR2BX4 U417 ( .AN(n108), .B(n342), .Y(n99) );
  NAND2X6 U418 ( .A(B[16]), .B(A[16]), .Y(n104) );
  NAND2X4 U419 ( .A(A[5]), .B(B[5]), .Y(n189) );
  INVX3 U420 ( .A(A[28]), .Y(n34) );
  NOR2X4 U421 ( .A(n124), .B(n90), .Y(n88) );
  NAND2X8 U422 ( .A(n108), .B(n92), .Y(n90) );
  NAND2XL U423 ( .A(n325), .B(n151), .Y(n8) );
  INVXL U424 ( .A(n38), .Y(n37) );
  OAI21X4 U425 ( .A0(n169), .A1(n161), .B0(n162), .Y(n160) );
  INVXL U426 ( .A(n81), .Y(n80) );
  NOR2X8 U427 ( .A(n121), .B(n114), .Y(n108) );
  INVX6 U428 ( .A(n55), .Y(n56) );
  NAND2X2 U429 ( .A(n69), .B(n65), .Y(n64) );
  BUFX20 U430 ( .A(n1), .Y(n359) );
  INVXL U431 ( .A(n144), .Y(n142) );
  NAND2X1 U432 ( .A(n201), .B(n115), .Y(n4) );
  INVXL U433 ( .A(n114), .Y(n201) );
  NAND2X1 U434 ( .A(n199), .B(n95), .Y(n2) );
  INVXL U435 ( .A(n328), .Y(n199) );
  NAND2X1 U436 ( .A(n211), .B(n189), .Y(n14) );
  INVXL U437 ( .A(n188), .Y(n211) );
  INVXL U438 ( .A(n122), .Y(n120) );
  CLKINVX1 U439 ( .A(n140), .Y(n138) );
  AND2XL U440 ( .A(n204), .B(n140), .Y(n358) );
  CLKINVX1 U441 ( .A(n61), .Y(n60) );
  INVXL U442 ( .A(n183), .Y(n181) );
  INVXL U443 ( .A(n177), .Y(n209) );
  INVXL U444 ( .A(n161), .Y(n207) );
  NAND2X6 U445 ( .A(A[4]), .B(B[4]), .Y(n192) );
  NAND2X4 U446 ( .A(B[7]), .B(A[7]), .Y(n178) );
  CLKINVX1 U447 ( .A(n43), .Y(n44) );
  NAND2XL U448 ( .A(n81), .B(n77), .Y(n76) );
  NAND2X1 U449 ( .A(n23), .B(n27), .Y(n22) );
  CLKINVX1 U450 ( .A(n39), .Y(n40) );
  CLKINVX1 U451 ( .A(n23), .Y(n24) );
  CLKINVX1 U452 ( .A(n27), .Y(n28) );
  NOR2X6 U453 ( .A(A[3]), .B(B[3]), .Y(n195) );
endmodule


module nextPCcalculator ( PCcur, PCplus4, PCplus4_regD, targetAddr, 
        branchOffset_I, branchOffset_regD, JumpRegAddr, PCsrc, PCnext );
  input [31:0] PCcur;
  input [31:0] PCplus4;
  input [31:0] PCplus4_regD;
  input [25:0] targetAddr;
  input [15:0] branchOffset_I;
  input [15:0] branchOffset_regD;
  input [31:0] JumpRegAddr;
  input [2:0] PCsrc;
  output [31:0] PCnext;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170;
  wire   [31:0] PCplus4_actual;
  wire   [17:2] branchOffset_actual;
  wire   [31:0] ADDresult;

  nextPCcalculator_DW01_add_1 add_1346 ( .A(PCplus4_actual), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        branchOffset_actual, 1'b0, 1'b0}), .CI(1'b0), .SUM(ADDresult) );
  MX2X8 U4 ( .A(PCplus4_regD[8]), .B(PCplus4[8]), .S0(n15), .Y(
        PCplus4_actual[8]) );
  MX2X8 U5 ( .A(branchOffset_regD[7]), .B(branchOffset_I[7]), .S0(n15), .Y(
        branchOffset_actual[9]) );
  CLKMX2X6 U6 ( .A(PCplus4_regD[9]), .B(PCplus4[9]), .S0(n15), .Y(
        PCplus4_actual[9]) );
  NAND2X2 U7 ( .A(n35), .B(n36), .Y(PCnext[0]) );
  AOI222X2 U8 ( .A0(JumpRegAddr[2]), .A1(n23), .B0(targetAddr[0]), .B1(n16), 
        .C0(ADDresult[2]), .C1(n25), .Y(n43) );
  AOI222X2 U9 ( .A0(JumpRegAddr[6]), .A1(n23), .B0(targetAddr[4]), .B1(n17), 
        .C0(ADDresult[6]), .C1(n25), .Y(n59) );
  AOI222X2 U10 ( .A0(JumpRegAddr[4]), .A1(n23), .B0(targetAddr[2]), .B1(n17), 
        .C0(ADDresult[4]), .C1(n25), .Y(n51) );
  OAI211X2 U11 ( .A0(n18), .A1(n65), .B0(n64), .C0(n63), .Y(PCnext[7]) );
  INVX1 U12 ( .A(n125), .Y(n12) );
  NOR2X6 U13 ( .A(n8), .B(n9), .Y(PCnext[26]) );
  INVX8 U14 ( .A(ADDresult[12]), .Y(n84) );
  MX2X8 U15 ( .A(PCplus4_regD[12]), .B(PCplus4[12]), .S0(n15), .Y(
        PCplus4_actual[12]) );
  CLKINVX20 U16 ( .A(n19), .Y(n18) );
  NAND3X4 U17 ( .A(n152), .B(n151), .C(n150), .Y(n153) );
  INVX8 U18 ( .A(n5), .Y(n1) );
  INVX2 U19 ( .A(n42), .Y(n5) );
  AOI222X2 U20 ( .A0(PCplus4_regD[22]), .A1(n143), .B0(targetAddr[20]), .B1(
        n16), .C0(JumpRegAddr[22]), .C1(n24), .Y(n124) );
  INVX20 U21 ( .A(n14), .Y(n143) );
  NAND2X4 U22 ( .A(n116), .B(n115), .Y(n117) );
  AOI222X4 U23 ( .A0(PCplus4_regD[20]), .A1(n143), .B0(targetAddr[18]), .B1(
        n16), .C0(JumpRegAddr[20]), .C1(n24), .Y(n116) );
  INVX8 U24 ( .A(PCsrc[1]), .Y(n42) );
  CLKINVX3 U25 ( .A(PCsrc[2]), .Y(n41) );
  MX2X4 U26 ( .A(PCplus4_regD[14]), .B(PCplus4[14]), .S0(n7), .Y(
        PCplus4_actual[14]) );
  CLKMX2X12 U27 ( .A(PCplus4_regD[10]), .B(PCplus4[10]), .S0(n30), .Y(
        PCplus4_actual[10]) );
  MX2X6 U28 ( .A(branchOffset_regD[6]), .B(branchOffset_I[6]), .S0(n15), .Y(
        branchOffset_actual[8]) );
  INVX6 U29 ( .A(n31), .Y(n6) );
  BUFX12 U30 ( .A(n20), .Y(n19) );
  INVX4 U31 ( .A(n26), .Y(n11) );
  INVXL U32 ( .A(PCcur[26]), .Y(n2) );
  NAND3BX1 U33 ( .AN(n6), .B(n41), .C(n5), .Y(n163) );
  NAND3BX1 U34 ( .AN(n1), .B(n13), .C(n31), .Y(n32) );
  NAND2X8 U35 ( .A(n1), .B(n13), .Y(n105) );
  INVX4 U36 ( .A(n32), .Y(n164) );
  INVX8 U37 ( .A(n105), .Y(n169) );
  NAND3BX1 U38 ( .AN(n6), .B(n1), .C(n41), .Y(n148) );
  NAND3BX2 U39 ( .AN(n1), .B(n6), .C(n41), .Y(n149) );
  CLKMX2X12 U40 ( .A(PCplus4_regD[17]), .B(PCplus4[17]), .S0(n7), .Y(
        PCplus4_actual[17]) );
  CLKMX2X12 U41 ( .A(branchOffset_regD[15]), .B(branchOffset_I[15]), .S0(n7), 
        .Y(branchOffset_actual[17]) );
  OAI211X2 U42 ( .A0(n18), .A1(n57), .B0(n56), .C0(n55), .Y(PCnext[5]) );
  MX2X8 U43 ( .A(PCplus4_regD[4]), .B(PCplus4[4]), .S0(n30), .Y(
        PCplus4_actual[4]) );
  OA22XL U44 ( .A0(n2), .A1(n33), .B0(n18), .B1(n138), .Y(n139) );
  NAND3BX2 U45 ( .AN(n5), .B(n6), .C(n41), .Y(n33) );
  MX2X8 U46 ( .A(branchOffset_regD[1]), .B(branchOffset_I[1]), .S0(n30), .Y(
        branchOffset_actual[3]) );
  MX2X6 U47 ( .A(PCplus4_regD[3]), .B(PCplus4[3]), .S0(n30), .Y(
        PCplus4_actual[3]) );
  CLKINVX3 U48 ( .A(n148), .Y(n20) );
  NAND3X2 U49 ( .A(n156), .B(n155), .C(n154), .Y(n157) );
  AOI22X1 U50 ( .A0(n165), .A1(PCplus4[29]), .B0(JumpRegAddr[29]), .B1(n23), 
        .Y(n154) );
  INVX8 U51 ( .A(ADDresult[17]), .Y(n104) );
  INVX6 U52 ( .A(ADDresult[11]), .Y(n80) );
  AOI222X4 U53 ( .A0(PCplus4_regD[23]), .A1(n143), .B0(targetAddr[21]), .B1(
        n16), .C0(JumpRegAddr[23]), .C1(n24), .Y(n128) );
  BUFX12 U54 ( .A(n142), .Y(n16) );
  AOI222X4 U55 ( .A0(PCplus4_regD[0]), .A1(n143), .B0(ADDresult[0]), .B1(n25), 
        .C0(JumpRegAddr[0]), .C1(n23), .Y(n36) );
  NOR2X6 U56 ( .A(ADDresult[26]), .B(n141), .Y(n8) );
  CLKINVX3 U57 ( .A(PCsrc[0]), .Y(n31) );
  MX2X8 U58 ( .A(branchOffset_regD[2]), .B(branchOffset_I[2]), .S0(n30), .Y(
        branchOffset_actual[4]) );
  NAND2X2 U59 ( .A(n39), .B(n38), .Y(PCnext[1]) );
  AOI222X4 U60 ( .A0(PCplus4_regD[1]), .A1(n143), .B0(ADDresult[1]), .B1(n25), 
        .C0(JumpRegAddr[1]), .C1(n23), .Y(n39) );
  AOI222X4 U61 ( .A0(PCplus4_regD[18]), .A1(n143), .B0(targetAddr[16]), .B1(
        n16), .C0(JumpRegAddr[18]), .C1(n24), .Y(n108) );
  MX2X6 U62 ( .A(branchOffset_regD[13]), .B(branchOffset_I[13]), .S0(n7), .Y(
        branchOffset_actual[15]) );
  AOI22X1 U63 ( .A0(n165), .A1(PCplus4[31]), .B0(JumpRegAddr[31]), .B1(n23), 
        .Y(n166) );
  AOI22X1 U64 ( .A0(n165), .A1(PCplus4[30]), .B0(JumpRegAddr[30]), .B1(n23), 
        .Y(n158) );
  CLKMX2X4 U65 ( .A(branchOffset_regD[8]), .B(branchOffset_I[8]), .S0(n30), 
        .Y(branchOffset_actual[10]) );
  MX2X6 U66 ( .A(PCplus4_regD[15]), .B(PCplus4[15]), .S0(n7), .Y(
        PCplus4_actual[15]) );
  MX2X8 U67 ( .A(branchOffset_regD[3]), .B(branchOffset_I[3]), .S0(n30), .Y(
        branchOffset_actual[5]) );
  MX2X8 U68 ( .A(PCplus4_regD[5]), .B(PCplus4[5]), .S0(n30), .Y(
        PCplus4_actual[5]) );
  AOI222X4 U69 ( .A0(JumpRegAddr[3]), .A1(n23), .B0(targetAddr[1]), .B1(n16), 
        .C0(ADDresult[3]), .C1(n25), .Y(n47) );
  NAND2X1 U70 ( .A(n124), .B(n123), .Y(n125) );
  CLKMX2X12 U71 ( .A(branchOffset_regD[14]), .B(branchOffset_I[14]), .S0(n7), 
        .Y(branchOffset_actual[16]) );
  CLKMX2X12 U72 ( .A(PCplus4_regD[16]), .B(PCplus4[16]), .S0(n7), .Y(
        PCplus4_actual[16]) );
  AOI222X2 U73 ( .A0(JumpRegAddr[5]), .A1(n23), .B0(targetAddr[3]), .B1(n17), 
        .C0(ADDresult[5]), .C1(n25), .Y(n55) );
  AOI222X4 U74 ( .A0(PCplus4_regD[19]), .A1(n143), .B0(targetAddr[17]), .B1(
        n16), .C0(JumpRegAddr[19]), .C1(n24), .Y(n112) );
  AOI222X4 U75 ( .A0(PCplus4_regD[25]), .A1(n143), .B0(targetAddr[23]), .B1(
        n16), .C0(JumpRegAddr[25]), .C1(n24), .Y(n136) );
  AOI2BB2X1 U76 ( .B0(PCcur[21]), .B1(n21), .A0N(n18), .A1N(n118), .Y(n119) );
  AOI222X4 U77 ( .A0(PCplus4_regD[21]), .A1(n143), .B0(targetAddr[19]), .B1(
        n16), .C0(JumpRegAddr[21]), .C1(n24), .Y(n120) );
  CLKMX2X3 U78 ( .A(PCplus4_regD[25]), .B(PCplus4[25]), .S0(n7), .Y(
        PCplus4_actual[25]) );
  OAI211X2 U79 ( .A0(n105), .A1(n88), .B0(n87), .C0(n86), .Y(PCnext[13]) );
  CLKMX2X3 U80 ( .A(PCplus4_regD[21]), .B(PCplus4[21]), .S0(n7), .Y(
        PCplus4_actual[21]) );
  AOI2BB2XL U81 ( .B0(PCcur[25]), .B1(n21), .A0N(n18), .A1N(n134), .Y(n135) );
  INVX4 U82 ( .A(n41), .Y(n13) );
  AOI222X1 U83 ( .A0(PCplus4_regD[24]), .A1(n143), .B0(targetAddr[22]), .B1(
        n16), .C0(JumpRegAddr[24]), .C1(n24), .Y(n132) );
  OA22X4 U84 ( .A0(ADDresult[30]), .A1(n161), .B0(n26), .B1(n161), .Y(
        PCnext[30]) );
  OA22X4 U85 ( .A0(ADDresult[31]), .A1(n170), .B0(n26), .B1(n170), .Y(
        PCnext[31]) );
  OA22X4 U86 ( .A0(ADDresult[28]), .A1(n153), .B0(n26), .B1(n153), .Y(
        PCnext[28]) );
  AOI2BB2X4 U87 ( .B0(n11), .B1(n12), .A0N(ADDresult[22]), .A1N(n125), .Y(
        PCnext[22]) );
  OAI211X2 U88 ( .A0(n105), .A1(n84), .B0(n83), .C0(n82), .Y(PCnext[12]) );
  INVX6 U89 ( .A(ADDresult[16]), .Y(n100) );
  OAI211X2 U90 ( .A0(n18), .A1(n73), .B0(n72), .C0(n71), .Y(PCnext[9]) );
  OA22X4 U91 ( .A0(ADDresult[29]), .A1(n157), .B0(n26), .B1(n157), .Y(
        PCnext[29]) );
  OAI211X2 U92 ( .A0(n105), .A1(n96), .B0(n95), .C0(n94), .Y(PCnext[15]) );
  INVX6 U93 ( .A(ADDresult[15]), .Y(n96) );
  CLKMX2X4 U94 ( .A(branchOffset_regD[5]), .B(branchOffset_I[5]), .S0(n30), 
        .Y(branchOffset_actual[7]) );
  OAI211X2 U95 ( .A0(n18), .A1(n53), .B0(n52), .C0(n51), .Y(PCnext[4]) );
  OA22X4 U96 ( .A0(ADDresult[25]), .A1(n137), .B0(n26), .B1(n137), .Y(
        PCnext[25]) );
  OAI211X2 U97 ( .A0(n92), .A1(n105), .B0(n91), .C0(n90), .Y(PCnext[14]) );
  INVX6 U98 ( .A(ADDresult[14]), .Y(n92) );
  CLKBUFX20 U99 ( .A(n29), .Y(n7) );
  BUFX20 U100 ( .A(n29), .Y(n15) );
  AOI2BB2X4 U101 ( .B0(n11), .B1(n10), .A0N(ADDresult[20]), .A1N(n117), .Y(
        PCnext[20]) );
  BUFX20 U102 ( .A(n164), .Y(n24) );
  MX2X8 U103 ( .A(branchOffset_regD[10]), .B(branchOffset_I[10]), .S0(n15), 
        .Y(branchOffset_actual[12]) );
  INVX4 U104 ( .A(ADDresult[13]), .Y(n88) );
  CLKMX2X4 U105 ( .A(PCplus4_regD[7]), .B(PCplus4[7]), .S0(n30), .Y(
        PCplus4_actual[7]) );
  CLKINVX8 U106 ( .A(n27), .Y(n29) );
  CLKINVX12 U107 ( .A(n28), .Y(n30) );
  AOI222X4 U108 ( .A0(PCplus4_regD[26]), .A1(n143), .B0(targetAddr[24]), .B1(
        n16), .C0(JumpRegAddr[26]), .C1(n24), .Y(n140) );
  INVX4 U109 ( .A(n149), .Y(n142) );
  BUFX20 U110 ( .A(n162), .Y(n21) );
  INVX4 U111 ( .A(n33), .Y(n162) );
  AOI22X1 U112 ( .A0(n165), .A1(PCplus4[28]), .B0(JumpRegAddr[28]), .B1(n23), 
        .Y(n150) );
  CLKMX2X8 U113 ( .A(PCplus4_regD[20]), .B(PCplus4[20]), .S0(n7), .Y(
        PCplus4_actual[20]) );
  AOI222X2 U114 ( .A0(JumpRegAddr[7]), .A1(n23), .B0(targetAddr[5]), .B1(n17), 
        .C0(ADDresult[7]), .C1(n25), .Y(n63) );
  CLKMX2X3 U115 ( .A(PCplus4_regD[19]), .B(PCplus4[19]), .S0(n7), .Y(
        PCplus4_actual[19]) );
  OAI211X2 U116 ( .A0(n100), .A1(n105), .B0(n99), .C0(n98), .Y(PCnext[16]) );
  NOR2X2 U117 ( .A(n26), .B(n141), .Y(n9) );
  NAND2X4 U118 ( .A(n140), .B(n139), .Y(n141) );
  OA22X4 U119 ( .A0(ADDresult[19]), .A1(n113), .B0(n25), .B1(n113), .Y(
        PCnext[19]) );
  OA22X4 U120 ( .A0(ADDresult[27]), .A1(n147), .B0(n26), .B1(n147), .Y(
        PCnext[27]) );
  OAI211X2 U121 ( .A0(n104), .A1(n105), .B0(n103), .C0(n102), .Y(PCnext[17])
         );
  CLKMX2X4 U122 ( .A(PCplus4_regD[6]), .B(PCplus4[6]), .S0(n30), .Y(
        PCplus4_actual[6]) );
  NAND3BX4 U123 ( .AN(PCsrc[0]), .B(n42), .C(PCsrc[2]), .Y(n28) );
  CLKMX2X6 U124 ( .A(branchOffset_regD[4]), .B(branchOffset_I[4]), .S0(n15), 
        .Y(branchOffset_actual[6]) );
  OAI211X2 U125 ( .A0(n18), .A1(n69), .B0(n67), .C0(n68), .Y(PCnext[8]) );
  CLKMX2X4 U126 ( .A(PCplus4_regD[2]), .B(PCplus4[2]), .S0(n30), .Y(
        PCplus4_actual[2]) );
  AOI222X2 U127 ( .A0(JumpRegAddr[8]), .A1(n23), .B0(targetAddr[6]), .B1(n17), 
        .C0(ADDresult[8]), .C1(n25), .Y(n67) );
  CLKMX2X4 U128 ( .A(branchOffset_regD[0]), .B(branchOffset_I[0]), .S0(n30), 
        .Y(branchOffset_actual[2]) );
  OAI211X2 U129 ( .A0(n105), .A1(n80), .B0(n79), .C0(n78), .Y(PCnext[11]) );
  BUFX20 U130 ( .A(n169), .Y(n26) );
  MX2X6 U131 ( .A(branchOffset_regD[11]), .B(branchOffset_I[11]), .S0(n15), 
        .Y(branchOffset_actual[13]) );
  MX2X6 U132 ( .A(PCplus4_regD[13]), .B(PCplus4[13]), .S0(n15), .Y(
        PCplus4_actual[13]) );
  AOI222X2 U133 ( .A0(JumpRegAddr[9]), .A1(n23), .B0(targetAddr[7]), .B1(n17), 
        .C0(ADDresult[9]), .C1(n25), .Y(n71) );
  BUFX20 U134 ( .A(n164), .Y(n23) );
  NAND3BX4 U135 ( .AN(PCsrc[0]), .B(n42), .C(PCsrc[2]), .Y(n27) );
  AOI222X1 U136 ( .A0(PCplus4_regD[27]), .A1(n143), .B0(targetAddr[25]), .B1(
        n17), .C0(JumpRegAddr[27]), .C1(n23), .Y(n146) );
  MX2X6 U137 ( .A(branchOffset_regD[9]), .B(branchOffset_I[9]), .S0(n15), .Y(
        branchOffset_actual[11]) );
  MX2X6 U138 ( .A(PCplus4_regD[11]), .B(PCplus4[11]), .S0(n30), .Y(
        PCplus4_actual[11]) );
  BUFX20 U139 ( .A(n169), .Y(n25) );
  BUFX16 U140 ( .A(n162), .Y(n22) );
  NAND2X2 U141 ( .A(n149), .B(n18), .Y(n165) );
  MX2XL U142 ( .A(PCplus4_regD[28]), .B(PCplus4[28]), .S0(n7), .Y(
        PCplus4_actual[28]) );
  MX2XL U143 ( .A(PCplus4_regD[30]), .B(PCplus4[30]), .S0(n7), .Y(
        PCplus4_actual[30]) );
  MX2XL U144 ( .A(PCplus4_regD[31]), .B(PCplus4[31]), .S0(n7), .Y(
        PCplus4_actual[31]) );
  BUFX12 U145 ( .A(n142), .Y(n17) );
  INVXL U146 ( .A(PCplus4[26]), .Y(n138) );
  INVXL U147 ( .A(PCplus4[19]), .Y(n110) );
  INVXL U148 ( .A(PCplus4[18]), .Y(n106) );
  NAND2X2 U149 ( .A(n25), .B(ADDresult[10]), .Y(n74) );
  INVXL U150 ( .A(PCplus4[14]), .Y(n89) );
  INVXL U151 ( .A(PCplus4[27]), .Y(n144) );
  INVX1 U152 ( .A(PCplus4[25]), .Y(n134) );
  INVXL U153 ( .A(PCplus4[24]), .Y(n130) );
  INVXL U154 ( .A(PCplus4[23]), .Y(n126) );
  INVXL U155 ( .A(PCplus4[21]), .Y(n118) );
  INVXL U156 ( .A(PCplus4[13]), .Y(n85) );
  INVXL U157 ( .A(PCplus4[16]), .Y(n97) );
  INVXL U158 ( .A(PCplus4[17]), .Y(n101) );
  INVXL U159 ( .A(PCplus4[15]), .Y(n93) );
  INVX1 U160 ( .A(PCplus4[11]), .Y(n77) );
  CLKMX2X4 U161 ( .A(PCplus4_regD[27]), .B(PCplus4[27]), .S0(n7), .Y(
        PCplus4_actual[27]) );
  CLKMX2X4 U162 ( .A(PCplus4_regD[22]), .B(PCplus4[22]), .S0(n7), .Y(
        PCplus4_actual[22]) );
  MX2X2 U163 ( .A(PCplus4_regD[18]), .B(PCplus4[18]), .S0(n7), .Y(
        PCplus4_actual[18]) );
  AOI2BB2XL U164 ( .B0(PCcur[27]), .B1(n21), .A0N(n18), .A1N(n144), .Y(n145)
         );
  NAND2XL U165 ( .A(PCcur[29]), .B(n21), .Y(n156) );
  AOI2BB2XL U166 ( .B0(PCcur[0]), .B1(n21), .A0N(n18), .A1N(n34), .Y(n35) );
  CLKMX2X4 U167 ( .A(PCplus4_regD[29]), .B(PCplus4[29]), .S0(n7), .Y(
        PCplus4_actual[29]) );
  AOI2BB2XL U168 ( .B0(PCcur[20]), .B1(n21), .A0N(n18), .A1N(n114), .Y(n115)
         );
  AOI2BB2XL U169 ( .B0(PCcur[22]), .B1(n21), .A0N(n18), .A1N(n122), .Y(n123)
         );
  INVXL U170 ( .A(PCplus4[22]), .Y(n122) );
  INVXL U171 ( .A(PCplus4[3]), .Y(n49) );
  AOI2BB2XL U172 ( .B0(PCcur[6]), .B1(n22), .A0N(n14), .A1N(n58), .Y(n60) );
  MX2X6 U173 ( .A(branchOffset_regD[12]), .B(branchOffset_I[12]), .S0(n15), 
        .Y(branchOffset_actual[14]) );
  NAND3BX2 U174 ( .AN(n76), .B(n74), .C(n75), .Y(PCnext[10]) );
  CLKMX2X4 U175 ( .A(PCplus4_regD[26]), .B(PCplus4[26]), .S0(n7), .Y(
        PCplus4_actual[26]) );
  NAND2X2 U176 ( .A(n120), .B(n119), .Y(n121) );
  NAND2X2 U177 ( .A(n107), .B(n108), .Y(n109) );
  AOI2BB2XL U178 ( .B0(PCcur[24]), .B1(n21), .A0N(n18), .A1N(n130), .Y(n131)
         );
  NAND2X2 U179 ( .A(n132), .B(n131), .Y(n133) );
  AOI2BB2XL U180 ( .B0(PCcur[23]), .B1(n22), .A0N(n18), .A1N(n126), .Y(n127)
         );
  NAND2X2 U181 ( .A(n128), .B(n127), .Y(n129) );
  INVXL U182 ( .A(PCplus4_regD[8]), .Y(n66) );
  INVXL U183 ( .A(PCplus4_regD[6]), .Y(n58) );
  INVXL U184 ( .A(PCplus4_regD[4]), .Y(n50) );
  INVXL U185 ( .A(PCplus4_regD[5]), .Y(n54) );
  INVXL U186 ( .A(PCplus4_regD[3]), .Y(n46) );
  INVXL U187 ( .A(PCplus4_regD[2]), .Y(n40) );
  INVXL U188 ( .A(PCplus4_regD[7]), .Y(n62) );
  INVXL U189 ( .A(PCplus4_regD[9]), .Y(n70) );
  CLKINVX1 U190 ( .A(PCplus4[12]), .Y(n81) );
  INVXL U191 ( .A(PCplus4[4]), .Y(n53) );
  AOI2BB2X1 U192 ( .B0(PCcur[4]), .B1(n21), .A0N(n14), .A1N(n50), .Y(n52) );
  CLKINVX1 U193 ( .A(n117), .Y(n10) );
  BUFX12 U194 ( .A(n163), .Y(n14) );
  INVXL U195 ( .A(PCplus4[5]), .Y(n57) );
  AOI2BB2XL U196 ( .B0(PCcur[5]), .B1(n22), .A0N(n14), .A1N(n54), .Y(n56) );
  CLKINVX1 U197 ( .A(PCplus4[0]), .Y(n34) );
  AOI2BB2XL U198 ( .B0(PCcur[1]), .B1(n21), .A0N(n18), .A1N(n37), .Y(n38) );
  CLKINVX1 U199 ( .A(PCplus4[1]), .Y(n37) );
  INVXL U200 ( .A(PCplus4[20]), .Y(n114) );
  AOI2BB2XL U201 ( .B0(PCcur[14]), .B1(n22), .A0N(n18), .A1N(n89), .Y(n90) );
  AOI2BB2XL U202 ( .B0(PCcur[16]), .B1(n22), .A0N(n18), .A1N(n97), .Y(n98) );
  AOI2BB2XL U203 ( .B0(PCcur[11]), .B1(n22), .A0N(n18), .A1N(n77), .Y(n78) );
  AOI2BB2XL U204 ( .B0(PCcur[12]), .B1(n22), .A0N(n18), .A1N(n81), .Y(n82) );
  OAI211X1 U205 ( .A0(n18), .A1(n49), .B0(n48), .C0(n47), .Y(PCnext[3]) );
  AOI2BB2XL U206 ( .B0(PCcur[3]), .B1(n21), .A0N(n14), .A1N(n46), .Y(n48) );
  INVXL U207 ( .A(PCplus4[7]), .Y(n65) );
  INVXL U208 ( .A(PCplus4[9]), .Y(n73) );
  OAI211X1 U209 ( .A0(n18), .A1(n45), .B0(n44), .C0(n43), .Y(PCnext[2]) );
  CLKINVX1 U210 ( .A(PCplus4[2]), .Y(n45) );
  AOI2BB2XL U211 ( .B0(PCcur[2]), .B1(n21), .A0N(n14), .A1N(n40), .Y(n44) );
  OAI211X1 U212 ( .A0(n18), .A1(n61), .B0(n59), .C0(n60), .Y(PCnext[6]) );
  INVXL U213 ( .A(PCplus4[6]), .Y(n61) );
  INVX1 U214 ( .A(PCplus4[8]), .Y(n69) );
  AOI2BB2X1 U215 ( .B0(PCcur[8]), .B1(n22), .A0N(n14), .A1N(n66), .Y(n68) );
  NAND2XL U216 ( .A(PCcur[28]), .B(n21), .Y(n152) );
  NAND2X1 U217 ( .A(n136), .B(n135), .Y(n137) );
  NAND2X1 U218 ( .A(n146), .B(n145), .Y(n147) );
  NAND3X1 U219 ( .A(n160), .B(n159), .C(n158), .Y(n161) );
  NAND2XL U220 ( .A(PCcur[30]), .B(n21), .Y(n160) );
  NAND3X1 U221 ( .A(n168), .B(n167), .C(n166), .Y(n170) );
  NAND2XL U222 ( .A(PCcur[31]), .B(n21), .Y(n168) );
  AOI222XL U223 ( .A0(PCplus4[10]), .A1(n19), .B0(PCplus4_regD[10]), .B1(n143), 
        .C0(PCcur[10]), .C1(n21), .Y(n75) );
  MX2XL U224 ( .A(PCplus4_regD[0]), .B(PCplus4[0]), .S0(n7), .Y(
        PCplus4_actual[0]) );
  MX2XL U225 ( .A(PCplus4_regD[1]), .B(PCplus4[1]), .S0(n7), .Y(
        PCplus4_actual[1]) );
  NAND2BXL U226 ( .AN(n14), .B(PCplus4_regD[31]), .Y(n167) );
  NAND2BXL U227 ( .AN(n14), .B(PCplus4_regD[28]), .Y(n151) );
  NAND2BXL U228 ( .AN(n14), .B(PCplus4_regD[30]), .Y(n159) );
  NAND2BXL U229 ( .AN(n14), .B(PCplus4_regD[29]), .Y(n155) );
  AOI2BB2XL U230 ( .B0(PCcur[13]), .B1(n22), .A0N(n18), .A1N(n85), .Y(n86) );
  NAND2X1 U231 ( .A(n112), .B(n111), .Y(n113) );
  AOI2BB2XL U232 ( .B0(PCcur[19]), .B1(n21), .A0N(n18), .A1N(n110), .Y(n111)
         );
  AOI2BB2XL U233 ( .B0(PCcur[18]), .B1(n22), .A0N(n18), .A1N(n106), .Y(n107)
         );
  AOI2BB2XL U234 ( .B0(PCcur[17]), .B1(n22), .A0N(n18), .A1N(n101), .Y(n102)
         );
  AOI222XL U235 ( .A0(PCplus4_regD[17]), .A1(n143), .B0(targetAddr[15]), .B1(
        n16), .C0(JumpRegAddr[17]), .C1(n24), .Y(n103) );
  AOI2BB2XL U236 ( .B0(PCcur[15]), .B1(n22), .A0N(n18), .A1N(n93), .Y(n94) );
  AOI222XL U237 ( .A0(PCplus4_regD[15]), .A1(n143), .B0(targetAddr[13]), .B1(
        n17), .C0(JumpRegAddr[15]), .C1(n24), .Y(n95) );
  AO22X1 U238 ( .A0(targetAddr[8]), .A1(n16), .B0(JumpRegAddr[10]), .B1(n23), 
        .Y(n76) );
  AOI222XL U239 ( .A0(PCplus4_regD[12]), .A1(n143), .B0(targetAddr[10]), .B1(
        n17), .C0(JumpRegAddr[12]), .C1(n24), .Y(n83) );
  AOI222XL U240 ( .A0(PCplus4_regD[16]), .A1(n143), .B0(targetAddr[14]), .B1(
        n16), .C0(JumpRegAddr[16]), .C1(n24), .Y(n99) );
  AOI222XL U241 ( .A0(PCplus4_regD[11]), .A1(n143), .B0(targetAddr[9]), .B1(
        n17), .C0(JumpRegAddr[11]), .C1(n24), .Y(n79) );
  AOI222XL U242 ( .A0(PCplus4_regD[13]), .A1(n143), .B0(targetAddr[11]), .B1(
        n17), .C0(JumpRegAddr[13]), .C1(n24), .Y(n87) );
  AOI222XL U243 ( .A0(PCplus4_regD[14]), .A1(n143), .B0(targetAddr[12]), .B1(
        n17), .C0(JumpRegAddr[14]), .C1(n24), .Y(n91) );
  CLKMX2X4 U244 ( .A(PCplus4_regD[24]), .B(PCplus4[24]), .S0(n7), .Y(
        PCplus4_actual[24]) );
  CLKMX2X4 U245 ( .A(PCplus4_regD[23]), .B(PCplus4[23]), .S0(n7), .Y(
        PCplus4_actual[23]) );
  AOI2BB2X2 U246 ( .B0(PCcur[7]), .B1(n22), .A0N(n14), .A1N(n62), .Y(n64) );
  AOI2BB2X2 U247 ( .B0(PCcur[9]), .B1(n22), .A0N(n14), .A1N(n70), .Y(n72) );
  OA22X4 U248 ( .A0(ADDresult[18]), .A1(n109), .B0(n25), .B1(n109), .Y(
        PCnext[18]) );
  OA22X4 U249 ( .A0(ADDresult[21]), .A1(n121), .B0(n26), .B1(n121), .Y(
        PCnext[21]) );
  OA22X4 U250 ( .A0(ADDresult[23]), .A1(n129), .B0(n26), .B1(n129), .Y(
        PCnext[23]) );
  OA22X4 U251 ( .A0(ADDresult[24]), .A1(n133), .B0(n26), .B1(n133), .Y(
        PCnext[24]) );
endmodule


module PCsrcLogic ( pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, 
        predict, stallcache, stall_lw_use, PCsrc );
  output [2:0] PCsrc;
  input pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, predict,
         stallcache, stall_lw_use;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  INVX12 U3 ( .A(Jump), .Y(n10) );
  INVX3 U4 ( .A(n12), .Y(n2) );
  AND3XL U5 ( .A(predict), .B(Branch_IF), .C(n10), .Y(n11) );
  CLKMX2X6 U6 ( .A(n11), .B(equal), .S0(n1), .Y(n13) );
  AND2X8 U7 ( .A(pred_cond), .B(Branch_EX), .Y(n1) );
  OAI2BB1X4 U8 ( .A0N(n7), .A1N(n6), .B0(n2), .Y(PCsrc[0]) );
  INVXL U9 ( .A(JumpReg), .Y(n6) );
  NAND2X8 U10 ( .A(n4), .B(n5), .Y(n12) );
  INVX4 U11 ( .A(equal), .Y(n8) );
  MXI2X4 U12 ( .A(equal), .B(n10), .S0(n3), .Y(n9) );
  NAND2X2 U13 ( .A(pred_cond), .B(Branch_EX), .Y(n3) );
  MXI2X4 U14 ( .A(n10), .B(n8), .S0(n1), .Y(n7) );
  AOI2BB1X4 U15 ( .A0N(n13), .A1N(JumpReg), .B0(n12), .Y(PCsrc[2]) );
  CLKINVX12 U16 ( .A(stallcache), .Y(n4) );
  AOI2BB1X4 U17 ( .A0N(n9), .A1N(JumpReg), .B0(n12), .Y(PCsrc[1]) );
  CLKINVX1 U18 ( .A(stall_lw_use), .Y(n5) );
endmodule


module ALU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45,
         n46, n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93,
         n94, n96, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109,
         n110, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n127, n128, n129, n130, n131, n132, n134, n137, n138,
         n140, n141, n143, n144, n145, n146, n147, n148, n149, n150, n153,
         n154, n155, n156, n157, n158, n159, n161, n162, n163, n164, n165,
         n166, n167, n168, n173, n174, n175, n176, n177, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n195, n196, n197, n198, n199, n200, n202, n205, n206, n207, n208,
         n209, n211, n212, n213, n214, n215, n216, n217, n218, n221, n222,
         n223, n224, n225, n226, n227, n229, n231, n232, n233, n234, n235,
         n236, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n260, n261, n262, n263,
         n264, n265, n268, n269, n270, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n306, n307, n308, n309, n310, n312, n313, n314,
         n315, n316, n317, n319, n320, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438;

  XNOR2X4 U38 ( .A(n72), .B(n10), .Y(SUM[28]) );
  AOI21X4 U57 ( .A0(n94), .A1(n77), .B0(n78), .Y(n5) );
  OAI21X4 U105 ( .A0(n148), .A1(n113), .B0(n114), .Y(n3) );
  NAND2XL U357 ( .A(B[24]), .B(A[24]), .Y(n107) );
  NOR2XL U358 ( .A(B[24]), .B(A[24]), .Y(n106) );
  AOI21X4 U359 ( .A0(n426), .A1(n44), .B0(n45), .Y(n43) );
  XOR2X4 U360 ( .A(n428), .B(n424), .Y(SUM[21]) );
  CLKINVX20 U361 ( .A(n17), .Y(n424) );
  INVX1 U362 ( .A(n200), .Y(n202) );
  NAND2X1 U363 ( .A(n4), .B(n55), .Y(n53) );
  OAI21X1 U364 ( .A0(n96), .A1(n86), .B0(n89), .Y(n85) );
  AOI21X2 U365 ( .A0(n426), .A1(n84), .B0(n85), .Y(n83) );
  NOR2BX2 U366 ( .AN(n93), .B(n86), .Y(n84) );
  AOI21X2 U367 ( .A0(n426), .A1(n55), .B0(n56), .Y(n54) );
  AND2X6 U368 ( .A(n432), .B(n433), .Y(n173) );
  INVX2 U369 ( .A(B[17]), .Y(n432) );
  AOI21X2 U370 ( .A0(n426), .A1(n297), .B0(n105), .Y(n103) );
  BUFX4 U371 ( .A(n79), .Y(n435) );
  CLKINVX8 U372 ( .A(n59), .Y(n57) );
  NOR2X4 U373 ( .A(n68), .B(n61), .Y(n59) );
  NAND2X2 U374 ( .A(n4), .B(n44), .Y(n42) );
  NOR2X4 U375 ( .A(n6), .B(n46), .Y(n44) );
  BUFX3 U376 ( .A(n118), .Y(n425) );
  BUFX20 U377 ( .A(n3), .Y(n426) );
  INVX3 U378 ( .A(n426), .Y(n110) );
  CLKINVX4 U379 ( .A(n236), .Y(n234) );
  AOI21X4 U380 ( .A0(n236), .A1(n431), .B0(n229), .Y(n227) );
  OAI21X4 U381 ( .A0(n241), .A1(n245), .B0(n242), .Y(n236) );
  NAND2X8 U382 ( .A(n153), .B(n167), .Y(n147) );
  CLKINVX2 U383 ( .A(n167), .Y(n165) );
  NAND2X2 U384 ( .A(n167), .B(n303), .Y(n158) );
  NOR2X4 U385 ( .A(n176), .B(n173), .Y(n167) );
  NAND2X1 U386 ( .A(n4), .B(n93), .Y(n91) );
  INVX1 U387 ( .A(n6), .Y(n75) );
  AOI21X2 U388 ( .A0(n218), .A1(n199), .B0(n200), .Y(n198) );
  INVX8 U389 ( .A(n247), .Y(n246) );
  OAI21X2 U390 ( .A0(n437), .A1(n82), .B0(n83), .Y(n81) );
  NOR2X6 U391 ( .A(n212), .B(n205), .Y(n199) );
  INVX8 U392 ( .A(n205), .Y(n308) );
  NOR2X6 U393 ( .A(B[13]), .B(A[13]), .Y(n205) );
  XNOR2X4 U394 ( .A(n157), .B(n19), .Y(SUM[19]) );
  OAI21X1 U395 ( .A0(n5), .A1(n57), .B0(n58), .Y(n56) );
  NAND2X4 U396 ( .A(B[3]), .B(A[3]), .Y(n280) );
  XNOR2X4 U397 ( .A(n63), .B(n9), .Y(SUM[29]) );
  XNOR2X4 U398 ( .A(n146), .B(n18), .Y(SUM[20]) );
  BUFX6 U399 ( .A(n253), .Y(n427) );
  NOR2X8 U400 ( .A(B[22]), .B(A[22]), .Y(n124) );
  NOR2X2 U401 ( .A(n117), .B(n124), .Y(n115) );
  INVX4 U402 ( .A(n124), .Y(n299) );
  OAI21X2 U403 ( .A0(n134), .A1(n124), .B0(n127), .Y(n123) );
  AOI21X2 U404 ( .A0(n426), .A1(n93), .B0(n94), .Y(n92) );
  OAI21X4 U405 ( .A0(n268), .A1(n274), .B0(n269), .Y(n263) );
  NAND2X8 U406 ( .A(B[4]), .B(A[4]), .Y(n274) );
  NAND2X4 U407 ( .A(B[5]), .B(A[5]), .Y(n269) );
  NAND2X4 U408 ( .A(n306), .B(n186), .Y(n23) );
  NAND2X4 U409 ( .A(B[15]), .B(A[15]), .Y(n186) );
  NOR2X8 U410 ( .A(B[4]), .B(A[4]), .Y(n273) );
  NOR2X8 U411 ( .A(n273), .B(n268), .Y(n262) );
  NOR2X6 U412 ( .A(B[5]), .B(A[5]), .Y(n268) );
  NOR2X2 U413 ( .A(B[12]), .B(A[12]), .Y(n212) );
  OR2X4 U414 ( .A(B[30]), .B(A[30]), .Y(n429) );
  OAI21X1 U415 ( .A0(n5), .A1(n46), .B0(n47), .Y(n45) );
  NAND2X2 U416 ( .A(n59), .B(n429), .Y(n46) );
  AOI21X1 U417 ( .A0(n60), .A1(n429), .B0(n49), .Y(n47) );
  NAND2X4 U418 ( .A(B[16]), .B(A[16]), .Y(n177) );
  OAI21X4 U419 ( .A0(n173), .A1(n177), .B0(n174), .Y(n168) );
  AOI21X2 U420 ( .A0(n426), .A1(n66), .B0(n67), .Y(n65) );
  NAND2X2 U421 ( .A(n434), .B(n177), .Y(n22) );
  INVX1 U422 ( .A(n51), .Y(n49) );
  AOI21X4 U423 ( .A0(n236), .A1(n221), .B0(n222), .Y(n216) );
  AND2X8 U424 ( .A(n431), .B(n310), .Y(n221) );
  XNOR2X4 U425 ( .A(n119), .B(n15), .Y(SUM[23]) );
  XNOR2X4 U426 ( .A(n90), .B(n12), .Y(SUM[26]) );
  OAI21X4 U427 ( .A0(n205), .A1(n213), .B0(n206), .Y(n200) );
  NAND2X6 U428 ( .A(n308), .B(n206), .Y(n25) );
  NAND2X4 U429 ( .A(B[13]), .B(A[13]), .Y(n206) );
  OAI21X2 U430 ( .A0(n246), .A1(n188), .B0(n189), .Y(n187) );
  XOR2X4 U431 ( .A(n261), .B(n32), .Y(SUM[6]) );
  AOI21X2 U432 ( .A0(n275), .A1(n262), .B0(n263), .Y(n261) );
  NAND2X4 U433 ( .A(B[22]), .B(A[22]), .Y(n127) );
  AOI21X4 U434 ( .A0(n132), .A1(n115), .B0(n116), .Y(n114) );
  NAND2X1 U435 ( .A(B[14]), .B(A[14]), .Y(n195) );
  OAI21X1 U436 ( .A0(n437), .A1(n140), .B0(n141), .Y(n428) );
  NOR2X2 U437 ( .A(B[28]), .B(A[28]), .Y(n68) );
  OR2XL U438 ( .A(B[31]), .B(A[31]), .Y(n430) );
  NAND2X4 U439 ( .A(n199), .B(n183), .Y(n181) );
  INVX4 U440 ( .A(n213), .Y(n211) );
  NAND2X1 U441 ( .A(n309), .B(n213), .Y(n26) );
  NAND2X2 U442 ( .A(B[12]), .B(A[12]), .Y(n213) );
  INVX3 U443 ( .A(n148), .Y(n150) );
  INVX2 U444 ( .A(n163), .Y(n161) );
  NOR2X4 U445 ( .A(n137), .B(n144), .Y(n131) );
  INVX2 U446 ( .A(n147), .Y(n149) );
  NAND2X2 U447 ( .A(n310), .B(n224), .Y(n27) );
  OAI21X1 U448 ( .A0(n437), .A1(n73), .B0(n74), .Y(n72) );
  NAND2X4 U449 ( .A(n93), .B(n77), .Y(n6) );
  OAI21XL U450 ( .A0(n265), .A1(n257), .B0(n260), .Y(n256) );
  INVX3 U451 ( .A(n436), .Y(n279) );
  INVX3 U452 ( .A(n285), .Y(n284) );
  INVX3 U453 ( .A(n215), .Y(n217) );
  INVX3 U454 ( .A(n155), .Y(n302) );
  INVX1 U455 ( .A(n117), .Y(n298) );
  OR2X8 U456 ( .A(B[10]), .B(A[10]), .Y(n431) );
  NAND2X4 U457 ( .A(B[11]), .B(A[11]), .Y(n224) );
  AOI21X2 U458 ( .A0(n218), .A1(n309), .B0(n211), .Y(n209) );
  INVX4 U459 ( .A(n216), .Y(n218) );
  OAI21X4 U460 ( .A0(n286), .A1(n289), .B0(n287), .Y(n285) );
  NOR2X6 U461 ( .A(B[19]), .B(A[19]), .Y(n155) );
  NOR2X4 U462 ( .A(n155), .B(n162), .Y(n153) );
  AOI21X1 U463 ( .A0(n426), .A1(n75), .B0(n76), .Y(n74) );
  XOR2X4 U464 ( .A(n246), .B(n30), .Y(SUM[8]) );
  NAND2X4 U465 ( .A(B[28]), .B(A[28]), .Y(n71) );
  NAND2X1 U466 ( .A(B[17]), .B(A[17]), .Y(n174) );
  INVX1 U467 ( .A(n274), .Y(n272) );
  NAND2XL U468 ( .A(B[7]), .B(A[7]), .Y(n253) );
  OAI21X1 U469 ( .A0(n252), .A1(n260), .B0(n427), .Y(n251) );
  INVXL U470 ( .A(A[17]), .Y(n433) );
  XNOR2X4 U471 ( .A(n196), .B(n24), .Y(SUM[14]) );
  OAI21X1 U472 ( .A0(n246), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U473 ( .A0(n275), .A1(n255), .B0(n256), .Y(n254) );
  XNOR2X2 U474 ( .A(n128), .B(n16), .Y(SUM[22]) );
  OAI21X1 U475 ( .A0(n437), .A1(n129), .B0(n130), .Y(n128) );
  NAND2X2 U476 ( .A(n4), .B(n66), .Y(n64) );
  NOR2X2 U477 ( .A(n6), .B(n68), .Y(n66) );
  NOR2X2 U478 ( .A(B[6]), .B(A[6]), .Y(n257) );
  OR2XL U479 ( .A(B[16]), .B(A[16]), .Y(n434) );
  OAI21X1 U480 ( .A0(n5), .A1(n68), .B0(n71), .Y(n67) );
  OAI21X2 U481 ( .A0(n246), .A1(n226), .B0(n227), .Y(n225) );
  NOR2X4 U482 ( .A(B[14]), .B(A[14]), .Y(n192) );
  NOR2X2 U483 ( .A(B[18]), .B(A[18]), .Y(n162) );
  NAND2X2 U484 ( .A(B[18]), .B(A[18]), .Y(n163) );
  CLKAND2X2 U485 ( .A(n131), .B(n299), .Y(n122) );
  NOR2XL U486 ( .A(B[27]), .B(A[27]), .Y(n79) );
  OAI21X2 U487 ( .A0(n246), .A1(n244), .B0(n245), .Y(n243) );
  OAI21X1 U488 ( .A0(n246), .A1(n215), .B0(n216), .Y(n214) );
  OAI21X4 U489 ( .A0(n137), .A1(n145), .B0(n138), .Y(n132) );
  NAND2X1 U490 ( .A(B[21]), .B(A[21]), .Y(n138) );
  OAI21X1 U491 ( .A0(n437), .A1(n102), .B0(n103), .Y(n101) );
  AND2X4 U492 ( .A(n199), .B(n307), .Y(n190) );
  INVX1 U493 ( .A(n192), .Y(n307) );
  OAI21X1 U494 ( .A0(n437), .A1(n176), .B0(n177), .Y(n175) );
  BUFX20 U495 ( .A(n2), .Y(n437) );
  OR2X4 U496 ( .A(B[3]), .B(A[3]), .Y(n436) );
  OAI21X1 U497 ( .A0(n117), .A1(n127), .B0(n425), .Y(n116) );
  NOR2X2 U498 ( .A(B[23]), .B(A[23]), .Y(n117) );
  OAI21X1 U499 ( .A0(n155), .A1(n163), .B0(n156), .Y(n154) );
  INVX1 U500 ( .A(n223), .Y(n310) );
  OAI21X1 U501 ( .A0(n223), .A1(n231), .B0(n224), .Y(n222) );
  NAND2X1 U502 ( .A(B[10]), .B(A[10]), .Y(n231) );
  NOR2X2 U503 ( .A(B[11]), .B(A[11]), .Y(n223) );
  NOR2X4 U504 ( .A(n99), .B(n106), .Y(n93) );
  INVX1 U505 ( .A(n107), .Y(n105) );
  XNOR2X4 U506 ( .A(n207), .B(n25), .Y(SUM[13]) );
  OAI21X2 U507 ( .A0(n246), .A1(n208), .B0(n209), .Y(n207) );
  NAND2X2 U508 ( .A(B[9]), .B(A[9]), .Y(n242) );
  NOR2X2 U509 ( .A(B[2]), .B(A[2]), .Y(n282) );
  NAND2X2 U510 ( .A(B[2]), .B(A[2]), .Y(n283) );
  NAND2X2 U511 ( .A(B[25]), .B(A[25]), .Y(n100) );
  NOR2X4 U512 ( .A(B[25]), .B(A[25]), .Y(n99) );
  NOR2X2 U513 ( .A(B[7]), .B(A[7]), .Y(n252) );
  NOR2X2 U514 ( .A(n282), .B(n279), .Y(n277) );
  XNOR2X4 U515 ( .A(n232), .B(n28), .Y(SUM[10]) );
  OAI21X2 U516 ( .A0(n246), .A1(n233), .B0(n234), .Y(n232) );
  AOI21X4 U517 ( .A0(n247), .A1(n179), .B0(n180), .Y(n2) );
  NOR2X2 U518 ( .A(n215), .B(n181), .Y(n179) );
  NOR2X6 U519 ( .A(n438), .B(A[1]), .Y(n286) );
  XNOR2X4 U520 ( .A(n108), .B(n14), .Y(SUM[24]) );
  NOR2X2 U521 ( .A(n6), .B(n57), .Y(n55) );
  NOR2X8 U522 ( .A(n147), .B(n113), .Y(n4) );
  OAI21X2 U523 ( .A0(n279), .A1(n283), .B0(n280), .Y(n278) );
  OAI21X1 U524 ( .A0(n437), .A1(n147), .B0(n148), .Y(n146) );
  NAND2X2 U525 ( .A(n303), .B(n163), .Y(n20) );
  NAND2X1 U526 ( .A(B[19]), .B(A[19]), .Y(n156) );
  NOR2X2 U527 ( .A(B[9]), .B(A[9]), .Y(n241) );
  XNOR2X4 U528 ( .A(n187), .B(n23), .Y(SUM[15]) );
  XNOR2X2 U529 ( .A(n225), .B(n27), .Y(SUM[11]) );
  NAND2X4 U530 ( .A(B[20]), .B(A[20]), .Y(n145) );
  XNOR2X4 U531 ( .A(n52), .B(n8), .Y(SUM[30]) );
  OAI21X2 U532 ( .A0(n437), .A1(n53), .B0(n54), .Y(n52) );
  OAI21X2 U533 ( .A0(n437), .A1(n165), .B0(n166), .Y(n164) );
  NAND2X2 U534 ( .A(B[6]), .B(A[6]), .Y(n260) );
  NOR2X6 U535 ( .A(B[29]), .B(A[29]), .Y(n61) );
  OAI21X1 U536 ( .A0(n437), .A1(n42), .B0(n43), .Y(n41) );
  OAI21X4 U537 ( .A0(n61), .A1(n71), .B0(n62), .Y(n60) );
  NAND2X4 U538 ( .A(B[29]), .B(A[29]), .Y(n62) );
  INVX1 U539 ( .A(n268), .Y(n316) );
  OAI21X1 U540 ( .A0(n185), .A1(n195), .B0(n186), .Y(n184) );
  OAI21X2 U541 ( .A0(n437), .A1(n158), .B0(n159), .Y(n157) );
  OAI21X2 U542 ( .A0(n99), .A1(n107), .B0(n100), .Y(n94) );
  NOR2X2 U543 ( .A(n185), .B(n192), .Y(n183) );
  NOR2X4 U544 ( .A(B[15]), .B(A[15]), .Y(n185) );
  NAND2X6 U545 ( .A(n438), .B(A[1]), .Y(n287) );
  BUFX20 U546 ( .A(B[1]), .Y(n438) );
  INVX1 U547 ( .A(n241), .Y(n312) );
  NOR2X2 U548 ( .A(n244), .B(n241), .Y(n235) );
  XOR2X1 U549 ( .A(n437), .B(n22), .Y(SUM[16]) );
  NOR2X4 U550 ( .A(B[20]), .B(A[20]), .Y(n144) );
  NOR2X2 U551 ( .A(n252), .B(n257), .Y(n250) );
  XNOR2X4 U552 ( .A(n41), .B(n7), .Y(SUM[31]) );
  XNOR2X4 U553 ( .A(n101), .B(n13), .Y(SUM[25]) );
  OAI21X2 U554 ( .A0(n437), .A1(n91), .B0(n92), .Y(n90) );
  XOR2X2 U555 ( .A(n254), .B(n31), .Y(SUM[7]) );
  INVX1 U556 ( .A(n273), .Y(n317) );
  NAND2X4 U557 ( .A(n235), .B(n221), .Y(n215) );
  XNOR2X4 U558 ( .A(n175), .B(n21), .Y(SUM[17]) );
  NOR2X4 U559 ( .A(B[8]), .B(A[8]), .Y(n244) );
  NAND2X4 U560 ( .A(B[8]), .B(A[8]), .Y(n245) );
  XNOR2X4 U561 ( .A(n81), .B(n11), .Y(SUM[27]) );
  NAND2X1 U562 ( .A(n4), .B(n84), .Y(n82) );
  INVX1 U563 ( .A(n106), .Y(n297) );
  NAND2X2 U564 ( .A(B[0]), .B(A[0]), .Y(n289) );
  OAI21X1 U565 ( .A0(n437), .A1(n120), .B0(n121), .Y(n119) );
  NAND2XL U566 ( .A(n122), .B(n149), .Y(n120) );
  AOI21X4 U567 ( .A0(n168), .A1(n153), .B0(n154), .Y(n148) );
  OAI21X2 U568 ( .A0(n437), .A1(n109), .B0(n110), .Y(n108) );
  AOI21X4 U569 ( .A0(n285), .A1(n277), .B0(n278), .Y(n276) );
  OAI21X4 U570 ( .A0(n276), .A1(n248), .B0(n249), .Y(n247) );
  NAND2X1 U571 ( .A(n217), .B(n309), .Y(n208) );
  NAND2X4 U572 ( .A(n115), .B(n131), .Y(n113) );
  NAND2XL U573 ( .A(n190), .B(n217), .Y(n188) );
  XOR2X1 U574 ( .A(n284), .B(n36), .Y(SUM[2]) );
  INVXL U575 ( .A(n282), .Y(n319) );
  INVXL U576 ( .A(n244), .Y(n313) );
  INVXL U577 ( .A(n252), .Y(n314) );
  OAI21XL U578 ( .A0(n284), .A1(n282), .B0(n283), .Y(n281) );
  INVXL U579 ( .A(n286), .Y(n320) );
  NAND2XL U580 ( .A(n293), .B(n71), .Y(n10) );
  OAI21X2 U581 ( .A0(n216), .A1(n181), .B0(n182), .Y(n180) );
  INVX3 U582 ( .A(n276), .Y(n275) );
  INVXL U583 ( .A(n5), .Y(n76) );
  NAND2XL U584 ( .A(n149), .B(n131), .Y(n129) );
  INVXL U585 ( .A(n168), .Y(n166) );
  NAND2XL U586 ( .A(n235), .B(n431), .Y(n226) );
  NAND2XL U587 ( .A(n429), .B(n51), .Y(n8) );
  NAND2XL U588 ( .A(n4), .B(n75), .Y(n73) );
  NAND2X2 U589 ( .A(n262), .B(n250), .Y(n248) );
  AOI21X2 U590 ( .A0(n263), .A1(n250), .B0(n251), .Y(n249) );
  INVXL U591 ( .A(n4), .Y(n109) );
  NAND2XL U592 ( .A(n302), .B(n156), .Y(n19) );
  NAND2XL U593 ( .A(n301), .B(n145), .Y(n18) );
  INVXL U594 ( .A(n263), .Y(n265) );
  INVXL U595 ( .A(n185), .Y(n306) );
  XNOR2XL U596 ( .A(n275), .B(n34), .Y(SUM[4]) );
  NAND2XL U597 ( .A(n431), .B(n231), .Y(n28) );
  INVX1 U598 ( .A(n94), .Y(n96) );
  INVXL U599 ( .A(n132), .Y(n134) );
  XOR2XL U600 ( .A(n37), .B(n289), .Y(SUM[1]) );
  INVXL U601 ( .A(n212), .Y(n309) );
  NAND2BXL U602 ( .AN(n288), .B(n289), .Y(n38) );
  NOR2X1 U603 ( .A(B[16]), .B(A[16]), .Y(n176) );
  NAND2XL U604 ( .A(B[27]), .B(A[27]), .Y(n80) );
  NAND2XL U605 ( .A(B[30]), .B(A[30]), .Y(n51) );
  NAND2XL U606 ( .A(B[23]), .B(A[23]), .Y(n118) );
  CLKINVX1 U607 ( .A(n60), .Y(n58) );
  AOI21X1 U608 ( .A0(n150), .A1(n131), .B0(n132), .Y(n130) );
  NAND2XL U609 ( .A(n4), .B(n297), .Y(n102) );
  NAND2XL U610 ( .A(n217), .B(n199), .Y(n197) );
  NAND2XL U611 ( .A(n149), .B(n301), .Y(n140) );
  NAND2X1 U612 ( .A(n292), .B(n62), .Y(n9) );
  OAI21X1 U613 ( .A0(n437), .A1(n64), .B0(n65), .Y(n63) );
  CLKINVX1 U614 ( .A(n61), .Y(n292) );
  CLKINVX1 U615 ( .A(n68), .Y(n293) );
  OAI21X1 U616 ( .A0(n435), .A1(n89), .B0(n80), .Y(n78) );
  XNOR2X1 U617 ( .A(n214), .B(n26), .Y(SUM[12]) );
  CLKINVX1 U618 ( .A(n235), .Y(n233) );
  NAND2X1 U619 ( .A(n307), .B(n195), .Y(n24) );
  XNOR2X1 U620 ( .A(n281), .B(n35), .Y(SUM[3]) );
  NAND2X1 U621 ( .A(n436), .B(n280), .Y(n35) );
  NAND2X1 U622 ( .A(n317), .B(n274), .Y(n34) );
  NAND2X1 U623 ( .A(n304), .B(n174), .Y(n21) );
  CLKINVX1 U624 ( .A(n173), .Y(n304) );
  NAND2X1 U625 ( .A(n299), .B(n127), .Y(n16) );
  XNOR2X1 U626 ( .A(n164), .B(n20), .Y(SUM[18]) );
  NAND2X1 U627 ( .A(n294), .B(n80), .Y(n11) );
  INVXL U628 ( .A(n435), .Y(n294) );
  NAND2X1 U629 ( .A(n296), .B(n100), .Y(n13) );
  INVXL U630 ( .A(n99), .Y(n296) );
  NAND2X1 U631 ( .A(n300), .B(n138), .Y(n17) );
  INVXL U632 ( .A(n137), .Y(n300) );
  NAND2X1 U633 ( .A(n298), .B(n425), .Y(n15) );
  XNOR2X1 U634 ( .A(n243), .B(n29), .Y(SUM[9]) );
  NAND2X1 U635 ( .A(n312), .B(n242), .Y(n29) );
  NOR2X2 U636 ( .A(n435), .B(n86), .Y(n77) );
  CLKINVX1 U637 ( .A(n144), .Y(n301) );
  CLKINVX1 U638 ( .A(n162), .Y(n303) );
  NAND2X1 U639 ( .A(n314), .B(n427), .Y(n31) );
  AOI21X1 U640 ( .A0(n200), .A1(n183), .B0(n184), .Y(n182) );
  CLKINVX1 U641 ( .A(n231), .Y(n229) );
  AOI21X1 U642 ( .A0(n218), .A1(n190), .B0(n191), .Y(n189) );
  OAI21XL U643 ( .A0(n202), .A1(n192), .B0(n195), .Y(n191) );
  AOI21X1 U644 ( .A0(n150), .A1(n301), .B0(n143), .Y(n141) );
  CLKINVX1 U645 ( .A(n145), .Y(n143) );
  AOI21XL U646 ( .A0(n168), .A1(n303), .B0(n161), .Y(n159) );
  AOI21X1 U647 ( .A0(n150), .A1(n122), .B0(n123), .Y(n121) );
  NAND2XL U648 ( .A(n297), .B(n107), .Y(n14) );
  NAND2XL U649 ( .A(n295), .B(n89), .Y(n12) );
  INVXL U650 ( .A(n86), .Y(n295) );
  NOR2X1 U651 ( .A(n264), .B(n257), .Y(n255) );
  INVXL U652 ( .A(n262), .Y(n264) );
  NAND2X1 U653 ( .A(n320), .B(n287), .Y(n37) );
  XOR2X1 U654 ( .A(n270), .B(n33), .Y(SUM[5]) );
  NAND2XL U655 ( .A(n316), .B(n269), .Y(n33) );
  AOI21X1 U656 ( .A0(n275), .A1(n317), .B0(n272), .Y(n270) );
  NAND2X1 U657 ( .A(n319), .B(n283), .Y(n36) );
  NAND2XL U658 ( .A(n315), .B(n260), .Y(n32) );
  CLKINVX1 U659 ( .A(n257), .Y(n315) );
  NAND2X1 U660 ( .A(n313), .B(n245), .Y(n30) );
  NAND2X1 U661 ( .A(n430), .B(n40), .Y(n7) );
  NAND2XL U662 ( .A(B[31]), .B(A[31]), .Y(n40) );
  INVX1 U663 ( .A(n38), .Y(SUM[0]) );
  NAND2X1 U664 ( .A(B[26]), .B(A[26]), .Y(n89) );
  NOR2X2 U665 ( .A(B[26]), .B(A[26]), .Y(n86) );
  NOR2XL U666 ( .A(B[0]), .B(A[0]), .Y(n288) );
  NOR2X2 U667 ( .A(B[21]), .B(A[21]), .Y(n137) );
endmodule


module ALU_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90,
         n91, n92, n93, n94, n95, n98, n99, n100, n101, n102, n104, n105, n106,
         n107, n108, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n127, n128, n129, n130, n131, n132, n133, n136,
         n137, n138, n139, n140, n143, n144, n145, n146, n147, n148, n149,
         n152, n153, n154, n155, n156, n157, n158, n160, n161, n162, n163,
         n164, n165, n166, n167, n172, n173, n174, n175, n176, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n194, n195, n196, n197, n198, n199, n201, n204, n205, n206,
         n207, n208, n210, n211, n212, n214, n215, n216, n217, n220, n221,
         n222, n223, n224, n225, n226, n228, n229, n230, n231, n232, n233,
         n234, n235, n240, n241, n242, n243, n244, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n259, n260, n261, n262,
         n263, n264, n267, n269, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n290,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472;

  NAND2X2 U386 ( .A(n326), .B(A[24]), .Y(n106) );
  XNOR2X4 U387 ( .A(n231), .B(n28), .Y(DIFF[10]) );
  NOR2X6 U388 ( .A(n116), .B(n123), .Y(n114) );
  OAI21X2 U389 ( .A0(n116), .A1(n455), .B0(n117), .Y(n115) );
  INVX3 U390 ( .A(n116), .Y(n296) );
  NOR2X8 U391 ( .A(n327), .B(A[23]), .Y(n116) );
  XNOR2X2 U392 ( .A(n174), .B(n21), .Y(DIFF[17]) );
  XNOR2X2 U393 ( .A(n40), .B(n7), .Y(DIFF[31]) );
  AOI21X4 U394 ( .A0(n3), .A1(n83), .B0(n84), .Y(n82) );
  NOR2X2 U395 ( .A(n94), .B(n462), .Y(n83) );
  OAI21X4 U396 ( .A0(n60), .A1(n70), .B0(n61), .Y(n59) );
  NAND2X4 U397 ( .A(n290), .B(n61), .Y(n9) );
  NAND2X6 U398 ( .A(n321), .B(A[29]), .Y(n61) );
  OAI21X2 U399 ( .A0(n5), .A1(n45), .B0(n46), .Y(n44) );
  OAI21X2 U400 ( .A0(n466), .A1(n52), .B0(n53), .Y(n51) );
  OAI21X2 U401 ( .A0(n466), .A1(n119), .B0(n120), .Y(n118) );
  OAI21X2 U402 ( .A0(n466), .A1(n157), .B0(n158), .Y(n156) );
  OAI21X2 U403 ( .A0(n466), .A1(n146), .B0(n147), .Y(n145) );
  OAI21X2 U404 ( .A0(n466), .A1(n139), .B0(n140), .Y(n138) );
  OAI21X1 U405 ( .A0(n95), .A1(n462), .B0(n88), .Y(n84) );
  XNOR2X2 U406 ( .A(n51), .B(n8), .Y(DIFF[30]) );
  OAI21X2 U407 ( .A0(n278), .A1(n282), .B0(n279), .Y(n277) );
  XOR2X2 U408 ( .A(n453), .B(n30), .Y(DIFF[8]) );
  OAI21X2 U409 ( .A0(n453), .A1(n187), .B0(n188), .Y(n186) );
  XNOR2X4 U410 ( .A(n100), .B(n13), .Y(DIFF[25]) );
  INVX8 U411 ( .A(B[21]), .Y(n329) );
  NAND2X2 U412 ( .A(n331), .B(A[19]), .Y(n155) );
  INVX8 U413 ( .A(B[19]), .Y(n331) );
  INVX6 U414 ( .A(n147), .Y(n149) );
  NAND2X2 U415 ( .A(n4), .B(n54), .Y(n52) );
  AOI21X2 U416 ( .A0(n3), .A1(n54), .B0(n55), .Y(n53) );
  OAI21X2 U417 ( .A0(n133), .A1(n123), .B0(n455), .Y(n122) );
  INVX8 U418 ( .A(n123), .Y(n297) );
  NOR2X4 U419 ( .A(n132), .B(n123), .Y(n121) );
  NOR2X8 U420 ( .A(n328), .B(A[22]), .Y(n123) );
  INVX1 U421 ( .A(n4), .Y(n108) );
  NAND2X1 U422 ( .A(n4), .B(n295), .Y(n101) );
  INVX4 U423 ( .A(n278), .Y(n316) );
  NOR2X6 U424 ( .A(n470), .B(A[3]), .Y(n278) );
  INVX8 U425 ( .A(n275), .Y(n274) );
  OAI21X4 U426 ( .A0(n267), .A1(n273), .B0(n460), .Y(n262) );
  NAND2X4 U427 ( .A(n471), .B(A[4]), .Y(n273) );
  NOR2X6 U428 ( .A(n472), .B(A[5]), .Y(n267) );
  AOI21X2 U429 ( .A0(n274), .A1(n254), .B0(n255), .Y(n253) );
  NOR2X1 U430 ( .A(n263), .B(n256), .Y(n254) );
  OA21X4 U431 ( .A0(n275), .A1(n247), .B0(n248), .Y(n453) );
  NAND2X4 U432 ( .A(n261), .B(n249), .Y(n247) );
  AOI21X4 U433 ( .A0(n262), .A1(n249), .B0(n250), .Y(n248) );
  NAND2X4 U434 ( .A(n470), .B(A[3]), .Y(n279) );
  INVX8 U435 ( .A(B[28]), .Y(n322) );
  NAND2X2 U436 ( .A(n58), .B(n47), .Y(n45) );
  XNOR2X2 U437 ( .A(n145), .B(n18), .Y(DIFF[20]) );
  BUFX16 U438 ( .A(n287), .Y(n464) );
  NOR2X6 U439 ( .A(n467), .B(A[0]), .Y(n287) );
  CLKXOR2X2 U440 ( .A(n260), .B(n32), .Y(DIFF[6]) );
  XOR2X4 U441 ( .A(n253), .B(n31), .Y(DIFF[7]) );
  OAI21X2 U442 ( .A0(n453), .A1(n207), .B0(n208), .Y(n206) );
  NAND2X4 U443 ( .A(n328), .B(A[22]), .Y(n455) );
  INVX12 U444 ( .A(B[22]), .Y(n328) );
  XNOR2X2 U445 ( .A(n62), .B(n9), .Y(DIFF[29]) );
  NAND2X4 U446 ( .A(n332), .B(A[18]), .Y(n162) );
  CLKINVX8 U447 ( .A(B[18]), .Y(n332) );
  AOI21X2 U448 ( .A0(n3), .A1(n43), .B0(n44), .Y(n42) );
  NAND2X2 U449 ( .A(n4), .B(n43), .Y(n41) );
  NOR2X2 U450 ( .A(n6), .B(n45), .Y(n43) );
  INVX8 U451 ( .A(B[7]), .Y(n343) );
  XNOR2X2 U452 ( .A(n118), .B(n15), .Y(DIFF[23]) );
  NAND2X2 U453 ( .A(n189), .B(n216), .Y(n187) );
  INVX6 U454 ( .A(n214), .Y(n216) );
  OAI21X4 U455 ( .A0(n98), .A1(n106), .B0(n99), .Y(n93) );
  AOI21X4 U456 ( .A0(n93), .A1(n76), .B0(n77), .Y(n5) );
  NOR2X8 U457 ( .A(n457), .B(n462), .Y(n76) );
  OAI21X2 U458 ( .A0(n457), .A1(n88), .B0(n79), .Y(n77) );
  NAND2X6 U459 ( .A(n318), .B(n286), .Y(n37) );
  NAND2X6 U460 ( .A(n468), .B(A[1]), .Y(n286) );
  NOR2X4 U461 ( .A(n154), .B(n161), .Y(n152) );
  NOR2X4 U462 ( .A(n332), .B(A[18]), .Y(n161) );
  NOR2X8 U463 ( .A(n146), .B(n112), .Y(n4) );
  NAND2X2 U464 ( .A(n114), .B(n130), .Y(n112) );
  NAND2X8 U465 ( .A(n152), .B(n166), .Y(n146) );
  NOR2X8 U466 ( .A(n211), .B(n204), .Y(n198) );
  CLKINVX8 U467 ( .A(n211), .Y(n307) );
  NOR2X6 U468 ( .A(n338), .B(A[12]), .Y(n211) );
  OAI21X4 U469 ( .A0(n215), .A1(n180), .B0(n181), .Y(n179) );
  NOR2X4 U470 ( .A(n214), .B(n180), .Y(n178) );
  NAND2X2 U471 ( .A(n198), .B(n182), .Y(n180) );
  XNOR2X4 U472 ( .A(n89), .B(n12), .Y(DIFF[26]) );
  XNOR2X4 U473 ( .A(n107), .B(n14), .Y(DIFF[24]) );
  AOI21X4 U474 ( .A0(n167), .A1(n152), .B0(n153), .Y(n147) );
  OAI21X2 U475 ( .A0(n154), .A1(n162), .B0(n155), .Y(n153) );
  AOI21X2 U476 ( .A0(n3), .A1(n92), .B0(n93), .Y(n91) );
  INVX8 U477 ( .A(n458), .Y(n3) );
  XNOR2X4 U478 ( .A(n127), .B(n16), .Y(DIFF[22]) );
  OAI21X2 U479 ( .A0(n466), .A1(n128), .B0(n129), .Y(n127) );
  OAI21X4 U480 ( .A0(n204), .A1(n212), .B0(n205), .Y(n199) );
  CLKINVX8 U481 ( .A(n212), .Y(n210) );
  NAND2X2 U482 ( .A(n307), .B(n212), .Y(n26) );
  NAND2X4 U483 ( .A(n338), .B(A[12]), .Y(n212) );
  CLKINVX4 U484 ( .A(n199), .Y(n201) );
  AOI21X2 U485 ( .A0(n217), .A1(n198), .B0(n199), .Y(n197) );
  AOI21X2 U486 ( .A0(n199), .A1(n182), .B0(n183), .Y(n181) );
  OAI21X1 U487 ( .A0(n201), .A1(n191), .B0(n194), .Y(n190) );
  INVX6 U488 ( .A(n215), .Y(n217) );
  NAND2X1 U489 ( .A(n472), .B(A[5]), .Y(n460) );
  NOR2X2 U490 ( .A(n339), .B(A[11]), .Y(n222) );
  NOR2X4 U491 ( .A(n344), .B(A[6]), .Y(n256) );
  NAND2X2 U492 ( .A(n334), .B(A[16]), .Y(n176) );
  NOR2X2 U493 ( .A(n281), .B(n278), .Y(n276) );
  NOR2BX2 U494 ( .AN(n74), .B(n56), .Y(n54) );
  CLKINVX6 U495 ( .A(B[4]), .Y(n471) );
  OAI2BB1X2 U496 ( .A0N(n75), .A1N(n58), .B0(n57), .Y(n55) );
  OAI21X2 U497 ( .A0(n453), .A1(n225), .B0(n226), .Y(n224) );
  XNOR2X2 U498 ( .A(n138), .B(n17), .Y(DIFF[21]) );
  INVX3 U499 ( .A(B[30]), .Y(n320) );
  CLKINVX6 U500 ( .A(B[6]), .Y(n344) );
  CLKINVX6 U501 ( .A(B[25]), .Y(n325) );
  CLKINVX6 U502 ( .A(B[12]), .Y(n338) );
  CLKINVX6 U503 ( .A(B[11]), .Y(n339) );
  INVX4 U504 ( .A(B[13]), .Y(n337) );
  INVX3 U505 ( .A(B[3]), .Y(n470) );
  INVX3 U506 ( .A(B[17]), .Y(n333) );
  INVX3 U507 ( .A(n146), .Y(n148) );
  NOR2X4 U508 ( .A(n336), .B(A[14]), .Y(n191) );
  CLKINVX6 U509 ( .A(n459), .Y(n172) );
  AOI21X4 U510 ( .A0(n246), .A1(n178), .B0(n179), .Y(n2) );
  OAI21X2 U511 ( .A0(n453), .A1(n243), .B0(n244), .Y(n242) );
  OAI21X2 U512 ( .A0(n453), .A1(n196), .B0(n197), .Y(n195) );
  OA21X4 U513 ( .A0(n453), .A1(n214), .B0(n215), .Y(n454) );
  OAI21X2 U514 ( .A0(n453), .A1(n232), .B0(n233), .Y(n231) );
  XOR2X4 U515 ( .A(n454), .B(n26), .Y(DIFF[12]) );
  NOR2X1 U516 ( .A(n471), .B(A[4]), .Y(n272) );
  INVX1 U517 ( .A(n273), .Y(n271) );
  INVX1 U518 ( .A(n272), .Y(n315) );
  NOR2X1 U519 ( .A(n343), .B(A[7]), .Y(n251) );
  XNOR2X2 U520 ( .A(n80), .B(n11), .Y(DIFF[27]) );
  OAI21X2 U521 ( .A0(n466), .A1(n81), .B0(n82), .Y(n80) );
  OAI21X4 U522 ( .A0(n172), .A1(n176), .B0(n173), .Y(n167) );
  OAI21X1 U523 ( .A0(n5), .A1(n67), .B0(n70), .Y(n66) );
  NOR2X6 U524 ( .A(n342), .B(A[8]), .Y(n243) );
  CLKINVX4 U525 ( .A(B[8]), .Y(n342) );
  NAND2X2 U526 ( .A(n330), .B(A[20]), .Y(n144) );
  INVX16 U527 ( .A(B[20]), .Y(n330) );
  NAND2X2 U528 ( .A(n339), .B(A[11]), .Y(n223) );
  NAND2X2 U529 ( .A(n323), .B(A[27]), .Y(n79) );
  CLKINVX4 U530 ( .A(B[27]), .Y(n323) );
  NOR2X2 U531 ( .A(n337), .B(A[13]), .Y(n204) );
  NAND2X2 U532 ( .A(n328), .B(A[22]), .Y(n456) );
  NAND2X4 U533 ( .A(n76), .B(n92), .Y(n6) );
  CLKINVX2 U534 ( .A(n6), .Y(n74) );
  NOR2X2 U535 ( .A(n331), .B(A[19]), .Y(n154) );
  NAND2X2 U536 ( .A(n333), .B(A[17]), .Y(n173) );
  NAND2X4 U537 ( .A(n327), .B(A[23]), .Y(n117) );
  INVX4 U538 ( .A(B[23]), .Y(n327) );
  INVX1 U539 ( .A(n5), .Y(n75) );
  INVXL U540 ( .A(n58), .Y(n56) );
  NOR2X4 U541 ( .A(n67), .B(n60), .Y(n58) );
  XNOR2X4 U542 ( .A(n195), .B(n24), .Y(DIFF[14]) );
  XNOR2X2 U543 ( .A(n206), .B(n25), .Y(DIFF[13]) );
  NOR2X4 U544 ( .A(n98), .B(n463), .Y(n92) );
  NOR2X6 U545 ( .A(n325), .B(A[25]), .Y(n98) );
  NAND2X6 U546 ( .A(n469), .B(A[2]), .Y(n282) );
  BUFX8 U547 ( .A(n78), .Y(n457) );
  NOR2X1 U548 ( .A(n324), .B(A[26]), .Y(n85) );
  OA21X4 U549 ( .A0(n147), .A1(n112), .B0(n113), .Y(n458) );
  OR2X8 U550 ( .A(n333), .B(A[17]), .Y(n459) );
  XNOR2X2 U551 ( .A(n242), .B(n29), .Y(DIFF[9]) );
  CLKINVX3 U552 ( .A(B[5]), .Y(n472) );
  CLKAND2X2 U553 ( .A(n330), .B(A[20]), .Y(n461) );
  INVX3 U554 ( .A(B[14]), .Y(n336) );
  BUFX8 U555 ( .A(n85), .Y(n462) );
  BUFX4 U556 ( .A(n105), .Y(n463) );
  OR2XL U557 ( .A(n469), .B(A[2]), .Y(n465) );
  CLKINVX8 U558 ( .A(B[2]), .Y(n469) );
  NAND2X1 U559 ( .A(n324), .B(A[26]), .Y(n88) );
  CLKINVX6 U560 ( .A(B[26]), .Y(n324) );
  INVX1 U561 ( .A(n222), .Y(n308) );
  NOR2X2 U562 ( .A(n229), .B(n222), .Y(n220) );
  NOR2X1 U563 ( .A(n323), .B(A[27]), .Y(n78) );
  INVX1 U564 ( .A(n463), .Y(n295) );
  NOR2X1 U565 ( .A(n334), .B(A[16]), .Y(n175) );
  INVX8 U566 ( .A(B[0]), .Y(n467) );
  NOR2X1 U567 ( .A(n469), .B(A[2]), .Y(n281) );
  NOR2X1 U568 ( .A(n340), .B(A[10]), .Y(n229) );
  NAND2X2 U569 ( .A(n340), .B(A[10]), .Y(n230) );
  NAND2X2 U570 ( .A(n325), .B(A[25]), .Y(n99) );
  AOI21X1 U571 ( .A0(n3), .A1(n74), .B0(n75), .Y(n73) );
  OAI21X2 U572 ( .A0(n466), .A1(n72), .B0(n73), .Y(n71) );
  BUFX20 U573 ( .A(n2), .Y(n466) );
  NAND2X4 U574 ( .A(n344), .B(A[6]), .Y(n259) );
  XNOR2X4 U575 ( .A(n186), .B(n23), .Y(DIFF[15]) );
  OAI21X4 U576 ( .A0(n285), .A1(n464), .B0(n286), .Y(n284) );
  NAND2X2 U577 ( .A(n329), .B(A[21]), .Y(n137) );
  OAI21X2 U578 ( .A0(n466), .A1(n164), .B0(n165), .Y(n163) );
  NAND2X6 U579 ( .A(n342), .B(A[8]), .Y(n244) );
  OAI21X1 U580 ( .A0(n184), .A1(n194), .B0(n185), .Y(n183) );
  NAND2X2 U581 ( .A(n336), .B(A[14]), .Y(n194) );
  NOR2X2 U582 ( .A(n184), .B(n191), .Y(n182) );
  OAI21X2 U583 ( .A0(n466), .A1(n63), .B0(n64), .Y(n62) );
  NOR2X4 U584 ( .A(n335), .B(A[15]), .Y(n184) );
  CLKINVX6 U585 ( .A(B[15]), .Y(n335) );
  NOR2X1 U586 ( .A(n320), .B(A[30]), .Y(n49) );
  OAI21X2 U587 ( .A0(n466), .A1(n41), .B0(n42), .Y(n40) );
  OAI21X1 U588 ( .A0(n466), .A1(n175), .B0(n176), .Y(n174) );
  AOI21X4 U589 ( .A0(n235), .A1(n220), .B0(n221), .Y(n215) );
  CLKINVX8 U590 ( .A(B[10]), .Y(n340) );
  NOR2X6 U591 ( .A(n468), .B(A[1]), .Y(n285) );
  CLKINVX12 U592 ( .A(B[1]), .Y(n468) );
  NOR2X2 U593 ( .A(n272), .B(n267), .Y(n261) );
  NOR2X4 U594 ( .A(n321), .B(A[29]), .Y(n60) );
  CLKINVX6 U595 ( .A(B[29]), .Y(n321) );
  INVX1 U596 ( .A(n243), .Y(n311) );
  NAND2XL U597 ( .A(n234), .B(n309), .Y(n225) );
  NAND2X4 U598 ( .A(n234), .B(n220), .Y(n214) );
  NOR2X4 U599 ( .A(n243), .B(n240), .Y(n234) );
  XNOR2X2 U600 ( .A(n156), .B(n19), .Y(DIFF[19]) );
  NAND2X4 U601 ( .A(n322), .B(A[28]), .Y(n70) );
  OAI21X2 U602 ( .A0(n466), .A1(n90), .B0(n91), .Y(n89) );
  NOR2X2 U603 ( .A(n330), .B(A[20]), .Y(n143) );
  CLKINVX6 U604 ( .A(B[24]), .Y(n326) );
  OAI21X2 U605 ( .A0(n466), .A1(n101), .B0(n102), .Y(n100) );
  AOI21X1 U606 ( .A0(n3), .A1(n295), .B0(n104), .Y(n102) );
  OAI21X2 U607 ( .A0(n466), .A1(n108), .B0(n458), .Y(n107) );
  AOI21X4 U608 ( .A0(n284), .A1(n276), .B0(n277), .Y(n275) );
  NAND2XL U609 ( .A(n216), .B(n307), .Y(n207) );
  NOR2X4 U610 ( .A(n136), .B(n143), .Y(n130) );
  OAI21X4 U611 ( .A0(n240), .A1(n244), .B0(n241), .Y(n235) );
  AOI21X1 U612 ( .A0(n131), .A1(n114), .B0(n115), .Y(n113) );
  CLKINVX1 U613 ( .A(B[9]), .Y(n341) );
  NOR2BX1 U614 ( .AN(n198), .B(n191), .Y(n189) );
  OAI21X2 U615 ( .A0(n136), .A1(n144), .B0(n137), .Y(n131) );
  INVXL U616 ( .A(n166), .Y(n164) );
  NAND2XL U617 ( .A(n294), .B(n99), .Y(n13) );
  NAND2XL U618 ( .A(n292), .B(n79), .Y(n11) );
  NOR2X2 U619 ( .A(n251), .B(n256), .Y(n249) );
  INVXL U620 ( .A(n131), .Y(n133) );
  INVXL U621 ( .A(n167), .Y(n165) );
  AOI21X1 U622 ( .A0(n3), .A1(n65), .B0(n66), .Y(n64) );
  NOR2X1 U623 ( .A(n6), .B(n67), .Y(n65) );
  NAND2XL U624 ( .A(n293), .B(n88), .Y(n12) );
  OAI21X1 U625 ( .A0(n222), .A1(n230), .B0(n223), .Y(n221) );
  NAND2XL U626 ( .A(n309), .B(n230), .Y(n28) );
  NAND2XL U627 ( .A(n301), .B(n162), .Y(n20) );
  OAI21X4 U628 ( .A0(n275), .A1(n247), .B0(n248), .Y(n246) );
  NAND2XL U629 ( .A(n304), .B(n185), .Y(n23) );
  NAND2XL U630 ( .A(n295), .B(n106), .Y(n14) );
  NAND2XL U631 ( .A(n299), .B(n144), .Y(n18) );
  OAI21X1 U632 ( .A0(n251), .A1(n259), .B0(n252), .Y(n250) );
  INVXL U633 ( .A(n262), .Y(n264) );
  NOR2X4 U634 ( .A(n175), .B(n172), .Y(n166) );
  NAND2XL U635 ( .A(n311), .B(n244), .Y(n30) );
  XOR2XL U636 ( .A(n466), .B(n22), .Y(DIFF[16]) );
  INVXL U637 ( .A(n462), .Y(n293) );
  NAND2XL U638 ( .A(n47), .B(n50), .Y(n8) );
  NOR2X1 U639 ( .A(n322), .B(A[28]), .Y(n67) );
  NOR2XL U640 ( .A(n326), .B(A[24]), .Y(n105) );
  NAND2XL U641 ( .A(n343), .B(A[7]), .Y(n252) );
  CLKINVX3 U642 ( .A(B[16]), .Y(n334) );
  NAND2XL U643 ( .A(n320), .B(A[30]), .Y(n50) );
  NAND2BX1 U644 ( .AN(n38), .B(n39), .Y(n7) );
  NAND2X1 U645 ( .A(n4), .B(n74), .Y(n72) );
  CLKINVX1 U646 ( .A(n59), .Y(n57) );
  XNOR2X1 U647 ( .A(n71), .B(n10), .Y(DIFF[28]) );
  NAND2XL U648 ( .A(n4), .B(n92), .Y(n90) );
  NAND2X1 U649 ( .A(n148), .B(n130), .Y(n128) );
  AOI21X1 U650 ( .A0(n149), .A1(n130), .B0(n131), .Y(n129) );
  NAND2XL U651 ( .A(n216), .B(n198), .Y(n196) );
  CLKINVX1 U652 ( .A(n92), .Y(n94) );
  CLKINVX1 U653 ( .A(n130), .Y(n132) );
  CLKINVX1 U654 ( .A(n235), .Y(n233) );
  NAND2X1 U655 ( .A(n166), .B(n301), .Y(n157) );
  CLKINVX1 U656 ( .A(n284), .Y(n283) );
  AOI21X1 U657 ( .A0(n59), .A1(n47), .B0(n48), .Y(n46) );
  CLKINVX1 U658 ( .A(n50), .Y(n48) );
  NAND2XL U659 ( .A(n4), .B(n65), .Y(n63) );
  NAND2BX1 U660 ( .AN(n67), .B(n70), .Y(n10) );
  NAND2X1 U661 ( .A(n297), .B(n456), .Y(n16) );
  NAND2X1 U662 ( .A(n298), .B(n137), .Y(n17) );
  NAND2X1 U663 ( .A(n296), .B(n117), .Y(n15) );
  INVXL U664 ( .A(n93), .Y(n95) );
  OAI21XL U665 ( .A0(n264), .A1(n256), .B0(n259), .Y(n255) );
  INVXL U666 ( .A(n261), .Y(n263) );
  CLKINVX1 U667 ( .A(n229), .Y(n309) );
  CLKINVX1 U668 ( .A(n161), .Y(n301) );
  CLKINVX1 U669 ( .A(n143), .Y(n299) );
  AOI21XL U670 ( .A0(n274), .A1(n261), .B0(n262), .Y(n260) );
  NAND2XL U671 ( .A(n313), .B(n259), .Y(n32) );
  INVXL U672 ( .A(n256), .Y(n313) );
  NAND2XL U673 ( .A(n306), .B(n205), .Y(n25) );
  INVXL U674 ( .A(n204), .Y(n306) );
  XNOR2X1 U675 ( .A(n224), .B(n27), .Y(DIFF[11]) );
  NAND2XL U676 ( .A(n308), .B(n223), .Y(n27) );
  INVXL U677 ( .A(n184), .Y(n304) );
  NAND2XL U678 ( .A(n310), .B(n241), .Y(n29) );
  INVXL U679 ( .A(n240), .Y(n310) );
  INVXL U680 ( .A(n234), .Y(n232) );
  NAND2X1 U681 ( .A(n305), .B(n194), .Y(n24) );
  INVXL U682 ( .A(n191), .Y(n305) );
  XNOR2X1 U683 ( .A(n163), .B(n20), .Y(DIFF[18]) );
  NAND2X1 U684 ( .A(n459), .B(n173), .Y(n21) );
  AOI21X1 U685 ( .A0(n217), .A1(n307), .B0(n210), .Y(n208) );
  NAND2X1 U686 ( .A(n312), .B(n252), .Y(n31) );
  INVXL U687 ( .A(n251), .Y(n312) );
  INVXL U688 ( .A(n136), .Y(n298) );
  AOI21XL U689 ( .A0(n235), .A1(n309), .B0(n228), .Y(n226) );
  CLKINVX1 U690 ( .A(n230), .Y(n228) );
  AOI21XL U691 ( .A0(n167), .A1(n301), .B0(n160), .Y(n158) );
  CLKINVX1 U692 ( .A(n162), .Y(n160) );
  AOI21X1 U693 ( .A0(n217), .A1(n189), .B0(n190), .Y(n188) );
  NAND2X1 U694 ( .A(n4), .B(n83), .Y(n81) );
  NAND2XL U695 ( .A(n300), .B(n155), .Y(n19) );
  INVXL U696 ( .A(n154), .Y(n300) );
  NAND2X1 U697 ( .A(n148), .B(n299), .Y(n139) );
  AOI21X1 U698 ( .A0(n149), .A1(n299), .B0(n461), .Y(n140) );
  CLKINVX1 U699 ( .A(n106), .Y(n104) );
  NAND2X1 U700 ( .A(n121), .B(n148), .Y(n119) );
  AOI21X1 U701 ( .A0(n149), .A1(n121), .B0(n122), .Y(n120) );
  XOR2X1 U702 ( .A(n269), .B(n33), .Y(DIFF[5]) );
  NAND2XL U703 ( .A(n314), .B(n460), .Y(n33) );
  AOI21X1 U704 ( .A0(n274), .A1(n315), .B0(n271), .Y(n269) );
  INVXL U705 ( .A(n267), .Y(n314) );
  NAND2X1 U706 ( .A(n303), .B(n176), .Y(n22) );
  INVXL U707 ( .A(n175), .Y(n303) );
  XNOR2XL U708 ( .A(n274), .B(n34), .Y(DIFF[4]) );
  NAND2X1 U709 ( .A(n315), .B(n273), .Y(n34) );
  INVXL U710 ( .A(n98), .Y(n294) );
  INVXL U711 ( .A(n457), .Y(n292) );
  XNOR2X1 U712 ( .A(n280), .B(n35), .Y(DIFF[3]) );
  NAND2X1 U713 ( .A(n316), .B(n279), .Y(n35) );
  OAI21XL U714 ( .A0(n283), .A1(n281), .B0(n282), .Y(n280) );
  CLKINVX1 U715 ( .A(n60), .Y(n290) );
  XOR2X1 U716 ( .A(n37), .B(n464), .Y(DIFF[1]) );
  CLKINVX1 U717 ( .A(n285), .Y(n318) );
  XOR2X1 U718 ( .A(n283), .B(n36), .Y(DIFF[2]) );
  NAND2X1 U719 ( .A(n465), .B(n282), .Y(n36) );
  CLKINVX1 U720 ( .A(n49), .Y(n47) );
  INVXL U721 ( .A(B[31]), .Y(n319) );
  NAND2XL U722 ( .A(n319), .B(A[31]), .Y(n39) );
  NOR2XL U723 ( .A(n319), .B(A[31]), .Y(n38) );
  NAND2XL U724 ( .A(n337), .B(A[13]), .Y(n205) );
  XNOR2XL U725 ( .A(n467), .B(A[0]), .Y(DIFF[0]) );
  NAND2XL U726 ( .A(n335), .B(A[15]), .Y(n185) );
  NOR2X2 U727 ( .A(n341), .B(A[9]), .Y(n240) );
  NAND2X1 U728 ( .A(n341), .B(A[9]), .Y(n241) );
  NOR2X2 U729 ( .A(n329), .B(A[21]), .Y(n136) );
endmodule


module ALU_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n1379, n1380, n1381, n1382,
         n1383, n1384;

  OAI21X1 U764 ( .A0(n45), .A1(n48), .B0(n46), .Y(n44) );
  NOR2X2 U765 ( .A(B[9]), .B(n129), .Y(n90) );
  CLKINVX2 U766 ( .A(A[9]), .Y(n129) );
  OAI21X2 U767 ( .A0(n90), .A1(n93), .B0(n91), .Y(n89) );
  NOR2X1 U768 ( .A(n92), .B(n90), .Y(n88) );
  OAI21X1 U769 ( .A0(n70), .A1(n73), .B0(n71), .Y(n69) );
  AOI21X4 U770 ( .A0(n34), .A1(n3), .B0(n4), .Y(n2) );
  OAI21X2 U771 ( .A0(n50), .A1(n35), .B0(n36), .Y(n34) );
  CLKINVX8 U772 ( .A(A[22]), .Y(n142) );
  NOR2X1 U773 ( .A(B[22]), .B(n142), .Y(n41) );
  NOR2X2 U774 ( .A(n1383), .B(n124), .Y(n107) );
  NAND2X2 U775 ( .A(n1383), .B(n124), .Y(n108) );
  CLKINVX2 U776 ( .A(A[4]), .Y(n124) );
  OAI21X4 U777 ( .A0(n63), .A1(n1), .B0(n2), .Y(GE_LT_GT_LE) );
  AOI21X2 U778 ( .A0(n94), .A1(n64), .B0(n65), .Y(n63) );
  NOR2X2 U779 ( .A(B[11]), .B(n131), .Y(n84) );
  CLKINVX1 U780 ( .A(A[11]), .Y(n131) );
  OAI21X1 U781 ( .A0(n84), .A1(n87), .B0(n85), .Y(n83) );
  NOR2X2 U782 ( .A(B[29]), .B(n149), .Y(n15) );
  INVX4 U783 ( .A(A[29]), .Y(n149) );
  NAND2X4 U784 ( .A(n13), .B(n7), .Y(n5) );
  NOR2X2 U785 ( .A(n9), .B(n11), .Y(n7) );
  NOR2X1 U786 ( .A(B[15]), .B(n135), .Y(n70) );
  NOR2X2 U787 ( .A(n70), .B(n72), .Y(n68) );
  OAI21X1 U788 ( .A0(n53), .A1(n56), .B0(n54), .Y(n52) );
  NOR2X4 U789 ( .A(n53), .B(n55), .Y(n51) );
  NOR2X1 U790 ( .A(B[19]), .B(n139), .Y(n53) );
  NOR2X1 U791 ( .A(B[26]), .B(n146), .Y(n25) );
  NAND2X2 U792 ( .A(B[26]), .B(n146), .Y(n26) );
  CLKINVX6 U793 ( .A(A[26]), .Y(n146) );
  NAND2X2 U794 ( .A(n3), .B(n33), .Y(n1) );
  NOR2X2 U795 ( .A(n5), .B(n19), .Y(n3) );
  INVX8 U796 ( .A(A[13]), .Y(n133) );
  CLKINVX4 U797 ( .A(A[30]), .Y(n150) );
  OAI21XL U798 ( .A0(n15), .A1(n18), .B0(n16), .Y(n14) );
  INVX1 U799 ( .A(A[7]), .Y(n127) );
  CLKINVX2 U800 ( .A(A[6]), .Y(n126) );
  BUFX3 U801 ( .A(n151), .Y(n1379) );
  INVX1 U802 ( .A(A[2]), .Y(n122) );
  CLKINVX6 U803 ( .A(A[14]), .Y(n134) );
  NOR2X4 U804 ( .A(B[23]), .B(n143), .Y(n39) );
  INVX6 U805 ( .A(A[23]), .Y(n143) );
  OAI21X1 U806 ( .A0(n59), .A1(n62), .B0(n60), .Y(n58) );
  NAND2X1 U807 ( .A(B[16]), .B(n136), .Y(n62) );
  NOR2X2 U808 ( .A(n80), .B(n66), .Y(n64) );
  NAND2X1 U809 ( .A(n88), .B(n82), .Y(n80) );
  NAND2X2 U810 ( .A(n74), .B(n68), .Y(n66) );
  CLKINVX2 U811 ( .A(A[27]), .Y(n147) );
  CLKINVX3 U812 ( .A(A[10]), .Y(n130) );
  CLKINVX6 U813 ( .A(A[25]), .Y(n145) );
  OAI21X1 U814 ( .A0(n81), .A1(n66), .B0(n67), .Y(n65) );
  NOR2X1 U815 ( .A(n1381), .B(n122), .Y(n114) );
  NAND2X1 U816 ( .A(n1380), .B(n121), .Y(n118) );
  NOR2XL U817 ( .A(B[21]), .B(n141), .Y(n45) );
  NOR2X1 U818 ( .A(n29), .B(n31), .Y(n27) );
  OAI21X1 U819 ( .A0(n20), .A1(n5), .B0(n6), .Y(n4) );
  OAI21X1 U820 ( .A0(n29), .A1(n32), .B0(n30), .Y(n28) );
  OAI21X1 U821 ( .A0(n117), .A1(n119), .B0(n118), .Y(n116) );
  OAI21X1 U822 ( .A0(n109), .A1(n95), .B0(n96), .Y(n94) );
  OAI21X1 U823 ( .A0(n112), .A1(n115), .B0(n113), .Y(n111) );
  NAND2XL U824 ( .A(n1382), .B(n123), .Y(n113) );
  OAI21X1 U825 ( .A0(n105), .A1(n108), .B0(n106), .Y(n104) );
  NOR2XL U826 ( .A(B[24]), .B(n144), .Y(n31) );
  NOR2X1 U827 ( .A(B[31]), .B(n1379), .Y(n9) );
  NAND2XL U828 ( .A(B[31]), .B(n1379), .Y(n10) );
  NOR2XL U829 ( .A(B[17]), .B(n137), .Y(n59) );
  INVXL U830 ( .A(A[31]), .Y(n151) );
  INVXL U831 ( .A(A[24]), .Y(n144) );
  OAI21XL U832 ( .A0(n76), .A1(n79), .B0(n77), .Y(n75) );
  INVXL U833 ( .A(A[21]), .Y(n141) );
  INVXL U834 ( .A(A[3]), .Y(n123) );
  INVXL U835 ( .A(A[1]), .Y(n121) );
  INVXL U836 ( .A(A[16]), .Y(n136) );
  INVXL U837 ( .A(A[18]), .Y(n138) );
  INVXL U838 ( .A(A[20]), .Y(n140) );
  AOI21X1 U839 ( .A0(n28), .A1(n21), .B0(n22), .Y(n20) );
  AOI21X1 U840 ( .A0(n14), .A1(n7), .B0(n8), .Y(n6) );
  NOR2X1 U841 ( .A(n1384), .B(n125), .Y(n105) );
  NAND2XL U842 ( .A(n1384), .B(n125), .Y(n106) );
  NOR2X1 U843 ( .A(n1380), .B(n121), .Y(n117) );
  NAND2X1 U844 ( .A(B[0]), .B(n120), .Y(n119) );
  AOI21X1 U845 ( .A0(n116), .A1(n110), .B0(n111), .Y(n109) );
  NAND2X1 U846 ( .A(n103), .B(n97), .Y(n95) );
  AOI21X1 U847 ( .A0(n104), .A1(n97), .B0(n98), .Y(n96) );
  AOI21X1 U848 ( .A0(n44), .A1(n37), .B0(n38), .Y(n36) );
  AOI21X1 U849 ( .A0(n58), .A1(n51), .B0(n52), .Y(n50) );
  OAI21XL U850 ( .A0(n39), .A1(n42), .B0(n40), .Y(n38) );
  AOI21X1 U851 ( .A0(n89), .A1(n82), .B0(n83), .Y(n81) );
  AOI21X1 U852 ( .A0(n75), .A1(n68), .B0(n69), .Y(n67) );
  NOR2X1 U853 ( .A(n107), .B(n105), .Y(n103) );
  NAND2X1 U854 ( .A(n1381), .B(n122), .Y(n115) );
  NOR2X1 U855 ( .A(n1382), .B(n123), .Y(n112) );
  NOR2X1 U856 ( .A(n114), .B(n112), .Y(n110) );
  CLKBUFX3 U857 ( .A(B[4]), .Y(n1383) );
  CLKBUFX3 U858 ( .A(B[2]), .Y(n1381) );
  CLKBUFX3 U859 ( .A(B[3]), .Y(n1382) );
  CLKBUFX3 U860 ( .A(B[1]), .Y(n1380) );
  CLKBUFX3 U861 ( .A(B[5]), .Y(n1384) );
  NAND2XL U862 ( .A(B[29]), .B(n149), .Y(n16) );
  NAND2XL U863 ( .A(B[28]), .B(n148), .Y(n18) );
  NAND2X1 U864 ( .A(n27), .B(n21), .Y(n19) );
  INVXL U865 ( .A(A[28]), .Y(n148) );
  NOR2X1 U866 ( .A(n17), .B(n15), .Y(n13) );
  NOR2X1 U867 ( .A(B[28]), .B(n148), .Y(n17) );
  NOR2XL U868 ( .A(B[13]), .B(n133), .Y(n76) );
  NAND2XL U869 ( .A(B[13]), .B(n133), .Y(n77) );
  NAND2XL U870 ( .A(B[12]), .B(n132), .Y(n79) );
  NAND2XL U871 ( .A(B[18]), .B(n138), .Y(n56) );
  NAND2XL U872 ( .A(B[19]), .B(n139), .Y(n54) );
  NAND2XL U873 ( .A(B[14]), .B(n134), .Y(n73) );
  NAND2XL U874 ( .A(B[15]), .B(n135), .Y(n71) );
  NAND2XL U875 ( .A(B[20]), .B(n140), .Y(n48) );
  NAND2XL U876 ( .A(B[21]), .B(n141), .Y(n46) );
  NOR2XL U877 ( .A(B[18]), .B(n138), .Y(n55) );
  NOR2XL U878 ( .A(B[14]), .B(n134), .Y(n72) );
  OAI21XL U879 ( .A0(n99), .A1(n102), .B0(n100), .Y(n98) );
  NAND2XL U880 ( .A(B[7]), .B(n127), .Y(n100) );
  NAND2XL U881 ( .A(B[6]), .B(n126), .Y(n102) );
  OAI21XL U882 ( .A0(n23), .A1(n26), .B0(n24), .Y(n22) );
  NAND2XL U883 ( .A(B[27]), .B(n147), .Y(n24) );
  NOR2X1 U884 ( .A(n23), .B(n25), .Y(n21) );
  NOR2X1 U885 ( .A(n99), .B(n101), .Y(n97) );
  NOR2XL U886 ( .A(B[6]), .B(n126), .Y(n101) );
  NOR2X1 U887 ( .A(n39), .B(n41), .Y(n37) );
  NOR2X1 U888 ( .A(n86), .B(n84), .Y(n82) );
  NOR2XL U889 ( .A(B[10]), .B(n130), .Y(n86) );
  NOR2X1 U890 ( .A(n78), .B(n76), .Y(n74) );
  NOR2XL U891 ( .A(B[12]), .B(n132), .Y(n78) );
  NAND2X1 U892 ( .A(n37), .B(n43), .Y(n35) );
  NOR2X1 U893 ( .A(n45), .B(n47), .Y(n43) );
  NOR2XL U894 ( .A(B[20]), .B(n140), .Y(n47) );
  NOR2XL U895 ( .A(B[8]), .B(n128), .Y(n92) );
  NOR2X1 U896 ( .A(n49), .B(n35), .Y(n33) );
  NAND2X1 U897 ( .A(n51), .B(n57), .Y(n49) );
  NOR2X1 U898 ( .A(n61), .B(n59), .Y(n57) );
  NOR2XL U899 ( .A(B[16]), .B(n136), .Y(n61) );
  NOR2X1 U900 ( .A(B[7]), .B(n127), .Y(n99) );
  NOR2X1 U901 ( .A(B[25]), .B(n145), .Y(n29) );
  NOR2X1 U902 ( .A(B[27]), .B(n147), .Y(n23) );
  NAND2XL U903 ( .A(B[17]), .B(n137), .Y(n60) );
  NAND2XL U904 ( .A(B[11]), .B(n131), .Y(n85) );
  NAND2XL U905 ( .A(B[10]), .B(n130), .Y(n87) );
  OAI21XL U906 ( .A0(n9), .A1(n12), .B0(n10), .Y(n8) );
  NAND2XL U907 ( .A(B[30]), .B(n150), .Y(n12) );
  NAND2XL U908 ( .A(B[8]), .B(n128), .Y(n93) );
  NAND2XL U909 ( .A(B[24]), .B(n144), .Y(n32) );
  NAND2XL U910 ( .A(B[22]), .B(n142), .Y(n42) );
  NOR2XL U911 ( .A(B[30]), .B(n150), .Y(n11) );
  NAND2XL U912 ( .A(B[9]), .B(n129), .Y(n91) );
  NAND2XL U913 ( .A(B[23]), .B(n143), .Y(n40) );
  NAND2XL U914 ( .A(B[25]), .B(n145), .Y(n30) );
  CLKINVX1 U915 ( .A(A[17]), .Y(n137) );
  CLKINVX1 U916 ( .A(A[8]), .Y(n128) );
  INVXL U917 ( .A(A[12]), .Y(n132) );
  INVXL U918 ( .A(A[19]), .Y(n139) );
  INVXL U919 ( .A(A[0]), .Y(n120) );
  INVXL U920 ( .A(A[5]), .Y(n125) );
  INVXL U921 ( .A(A[15]), .Y(n135) );
endmodule


module ALU_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346;

  MXI2X4 U255 ( .A(n112), .B(n108), .S0(n337), .Y(n80) );
  MXI2X1 U256 ( .A(n116), .B(n112), .S0(n338), .Y(n84) );
  MXI2X4 U257 ( .A(n144), .B(n142), .S0(n335), .Y(n112) );
  MXI2X4 U258 ( .A(n109), .B(n105), .S0(n337), .Y(n77) );
  MXI2X4 U259 ( .A(n105), .B(n101), .S0(n337), .Y(n73) );
  NAND2BX4 U260 ( .AN(n346), .B(n73), .Y(n41) );
  NOR2BX4 U261 ( .AN(n35), .B(n328), .Y(B[31]) );
  NAND2BX2 U262 ( .AN(n344), .B(n96), .Y(n64) );
  NOR2BX4 U263 ( .AN(n25), .B(n328), .Y(B[21]) );
  MXI2X2 U264 ( .A(n57), .B(n41), .S0(n342), .Y(n25) );
  CLKAND2X6 U265 ( .A(n28), .B(n322), .Y(B[24]) );
  CLKINVX2 U266 ( .A(n3), .Y(n322) );
  MXI2X2 U267 ( .A(n63), .B(n47), .S0(n340), .Y(n31) );
  NAND2BX2 U268 ( .AN(n344), .B(n95), .Y(n63) );
  NOR2BX2 U269 ( .AN(n9), .B(n329), .Y(B[5]) );
  MXI2X2 U270 ( .A(n162), .B(n160), .S0(n334), .Y(n130) );
  MXI2X1 U271 ( .A(n194), .B(n193), .S0(n332), .Y(n162) );
  MXI2X2 U272 ( .A(n130), .B(n126), .S0(n338), .Y(n98) );
  NOR2BX4 U273 ( .AN(n7), .B(n329), .Y(B[3]) );
  NAND2BX2 U274 ( .AN(n344), .B(n93), .Y(n61) );
  OR2X8 U275 ( .A(n219), .B(n220), .Y(n207) );
  OR2X4 U276 ( .A(SH[30]), .B(SH[26]), .Y(n219) );
  NOR2BX4 U277 ( .AN(n20), .B(n330), .Y(B[16]) );
  NOR2BX4 U278 ( .AN(n21), .B(n330), .Y(B[17]) );
  NOR2BX4 U279 ( .AN(n22), .B(n330), .Y(B[18]) );
  NOR2BX4 U280 ( .AN(n23), .B(n330), .Y(B[19]) );
  NOR2BX4 U281 ( .AN(n19), .B(n330), .Y(B[15]) );
  BUFX3 U282 ( .A(n3), .Y(n330) );
  MXI2X4 U283 ( .A(n169), .B(n168), .S0(n331), .Y(n137) );
  NAND2BX4 U284 ( .AN(n345), .B(n79), .Y(n47) );
  MXI2X4 U285 ( .A(n108), .B(n104), .S0(n337), .Y(n76) );
  NOR2BX4 U286 ( .AN(n12), .B(n328), .Y(B[8]) );
  OR2X4 U287 ( .A(n217), .B(n218), .Y(n206) );
  OR2X1 U288 ( .A(SH[24]), .B(SH[14]), .Y(n218) );
  MXI2X2 U289 ( .A(n321), .B(n125), .S0(n338), .Y(n97) );
  NAND2BX4 U290 ( .AN(n345), .B(n76), .Y(n44) );
  CLKBUFX20 U291 ( .A(SH[3]), .Y(n339) );
  MXI2X2 U292 ( .A(n163), .B(n161), .S0(n334), .Y(n131) );
  MXI2X2 U293 ( .A(n195), .B(n194), .S0(n332), .Y(n163) );
  NAND2BX4 U294 ( .AN(n345), .B(n77), .Y(n45) );
  NOR2BX4 U295 ( .AN(n33), .B(n328), .Y(B[29]) );
  NOR2BX4 U296 ( .AN(n8), .B(n329), .Y(B[4]) );
  NOR2BX4 U297 ( .AN(n30), .B(n328), .Y(B[26]) );
  MXI2X4 U298 ( .A(n185), .B(n184), .S0(n332), .Y(n153) );
  MXI2X4 U299 ( .A(n107), .B(n103), .S0(n337), .Y(n75) );
  NOR2BX4 U300 ( .AN(n11), .B(n329), .Y(B[7]) );
  MXI2X4 U301 ( .A(n171), .B(n170), .S0(n331), .Y(n139) );
  NAND2BX4 U302 ( .AN(n339), .B(A[6]), .Y(n170) );
  NOR2X4 U303 ( .A(n101), .B(n337), .Y(n69) );
  NAND2BX4 U304 ( .AN(n336), .B(n133), .Y(n101) );
  MXI2X2 U305 ( .A(n53), .B(n37), .S0(n342), .Y(n21) );
  NAND2BX4 U306 ( .AN(n346), .B(n69), .Y(n37) );
  NOR2X2 U307 ( .A(n102), .B(n337), .Y(n70) );
  NAND2BX4 U308 ( .AN(n345), .B(n75), .Y(n43) );
  NAND2BX2 U309 ( .AN(n344), .B(n90), .Y(n58) );
  MXI2X2 U310 ( .A(n122), .B(n118), .S0(n338), .Y(n90) );
  NOR2BX4 U311 ( .AN(n26), .B(n328), .Y(B[22]) );
  MXI2X2 U312 ( .A(n58), .B(n42), .S0(n342), .Y(n26) );
  MXI2X4 U313 ( .A(n114), .B(n110), .S0(n337), .Y(n82) );
  MXI2X4 U314 ( .A(n142), .B(n140), .S0(n335), .Y(n110) );
  NOR2BX4 U315 ( .AN(n13), .B(n328), .Y(B[9]) );
  MXI2X2 U316 ( .A(n54), .B(n38), .S0(n342), .Y(n22) );
  OR2X4 U317 ( .A(SH[12]), .B(SH[28]), .Y(n212) );
  NAND2BX2 U318 ( .AN(n344), .B(n92), .Y(n60) );
  MXI2X2 U319 ( .A(n124), .B(n120), .S0(n338), .Y(n92) );
  OR2X8 U320 ( .A(n215), .B(n216), .Y(n205) );
  OR2X2 U321 ( .A(SH[13]), .B(SH[29]), .Y(n215) );
  MXI2X4 U322 ( .A(n106), .B(n102), .S0(n337), .Y(n74) );
  MXI2X4 U323 ( .A(n134), .B(n132), .S0(n336), .Y(n102) );
  NAND2BX4 U324 ( .AN(n345), .B(n74), .Y(n42) );
  NAND2BX4 U325 ( .AN(n339), .B(A[3]), .Y(n167) );
  NAND2BX4 U326 ( .AN(n346), .B(n72), .Y(n40) );
  MXI2X4 U327 ( .A(n104), .B(n100), .S0(n337), .Y(n72) );
  MXI2X2 U328 ( .A(A[27]), .B(A[19]), .S0(n339), .Y(n191) );
  MXI2X4 U329 ( .A(n170), .B(n169), .S0(n331), .Y(n138) );
  INVXL U330 ( .A(A[1]), .Y(n324) );
  CLKINVX1 U331 ( .A(A[0]), .Y(n325) );
  INVX3 U332 ( .A(A[5]), .Y(n327) );
  MXI2X2 U333 ( .A(n161), .B(n159), .S0(n334), .Y(n321) );
  NOR2BX2 U334 ( .AN(n14), .B(n329), .Y(B[10]) );
  MXI2X4 U335 ( .A(n323), .B(n326), .S0(n331), .Y(n144) );
  BUFX6 U336 ( .A(n175), .Y(n326) );
  MXI2X4 U337 ( .A(n153), .B(n151), .S0(n334), .Y(n121) );
  NOR2BX2 U338 ( .AN(n6), .B(n329), .Y(B[2]) );
  NAND2BX2 U339 ( .AN(n339), .B(A[7]), .Y(n171) );
  NOR2BX4 U340 ( .AN(n31), .B(n328), .Y(B[27]) );
  AND2X4 U341 ( .A(n24), .B(n322), .Y(B[20]) );
  CLKBUFX6 U342 ( .A(n176), .Y(n323) );
  MXI2X2 U343 ( .A(A[12]), .B(A[4]), .S0(SH[3]), .Y(n176) );
  MXI2X2 U344 ( .A(A[14]), .B(A[6]), .S0(SH[3]), .Y(n178) );
  MXI2X2 U345 ( .A(A[19]), .B(A[11]), .S0(SH[3]), .Y(n183) );
  MXI2X2 U346 ( .A(n186), .B(n185), .S0(n332), .Y(n154) );
  MXI2X2 U347 ( .A(n115), .B(n111), .S0(n338), .Y(n83) );
  MXI2X4 U348 ( .A(n147), .B(n145), .S0(n335), .Y(n115) );
  NOR2BX2 U349 ( .AN(n34), .B(n328), .Y(B[30]) );
  MXI2X1 U350 ( .A(n66), .B(n50), .S0(n340), .Y(n34) );
  OR2X8 U351 ( .A(n339), .B(n324), .Y(n165) );
  NAND2BX4 U352 ( .AN(n345), .B(n81), .Y(n49) );
  MXI2X4 U353 ( .A(n113), .B(n109), .S0(n337), .Y(n81) );
  OR2X8 U354 ( .A(n339), .B(n325), .Y(n164) );
  MXI2X4 U355 ( .A(n179), .B(n178), .S0(n332), .Y(n147) );
  MXI2X4 U356 ( .A(n178), .B(n177), .S0(n331), .Y(n146) );
  MXI2X4 U357 ( .A(n326), .B(n174), .S0(n331), .Y(n143) );
  MXI2X4 U358 ( .A(n174), .B(n173), .S0(n331), .Y(n142) );
  MXI2X2 U359 ( .A(A[10]), .B(A[2]), .S0(SH[3]), .Y(n174) );
  MXI2X2 U360 ( .A(A[13]), .B(A[5]), .S0(SH[3]), .Y(n177) );
  MXI2X1 U361 ( .A(n118), .B(n114), .S0(n338), .Y(n86) );
  MXI2X4 U362 ( .A(n146), .B(n144), .S0(n335), .Y(n114) );
  NAND2BX2 U363 ( .AN(n345), .B(n85), .Y(n53) );
  MXI2X1 U364 ( .A(n117), .B(n113), .S0(n338), .Y(n85) );
  NOR2X4 U365 ( .A(n164), .B(n331), .Y(n132) );
  NAND2BX2 U366 ( .AN(n344), .B(n88), .Y(n56) );
  NAND2BX2 U367 ( .AN(n344), .B(n98), .Y(n66) );
  NAND2BX2 U368 ( .AN(n344), .B(n99), .Y(n67) );
  NAND2BX2 U369 ( .AN(n344), .B(n91), .Y(n59) );
  NAND2BX2 U370 ( .AN(n344), .B(n89), .Y(n57) );
  NAND2BX2 U371 ( .AN(n344), .B(n97), .Y(n65) );
  BUFX16 U372 ( .A(n343), .Y(n344) );
  NOR2BX4 U373 ( .AN(n29), .B(n328), .Y(B[25]) );
  MXI2X2 U374 ( .A(n61), .B(n45), .S0(n342), .Y(n29) );
  MXI2X4 U375 ( .A(n173), .B(n172), .S0(n331), .Y(n141) );
  MXI2X2 U376 ( .A(A[9]), .B(A[1]), .S0(SH[3]), .Y(n173) );
  MXI2X2 U377 ( .A(A[18]), .B(A[10]), .S0(SH[3]), .Y(n182) );
  MXI2X2 U378 ( .A(n160), .B(n158), .S0(n334), .Y(n128) );
  MXI2X2 U379 ( .A(n192), .B(n191), .S0(n332), .Y(n160) );
  MXI2X4 U380 ( .A(A[16]), .B(A[8]), .S0(SH[3]), .Y(n180) );
  MXI2X1 U381 ( .A(n121), .B(n117), .S0(n338), .Y(n89) );
  MXI2X4 U382 ( .A(n136), .B(n134), .S0(n336), .Y(n104) );
  MXI2X4 U383 ( .A(n166), .B(n165), .S0(n331), .Y(n134) );
  OR2X8 U384 ( .A(n339), .B(n327), .Y(n169) );
  MXI2X4 U385 ( .A(n158), .B(n156), .S0(n334), .Y(n126) );
  MXI2X2 U386 ( .A(n190), .B(n189), .S0(n332), .Y(n158) );
  OR2X2 U387 ( .A(SH[21]), .B(SH[19]), .Y(n211) );
  BUFX20 U388 ( .A(n3), .Y(n328) );
  MXI2X1 U389 ( .A(A[24]), .B(A[16]), .S0(SH[3]), .Y(n188) );
  MXI2X4 U390 ( .A(A[30]), .B(A[22]), .S0(n339), .Y(n194) );
  MXI2X2 U391 ( .A(n131), .B(n127), .S0(n338), .Y(n99) );
  MXI2X4 U392 ( .A(n159), .B(n157), .S0(n334), .Y(n127) );
  MXI2X4 U393 ( .A(n157), .B(n155), .S0(n334), .Y(n125) );
  MXI2X2 U394 ( .A(n189), .B(n188), .S0(n332), .Y(n157) );
  BUFX20 U395 ( .A(n3), .Y(n329) );
  NOR2X4 U396 ( .A(n103), .B(n337), .Y(n71) );
  MXI2X4 U397 ( .A(n135), .B(n133), .S0(n336), .Y(n103) );
  NAND2BX4 U398 ( .AN(n346), .B(n71), .Y(n39) );
  MXI2X4 U399 ( .A(n165), .B(n164), .S0(n331), .Y(n133) );
  MXI2X1 U400 ( .A(A[11]), .B(A[3]), .S0(SH[3]), .Y(n175) );
  MXI2X2 U401 ( .A(n183), .B(n182), .S0(n332), .Y(n151) );
  OR2X4 U402 ( .A(SH[22]), .B(SH[20]), .Y(n220) );
  MXI2X2 U403 ( .A(n177), .B(n176), .S0(n331), .Y(n145) );
  MXI2X4 U404 ( .A(n152), .B(n150), .S0(n334), .Y(n120) );
  MXI2X4 U405 ( .A(n182), .B(n181), .S0(n332), .Y(n150) );
  MXI2X2 U406 ( .A(A[17]), .B(A[9]), .S0(SH[3]), .Y(n181) );
  MXI2X2 U407 ( .A(n145), .B(n143), .S0(n335), .Y(n113) );
  MXI2XL U408 ( .A(A[31]), .B(A[23]), .S0(n339), .Y(n195) );
  MXI2X4 U409 ( .A(n140), .B(n138), .S0(n335), .Y(n108) );
  NAND2BX2 U410 ( .AN(n345), .B(n84), .Y(n52) );
  MXI2X2 U411 ( .A(n148), .B(n146), .S0(n335), .Y(n116) );
  MXI2X2 U412 ( .A(n55), .B(n39), .S0(n342), .Y(n23) );
  MXI2X1 U413 ( .A(n119), .B(n115), .S0(n338), .Y(n87) );
  MXI2X4 U414 ( .A(n141), .B(n139), .S0(n335), .Y(n109) );
  MXI2X4 U415 ( .A(n139), .B(n137), .S0(n336), .Y(n107) );
  MXI2X1 U416 ( .A(n65), .B(n49), .S0(n340), .Y(n33) );
  MXI2X4 U417 ( .A(n137), .B(n135), .S0(n336), .Y(n105) );
  BUFX12 U418 ( .A(n333), .Y(n336) );
  MXI2X4 U419 ( .A(n167), .B(n166), .S0(n331), .Y(n135) );
  NAND2BX1 U420 ( .AN(n339), .B(A[2]), .Y(n166) );
  NAND2BX2 U421 ( .AN(n346), .B(n70), .Y(n38) );
  MXI2X2 U422 ( .A(n126), .B(n122), .S0(n338), .Y(n94) );
  MXI2X4 U423 ( .A(n154), .B(n152), .S0(n334), .Y(n122) );
  MXI2X1 U424 ( .A(A[21]), .B(A[13]), .S0(SH[3]), .Y(n185) );
  MXI2X4 U425 ( .A(n155), .B(n153), .S0(n334), .Y(n123) );
  MXI2X1 U426 ( .A(n127), .B(n123), .S0(n338), .Y(n95) );
  MXI2X2 U427 ( .A(n111), .B(n107), .S0(n337), .Y(n79) );
  NOR2X4 U428 ( .A(n100), .B(n337), .Y(n68) );
  NAND2BX2 U429 ( .AN(n336), .B(n132), .Y(n100) );
  MXI2X2 U430 ( .A(n187), .B(n186), .S0(n332), .Y(n155) );
  MXI2X2 U431 ( .A(n188), .B(n187), .S0(n332), .Y(n156) );
  MXI2X4 U432 ( .A(n156), .B(n154), .S0(n334), .Y(n124) );
  MXI2X2 U433 ( .A(n60), .B(n44), .S0(n342), .Y(n28) );
  MXI2X1 U434 ( .A(A[23]), .B(A[15]), .S0(SH[3]), .Y(n187) );
  MXI2X4 U435 ( .A(n168), .B(n167), .S0(n331), .Y(n136) );
  NAND2BX4 U436 ( .AN(n339), .B(A[4]), .Y(n168) );
  NAND2BX2 U437 ( .AN(n345), .B(n78), .Y(n46) );
  MXI2X2 U438 ( .A(n110), .B(n106), .S0(n337), .Y(n78) );
  MXI2X2 U439 ( .A(n138), .B(n136), .S0(n336), .Y(n106) );
  BUFX20 U440 ( .A(SH[2]), .Y(n337) );
  MXI2X4 U441 ( .A(n180), .B(n179), .S0(n332), .Y(n148) );
  MXI2X4 U442 ( .A(A[15]), .B(A[7]), .S0(SH[3]), .Y(n179) );
  MXI2X4 U443 ( .A(n193), .B(n192), .S0(n332), .Y(n161) );
  MXI2X2 U444 ( .A(A[29]), .B(A[21]), .S0(n339), .Y(n193) );
  MXI2X4 U445 ( .A(A[28]), .B(A[20]), .S0(n339), .Y(n192) );
  MXI2X4 U446 ( .A(n191), .B(n190), .S0(n332), .Y(n159) );
  MXI2X2 U447 ( .A(A[26]), .B(A[18]), .S0(n339), .Y(n190) );
  MXI2X2 U448 ( .A(n149), .B(n147), .S0(n335), .Y(n117) );
  MXI2X2 U449 ( .A(n151), .B(n149), .S0(n335), .Y(n119) );
  MXI2X2 U450 ( .A(n181), .B(n180), .S0(n332), .Y(n149) );
  MXI2X1 U451 ( .A(A[25]), .B(A[17]), .S0(SH[3]), .Y(n189) );
  MXI2X2 U452 ( .A(n150), .B(n148), .S0(n335), .Y(n118) );
  NAND2BX2 U453 ( .AN(n345), .B(n83), .Y(n51) );
  MXI2X4 U454 ( .A(n184), .B(n183), .S0(n332), .Y(n152) );
  MXI2X2 U455 ( .A(A[20]), .B(A[12]), .S0(n339), .Y(n184) );
  NAND2BX2 U456 ( .AN(n345), .B(n82), .Y(n50) );
  CLKBUFX2 U457 ( .A(SH[4]), .Y(n340) );
  MXI2X2 U458 ( .A(n143), .B(n141), .S0(n335), .Y(n111) );
  MXI2X1 U459 ( .A(n62), .B(n46), .S0(n342), .Y(n30) );
  NAND2BX2 U460 ( .AN(n344), .B(n94), .Y(n62) );
  MXI2X1 U461 ( .A(n59), .B(n43), .S0(n342), .Y(n27) );
  MXI2X1 U462 ( .A(n123), .B(n119), .S0(n338), .Y(n91) );
  BUFX20 U463 ( .A(SH[1]), .Y(n334) );
  MXI2X4 U464 ( .A(n172), .B(n171), .S0(n331), .Y(n140) );
  MXI2X2 U465 ( .A(n64), .B(n48), .S0(n340), .Y(n32) );
  NAND2BX2 U466 ( .AN(n345), .B(n80), .Y(n48) );
  NOR2BX1 U467 ( .AN(n32), .B(n328), .Y(B[28]) );
  BUFX20 U468 ( .A(SH[0]), .Y(n332) );
  BUFX20 U469 ( .A(SH[0]), .Y(n331) );
  MXI2X2 U470 ( .A(A[8]), .B(A[0]), .S0(SH[3]), .Y(n172) );
  BUFX8 U471 ( .A(n343), .Y(n345) );
  BUFX12 U472 ( .A(SH[2]), .Y(n338) );
  BUFX8 U473 ( .A(SH[1]), .Y(n335) );
  BUFX12 U474 ( .A(SH[4]), .Y(n342) );
  CLKBUFX3 U475 ( .A(SH[4]), .Y(n341) );
  NOR2X1 U476 ( .A(n36), .B(n341), .Y(n4) );
  MXI2X1 U477 ( .A(n128), .B(n124), .S0(n338), .Y(n96) );
  NOR2BX1 U478 ( .AN(n27), .B(n328), .Y(B[23]) );
  OR2X8 U479 ( .A(n197), .B(n198), .Y(n3) );
  OR2X8 U480 ( .A(n201), .B(n202), .Y(n198) );
  OR2X8 U481 ( .A(n199), .B(n200), .Y(n197) );
  OR2XL U482 ( .A(SH[18]), .B(SH[16]), .Y(n216) );
  OR2X4 U483 ( .A(n209), .B(n210), .Y(n202) );
  NOR2BX1 U484 ( .AN(n4), .B(n329), .Y(B[0]) );
  OR2X2 U485 ( .A(n203), .B(n204), .Y(n199) );
  OR2XL U486 ( .A(SH[8]), .B(SH[9]), .Y(n213) );
  NOR2X1 U487 ( .A(n46), .B(n341), .Y(n14) );
  NOR2BX1 U488 ( .AN(n17), .B(n329), .Y(B[13]) );
  NOR2X1 U489 ( .A(n49), .B(n342), .Y(n17) );
  NOR2X1 U490 ( .A(n44), .B(n341), .Y(n12) );
  NOR2X1 U491 ( .A(n41), .B(n341), .Y(n9) );
  NOR2BX1 U492 ( .AN(n5), .B(n329), .Y(B[1]) );
  NOR2X1 U493 ( .A(n37), .B(n341), .Y(n5) );
  NOR2X1 U494 ( .A(n38), .B(n341), .Y(n6) );
  NOR2X1 U495 ( .A(n39), .B(n341), .Y(n7) );
  NOR2X1 U496 ( .A(n40), .B(n341), .Y(n8) );
  NOR2BX1 U497 ( .AN(n10), .B(n329), .Y(B[6]) );
  NOR2X1 U498 ( .A(n42), .B(n341), .Y(n10) );
  NOR2X1 U499 ( .A(n43), .B(n341), .Y(n11) );
  NOR2X1 U500 ( .A(n45), .B(n341), .Y(n13) );
  NOR2BX1 U501 ( .AN(n15), .B(n329), .Y(B[11]) );
  NOR2X1 U502 ( .A(n47), .B(n341), .Y(n15) );
  NOR2BX1 U503 ( .AN(n16), .B(n329), .Y(B[12]) );
  NOR2X1 U504 ( .A(n48), .B(n342), .Y(n16) );
  NOR2BX1 U505 ( .AN(n18), .B(n329), .Y(B[14]) );
  NOR2X1 U506 ( .A(n50), .B(n342), .Y(n18) );
  MXI2X1 U507 ( .A(n56), .B(n40), .S0(n342), .Y(n24) );
  MXI2X1 U508 ( .A(n120), .B(n116), .S0(n338), .Y(n88) );
  NAND2BX1 U509 ( .AN(n344), .B(n87), .Y(n55) );
  NAND2BX1 U510 ( .AN(n345), .B(n86), .Y(n54) );
  MXI2X1 U511 ( .A(n52), .B(n36), .S0(n342), .Y(n20) );
  NOR2X1 U512 ( .A(n51), .B(n342), .Y(n19) );
  MXI2X1 U513 ( .A(n125), .B(n121), .S0(n338), .Y(n93) );
  NAND2BX1 U514 ( .AN(n346), .B(n68), .Y(n36) );
  MXI2X1 U515 ( .A(n67), .B(n51), .S0(n340), .Y(n35) );
  CLKBUFX3 U516 ( .A(SH[1]), .Y(n333) );
  CLKBUFX3 U517 ( .A(SH[5]), .Y(n343) );
  CLKBUFX3 U518 ( .A(SH[5]), .Y(n346) );
  OR2X4 U519 ( .A(n213), .B(n214), .Y(n204) );
  OR2X2 U520 ( .A(n211), .B(n212), .Y(n203) );
  OR2XL U521 ( .A(SH[27]), .B(SH[23]), .Y(n210) );
  OR2XL U522 ( .A(SH[10]), .B(SH[11]), .Y(n214) );
  OR2XL U523 ( .A(SH[15]), .B(SH[31]), .Y(n209) );
  OR2X2 U524 ( .A(n205), .B(n206), .Y(n200) );
  OR2XL U525 ( .A(SH[17]), .B(SH[6]), .Y(n217) );
  OR2X2 U526 ( .A(n207), .B(n208), .Y(n201) );
  OR2XL U527 ( .A(SH[7]), .B(SH[25]), .Y(n208) );
  MXI2X1 U528 ( .A(A[22]), .B(A[14]), .S0(SH[3]), .Y(n186) );
endmodule


module ALU_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348;

  NOR2BX2 U256 ( .AN(n34), .B(n334), .Y(B[30]) );
  MXI2X2 U257 ( .A(n167), .B(n168), .S0(n337), .Y(n135) );
  INVX6 U258 ( .A(n324), .Y(n168) );
  MXI2X2 U259 ( .A(n135), .B(n137), .S0(n339), .Y(n103) );
  MXI2X4 U260 ( .A(n121), .B(n125), .S0(n342), .Y(n89) );
  NAND2BX2 U261 ( .AN(n348), .B(n76), .Y(n44) );
  NOR2X6 U262 ( .A(n195), .B(n336), .Y(n163) );
  MXI2X4 U263 ( .A(n125), .B(n129), .S0(n342), .Y(n93) );
  NOR2X4 U264 ( .A(n131), .B(n342), .Y(n99) );
  NOR2X1 U265 ( .A(n59), .B(n345), .Y(n27) );
  NAND2BX2 U266 ( .AN(n347), .B(n91), .Y(n59) );
  NOR2BX4 U267 ( .AN(n18), .B(n334), .Y(B[14]) );
  MXI2X2 U268 ( .A(n50), .B(n66), .S0(n346), .Y(n18) );
  MXI2X2 U269 ( .A(n37), .B(n53), .S0(n346), .Y(n5) );
  MXI2X2 U270 ( .A(n112), .B(n116), .S0(n343), .Y(n80) );
  MXI2X4 U271 ( .A(n148), .B(n150), .S0(n340), .Y(n116) );
  NAND2BX2 U272 ( .AN(n348), .B(n80), .Y(n48) );
  MXI2X4 U273 ( .A(A[25]), .B(A[17]), .S0(n331), .Y(n181) );
  MXI2X4 U274 ( .A(n139), .B(n141), .S0(n339), .Y(n107) );
  NOR2X1 U275 ( .A(n67), .B(n345), .Y(n35) );
  NAND2BX2 U276 ( .AN(n347), .B(n99), .Y(n67) );
  CLKMX2X4 U277 ( .A(n42), .B(n58), .S0(n346), .Y(n323) );
  MXI2X2 U278 ( .A(n102), .B(n106), .S0(n343), .Y(n70) );
  MXI2X2 U279 ( .A(n134), .B(n136), .S0(n339), .Y(n102) );
  NOR2X1 U280 ( .A(n57), .B(n345), .Y(n25) );
  NOR2X1 U281 ( .A(n58), .B(n345), .Y(n26) );
  NAND2BX2 U282 ( .AN(n347), .B(n90), .Y(n58) );
  NAND2BX2 U283 ( .AN(n347), .B(n88), .Y(n56) );
  MXI2X2 U284 ( .A(n169), .B(n170), .S0(n337), .Y(n137) );
  MXI2X2 U285 ( .A(n104), .B(n108), .S0(n343), .Y(n72) );
  NOR2BX2 U286 ( .AN(n33), .B(n334), .Y(B[29]) );
  INVX12 U287 ( .A(n331), .Y(n332) );
  CLKMX2X4 U288 ( .A(A[12]), .B(A[4]), .S0(n331), .Y(n324) );
  MX2X8 U289 ( .A(A[19]), .B(A[11]), .S0(n331), .Y(n325) );
  MX2X8 U290 ( .A(A[23]), .B(A[15]), .S0(n331), .Y(n328) );
  NOR2X2 U291 ( .A(n323), .B(n335), .Y(B[6]) );
  MXI2X2 U292 ( .A(n101), .B(n105), .S0(n343), .Y(n69) );
  MXI2X2 U293 ( .A(n133), .B(n135), .S0(n339), .Y(n101) );
  MXI2X2 U294 ( .A(n49), .B(n65), .S0(n346), .Y(n17) );
  NOR2BX4 U295 ( .AN(n17), .B(n335), .Y(B[13]) );
  BUFX8 U296 ( .A(n187), .Y(n330) );
  NOR2BX4 U297 ( .AN(n23), .B(n335), .Y(B[19]) );
  MXI2X2 U298 ( .A(n40), .B(n56), .S0(n346), .Y(n8) );
  NAND2BX2 U299 ( .AN(SH[5]), .B(n72), .Y(n40) );
  MXI2X4 U300 ( .A(n177), .B(n178), .S0(n337), .Y(n145) );
  MXI2X2 U301 ( .A(n111), .B(n115), .S0(n343), .Y(n79) );
  NOR2BX4 U302 ( .AN(n9), .B(n335), .Y(B[5]) );
  MXI2X2 U303 ( .A(n41), .B(n57), .S0(n346), .Y(n9) );
  MXI2X4 U304 ( .A(n142), .B(n144), .S0(n339), .Y(n110) );
  MXI2X4 U305 ( .A(n144), .B(n326), .S0(n340), .Y(n112) );
  MXI2X4 U306 ( .A(n176), .B(n177), .S0(n337), .Y(n144) );
  MXI2X2 U307 ( .A(n110), .B(n114), .S0(n343), .Y(n78) );
  MXI2X4 U308 ( .A(n190), .B(n191), .S0(n336), .Y(n158) );
  NOR2BX2 U309 ( .AN(n28), .B(n334), .Y(B[24]) );
  NOR2X1 U310 ( .A(n60), .B(n345), .Y(n28) );
  MXI2X2 U311 ( .A(n44), .B(n60), .S0(n346), .Y(n12) );
  MXI2X4 U312 ( .A(n182), .B(n183), .S0(n336), .Y(n150) );
  INVX8 U313 ( .A(n329), .Y(n183) );
  MXI2X2 U314 ( .A(n114), .B(n118), .S0(n343), .Y(n82) );
  MXI2X4 U315 ( .A(n150), .B(n152), .S0(n340), .Y(n118) );
  MXI2X4 U316 ( .A(n326), .B(n148), .S0(n340), .Y(n114) );
  MXI2X2 U317 ( .A(n115), .B(n119), .S0(n343), .Y(n83) );
  NOR2BX4 U318 ( .AN(n19), .B(n334), .Y(B[15]) );
  MXI2X2 U319 ( .A(n51), .B(n67), .S0(n346), .Y(n19) );
  MXI2X4 U320 ( .A(n141), .B(n143), .S0(n339), .Y(n109) );
  MXI2X4 U321 ( .A(n143), .B(n145), .S0(n339), .Y(n111) );
  MXI2X4 U322 ( .A(n175), .B(n176), .S0(n337), .Y(n143) );
  MXI2X2 U323 ( .A(n105), .B(n109), .S0(n343), .Y(n73) );
  NOR2BX4 U324 ( .AN(n20), .B(n335), .Y(B[16]) );
  NOR2X2 U325 ( .A(n52), .B(n346), .Y(n20) );
  NOR2BX4 U326 ( .AN(n22), .B(n334), .Y(B[18]) );
  NOR2X2 U327 ( .A(n54), .B(n346), .Y(n22) );
  MXI2X4 U328 ( .A(A[22]), .B(A[30]), .S0(n333), .Y(n186) );
  MXI2X4 U329 ( .A(n152), .B(n154), .S0(n340), .Y(n120) );
  MXI2X4 U330 ( .A(n186), .B(n187), .S0(n336), .Y(n154) );
  MXI2X2 U331 ( .A(n166), .B(n167), .S0(n337), .Y(n134) );
  NAND2BX2 U332 ( .AN(SH[5]), .B(n68), .Y(n36) );
  NAND2BX2 U333 ( .AN(n333), .B(A[31]), .Y(n195) );
  MXI2X4 U334 ( .A(n178), .B(n179), .S0(n337), .Y(n326) );
  MXI2X4 U335 ( .A(n192), .B(n193), .S0(n336), .Y(n160) );
  INVX20 U336 ( .A(n331), .Y(n333) );
  MXI2X4 U337 ( .A(n194), .B(n195), .S0(n336), .Y(n162) );
  MXI2X4 U338 ( .A(n117), .B(n121), .S0(n342), .Y(n85) );
  NOR2X2 U339 ( .A(n53), .B(n346), .Y(n21) );
  MXI2X4 U340 ( .A(n181), .B(n182), .S0(n336), .Y(n149) );
  MXI2X4 U341 ( .A(n185), .B(n186), .S0(n336), .Y(n153) );
  MXI2X2 U342 ( .A(A[8]), .B(A[16]), .S0(n332), .Y(n172) );
  NAND2BX1 U343 ( .AN(n348), .B(n79), .Y(n47) );
  BUFX2 U344 ( .A(SH[5]), .Y(n348) );
  INVX20 U345 ( .A(SH[3]), .Y(n331) );
  MXI2X2 U346 ( .A(n100), .B(n104), .S0(n342), .Y(n68) );
  NOR2BX4 U347 ( .AN(n8), .B(n335), .Y(B[4]) );
  MXI2X4 U348 ( .A(n137), .B(n139), .S0(n339), .Y(n105) );
  NOR2BX4 U349 ( .AN(n5), .B(n335), .Y(B[1]) );
  MXI2X4 U350 ( .A(n140), .B(n142), .S0(n339), .Y(n108) );
  NOR2BX4 U351 ( .AN(n12), .B(n335), .Y(B[8]) );
  MXI2X1 U352 ( .A(A[5]), .B(A[13]), .S0(SH[3]), .Y(n169) );
  NOR2X1 U353 ( .A(n55), .B(n346), .Y(n23) );
  NAND2BX2 U354 ( .AN(n347), .B(n87), .Y(n55) );
  MXI2X1 U355 ( .A(n165), .B(n166), .S0(n337), .Y(n133) );
  MXI2X2 U356 ( .A(n116), .B(n120), .S0(SH[2]), .Y(n84) );
  NAND2BX2 U357 ( .AN(SH[3]), .B(A[29]), .Y(n193) );
  MXI2X4 U358 ( .A(n151), .B(n153), .S0(n340), .Y(n119) );
  MXI2X4 U359 ( .A(n174), .B(n175), .S0(n337), .Y(n142) );
  MXI2X4 U360 ( .A(n173), .B(n174), .S0(n337), .Y(n141) );
  MXI2X2 U361 ( .A(A[10]), .B(A[18]), .S0(SH[3]), .Y(n174) );
  CLKINVX20 U362 ( .A(n325), .Y(n175) );
  NOR2BX2 U363 ( .AN(n26), .B(n334), .Y(B[22]) );
  MXI2X4 U364 ( .A(A[13]), .B(A[21]), .S0(n332), .Y(n177) );
  MXI2X2 U365 ( .A(A[14]), .B(A[22]), .S0(SH[3]), .Y(n178) );
  MXI2X4 U366 ( .A(n180), .B(n181), .S0(n337), .Y(n148) );
  MXI2X4 U367 ( .A(n179), .B(n180), .S0(n337), .Y(n147) );
  MXI2X2 U368 ( .A(A[16]), .B(A[24]), .S0(n333), .Y(n180) );
  MXI2X4 U369 ( .A(n330), .B(n188), .S0(n336), .Y(n155) );
  MXI2X4 U370 ( .A(A[3]), .B(A[11]), .S0(n333), .Y(n167) );
  BUFX8 U371 ( .A(n184), .Y(n327) );
  CLKINVX20 U372 ( .A(n328), .Y(n179) );
  CLKMX2X8 U373 ( .A(A[27]), .B(A[19]), .S0(n331), .Y(n329) );
  MXI2X1 U374 ( .A(A[2]), .B(A[10]), .S0(n333), .Y(n166) );
  NAND2BX2 U375 ( .AN(SH[3]), .B(A[30]), .Y(n194) );
  MXI2X2 U376 ( .A(A[23]), .B(A[31]), .S0(n333), .Y(n187) );
  NOR2BX4 U377 ( .AN(n11), .B(n334), .Y(B[7]) );
  NOR2BX2 U378 ( .AN(n35), .B(n334), .Y(B[31]) );
  NOR2BX4 U379 ( .AN(n29), .B(n334), .Y(B[25]) );
  NOR2BX2 U380 ( .AN(n32), .B(n334), .Y(B[28]) );
  NOR2BX2 U381 ( .AN(n25), .B(n334), .Y(B[21]) );
  NOR2BX4 U382 ( .AN(n24), .B(n334), .Y(B[20]) );
  BUFX20 U383 ( .A(n3), .Y(n334) );
  NAND2BX4 U384 ( .AN(n333), .B(A[27]), .Y(n191) );
  NOR2X1 U385 ( .A(n66), .B(n345), .Y(n34) );
  NAND2BX2 U386 ( .AN(n347), .B(n98), .Y(n66) );
  MXI2X4 U387 ( .A(n147), .B(n149), .S0(n340), .Y(n115) );
  MXI2X4 U388 ( .A(n145), .B(n147), .S0(n340), .Y(n113) );
  NOR2X1 U389 ( .A(n65), .B(n345), .Y(n33) );
  NAND2BX2 U390 ( .AN(n347), .B(n97), .Y(n65) );
  MXI2X4 U391 ( .A(A[6]), .B(A[14]), .S0(n332), .Y(n170) );
  NAND2BX4 U392 ( .AN(SH[3]), .B(A[26]), .Y(n190) );
  MXI2X4 U393 ( .A(n327), .B(n185), .S0(n336), .Y(n152) );
  MXI2X1 U394 ( .A(A[20]), .B(A[28]), .S0(SH[3]), .Y(n184) );
  MXI2X4 U395 ( .A(n168), .B(n169), .S0(n337), .Y(n136) );
  MXI2X4 U396 ( .A(A[12]), .B(A[20]), .S0(n332), .Y(n176) );
  NOR2BX4 U397 ( .AN(n7), .B(n335), .Y(B[3]) );
  NAND2BX2 U398 ( .AN(SH[5]), .B(n71), .Y(n39) );
  OR2X4 U399 ( .A(n211), .B(n212), .Y(n203) );
  OR2X2 U400 ( .A(SH[21]), .B(SH[19]), .Y(n211) );
  MXI2X2 U401 ( .A(n123), .B(n127), .S0(n342), .Y(n91) );
  NAND2BX4 U402 ( .AN(SH[3]), .B(A[25]), .Y(n189) );
  NAND2BX2 U403 ( .AN(n348), .B(n74), .Y(n42) );
  MXI2X2 U404 ( .A(n138), .B(n140), .S0(n339), .Y(n106) );
  MXI2X4 U405 ( .A(n172), .B(n173), .S0(n337), .Y(n140) );
  NAND2BX2 U406 ( .AN(n347), .B(n89), .Y(n57) );
  MXI2X4 U407 ( .A(n157), .B(n159), .S0(n341), .Y(n125) );
  MXI2X4 U408 ( .A(n189), .B(n190), .S0(n336), .Y(n157) );
  OR2X4 U409 ( .A(SH[22]), .B(SH[20]), .Y(n220) );
  NOR2BX1 U410 ( .AN(n27), .B(n334), .Y(B[23]) );
  MXI2X4 U411 ( .A(n193), .B(n194), .S0(n336), .Y(n161) );
  MXI2X4 U412 ( .A(n154), .B(n156), .S0(n340), .Y(n122) );
  MXI2X4 U413 ( .A(n188), .B(n189), .S0(n336), .Y(n156) );
  MXI2X2 U414 ( .A(n118), .B(n122), .S0(n342), .Y(n86) );
  MXI2X4 U415 ( .A(n158), .B(n160), .S0(n341), .Y(n126) );
  NOR2BX4 U416 ( .AN(n13), .B(n335), .Y(B[9]) );
  BUFX20 U417 ( .A(n3), .Y(n335) );
  MXI2X2 U418 ( .A(n45), .B(n61), .S0(n346), .Y(n13) );
  NOR2X1 U419 ( .A(n61), .B(n345), .Y(n29) );
  NAND2BX2 U420 ( .AN(n347), .B(n93), .Y(n61) );
  MXI2X4 U421 ( .A(n156), .B(n158), .S0(n341), .Y(n124) );
  MXI2X4 U422 ( .A(n120), .B(n124), .S0(n342), .Y(n88) );
  NOR2X1 U423 ( .A(n56), .B(n345), .Y(n24) );
  NOR2BX4 U424 ( .AN(n6), .B(n335), .Y(B[2]) );
  MXI2XL U425 ( .A(n106), .B(n110), .S0(n343), .Y(n74) );
  NAND2BX2 U426 ( .AN(SH[5]), .B(n69), .Y(n37) );
  MXI2X4 U427 ( .A(n171), .B(n172), .S0(n337), .Y(n139) );
  MXI2X4 U428 ( .A(A[7]), .B(A[15]), .S0(n333), .Y(n171) );
  NAND2BX2 U429 ( .AN(n348), .B(n77), .Y(n45) );
  MXI2X4 U430 ( .A(n155), .B(n157), .S0(n340), .Y(n123) );
  NAND2BX1 U431 ( .AN(SH[3]), .B(A[24]), .Y(n188) );
  NAND2BX2 U432 ( .AN(n347), .B(n96), .Y(n64) );
  NOR2X4 U433 ( .A(n128), .B(n342), .Y(n96) );
  NAND2BX4 U434 ( .AN(SH[3]), .B(A[28]), .Y(n192) );
  MXI2X4 U435 ( .A(n160), .B(n162), .S0(n341), .Y(n128) );
  MXI2X4 U436 ( .A(n183), .B(n327), .S0(n336), .Y(n151) );
  NAND2BX2 U437 ( .AN(n348), .B(n86), .Y(n54) );
  NAND2BX2 U438 ( .AN(SH[5]), .B(n70), .Y(n38) );
  MXI2X2 U439 ( .A(n170), .B(n171), .S0(n337), .Y(n138) );
  MXI2X4 U440 ( .A(n149), .B(n151), .S0(n340), .Y(n117) );
  MXI2X2 U441 ( .A(A[21]), .B(A[29]), .S0(SH[3]), .Y(n185) );
  MXI2X4 U442 ( .A(n127), .B(n131), .S0(n342), .Y(n95) );
  MXI2X4 U443 ( .A(n159), .B(n161), .S0(n341), .Y(n127) );
  NOR2X1 U444 ( .A(n63), .B(n345), .Y(n31) );
  NAND2BX2 U445 ( .AN(n347), .B(n95), .Y(n63) );
  NAND2BX2 U446 ( .AN(n341), .B(n163), .Y(n131) );
  BUFX12 U447 ( .A(n338), .Y(n341) );
  MXI2X2 U448 ( .A(n191), .B(n192), .S0(n336), .Y(n159) );
  MXI2X2 U449 ( .A(n113), .B(n117), .S0(n343), .Y(n81) );
  NAND2BX2 U450 ( .AN(n348), .B(n84), .Y(n52) );
  MXI2X4 U451 ( .A(n153), .B(n155), .S0(n340), .Y(n121) );
  NAND2BX2 U452 ( .AN(n347), .B(n92), .Y(n60) );
  MXI2X2 U453 ( .A(n124), .B(n128), .S0(n342), .Y(n92) );
  BUFX20 U454 ( .A(SH[2]), .Y(n342) );
  MXI2X2 U455 ( .A(n136), .B(n138), .S0(n339), .Y(n104) );
  NAND2BX2 U456 ( .AN(n348), .B(n85), .Y(n53) );
  MXI2X2 U457 ( .A(A[18]), .B(A[26]), .S0(SH[3]), .Y(n182) );
  CLKBUFX2 U458 ( .A(SH[4]), .Y(n344) );
  NOR2X1 U459 ( .A(n62), .B(n345), .Y(n30) );
  NAND2BX2 U460 ( .AN(n347), .B(n94), .Y(n62) );
  NAND2BX2 U461 ( .AN(n341), .B(n162), .Y(n130) );
  MXI2X2 U462 ( .A(n126), .B(n130), .S0(n342), .Y(n94) );
  MXI2X2 U463 ( .A(n122), .B(n126), .S0(n342), .Y(n90) );
  MXI2X2 U464 ( .A(n161), .B(n163), .S0(n341), .Y(n129) );
  BUFX20 U465 ( .A(SH[0]), .Y(n336) );
  BUFX16 U466 ( .A(SH[1]), .Y(n340) );
  BUFX20 U467 ( .A(SH[0]), .Y(n337) );
  BUFX8 U468 ( .A(SH[1]), .Y(n339) );
  BUFX12 U469 ( .A(SH[2]), .Y(n343) );
  BUFX12 U470 ( .A(n344), .Y(n346) );
  CLKBUFX2 U471 ( .A(SH[4]), .Y(n345) );
  NOR2BX1 U472 ( .AN(n30), .B(n334), .Y(B[26]) );
  NOR2BX1 U473 ( .AN(n31), .B(n334), .Y(B[27]) );
  OR2X8 U474 ( .A(n197), .B(n198), .Y(n3) );
  OR2X8 U475 ( .A(n201), .B(n202), .Y(n198) );
  OR2X8 U476 ( .A(n199), .B(n200), .Y(n197) );
  OR2XL U477 ( .A(SH[18]), .B(SH[16]), .Y(n216) );
  NOR2XL U478 ( .A(n64), .B(n345), .Y(n32) );
  MXI2X1 U479 ( .A(n103), .B(n107), .S0(n343), .Y(n71) );
  NOR2BX1 U480 ( .AN(n4), .B(n335), .Y(B[0]) );
  OR2X4 U481 ( .A(n209), .B(n210), .Y(n202) );
  OR2X2 U482 ( .A(n203), .B(n204), .Y(n199) );
  OR2XL U483 ( .A(SH[8]), .B(SH[9]), .Y(n213) );
  MXI2X1 U484 ( .A(n119), .B(n123), .S0(n342), .Y(n87) );
  NOR2X1 U485 ( .A(n130), .B(n342), .Y(n98) );
  NOR2X1 U486 ( .A(n129), .B(n342), .Y(n97) );
  MXI2X1 U487 ( .A(n107), .B(n111), .S0(n343), .Y(n75) );
  MXI2X1 U488 ( .A(n109), .B(n113), .S0(n343), .Y(n77) );
  MXI2X1 U489 ( .A(n108), .B(n112), .S0(n343), .Y(n76) );
  CLKBUFX3 U490 ( .A(SH[5]), .Y(n347) );
  NOR2BX1 U491 ( .AN(n14), .B(n335), .Y(B[10]) );
  MXI2X1 U492 ( .A(n46), .B(n62), .S0(n346), .Y(n14) );
  NAND2BX1 U493 ( .AN(n348), .B(n78), .Y(n46) );
  MXI2X1 U494 ( .A(n36), .B(n52), .S0(n346), .Y(n4) );
  NAND2BX1 U495 ( .AN(n348), .B(n83), .Y(n51) );
  NAND2BX1 U496 ( .AN(n348), .B(n81), .Y(n49) );
  NOR2BX1 U497 ( .AN(n16), .B(n335), .Y(B[12]) );
  MXI2X1 U498 ( .A(n48), .B(n64), .S0(n346), .Y(n16) );
  NOR2BX1 U499 ( .AN(n15), .B(n335), .Y(B[11]) );
  MXI2X1 U500 ( .A(n47), .B(n63), .S0(n346), .Y(n15) );
  NAND2BX1 U501 ( .AN(n348), .B(n82), .Y(n50) );
  MXI2X1 U502 ( .A(n39), .B(n55), .S0(n346), .Y(n7) );
  MXI2X1 U503 ( .A(n38), .B(n54), .S0(n346), .Y(n6) );
  MXI2X1 U504 ( .A(n43), .B(n59), .S0(n346), .Y(n11) );
  NAND2BX1 U505 ( .AN(n348), .B(n75), .Y(n43) );
  NAND2BX1 U506 ( .AN(n348), .B(n73), .Y(n41) );
  NOR2BX1 U507 ( .AN(n21), .B(n334), .Y(B[17]) );
  CLKBUFX3 U508 ( .A(SH[1]), .Y(n338) );
  OR2XL U509 ( .A(SH[12]), .B(SH[28]), .Y(n212) );
  OR2X4 U510 ( .A(n213), .B(n214), .Y(n204) );
  MXI2X1 U511 ( .A(n132), .B(n134), .S0(n339), .Y(n100) );
  MXI2X1 U512 ( .A(n164), .B(n165), .S0(n337), .Y(n132) );
  OR2XL U513 ( .A(SH[24]), .B(SH[14]), .Y(n218) );
  OR2XL U514 ( .A(SH[30]), .B(SH[26]), .Y(n219) );
  OR2XL U515 ( .A(SH[13]), .B(SH[29]), .Y(n215) );
  OR2XL U516 ( .A(SH[27]), .B(SH[23]), .Y(n210) );
  OR2XL U517 ( .A(SH[10]), .B(SH[11]), .Y(n214) );
  OR2XL U518 ( .A(SH[15]), .B(SH[31]), .Y(n209) );
  OR2X4 U519 ( .A(n205), .B(n206), .Y(n200) );
  OR2X4 U520 ( .A(n217), .B(n218), .Y(n206) );
  OR2X4 U521 ( .A(n215), .B(n216), .Y(n205) );
  OR2XL U522 ( .A(SH[17]), .B(SH[6]), .Y(n217) );
  OR2X4 U523 ( .A(n207), .B(n208), .Y(n201) );
  OR2XL U524 ( .A(SH[7]), .B(SH[25]), .Y(n208) );
  OR2X1 U525 ( .A(n219), .B(n220), .Y(n207) );
  MXI2XL U526 ( .A(A[0]), .B(A[8]), .S0(n333), .Y(n164) );
  MXI2X1 U527 ( .A(A[1]), .B(A[9]), .S0(n333), .Y(n165) );
  MXI2X1 U528 ( .A(A[9]), .B(A[17]), .S0(SH[3]), .Y(n173) );
endmodule


module ALU ( ALUOp_regD, funct_regD, ALUinA, ALUinB, ALUout );
  input [5:0] ALUOp_regD;
  input [5:0] funct_regD;
  input [31:0] ALUinA;
  input [31:0] ALUinB;
  output [31:0] ALUout;
  wire   N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N441, n429, n444, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542;

  ALU_DW01_add_1 r319 ( .A(ALUinA), .B({ALUinB[31:6], n123, n121, n119, n117, 
        n115, n113}), .CI(1'b0), .SUM({N280, N279, N278, N277, N276, N275, 
        N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, 
        N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, 
        N250, N249}) );
  ALU_DW01_sub_1 sub_1145 ( .A(ALUinA), .B({ALUinB[31:6], n123, n121, n119, 
        n117, n115, n113}), .CI(1'b0), .DIFF({N312, N311, N310, N309, N308, 
        N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281}) );
  ALU_DW_cmp_1 r323 ( .A(ALUinA), .B({ALUinB[31:6], n123, n121, n6, n117, n115, 
        n113}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N441)
         );
  ALU_DW_leftsh_1 sll_1160 ( .A(ALUinA), .SH({ALUinB[31:6], n123, n121, n7, 
        n117, n115, n113}), .B({N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345}) );
  ALU_DW_rightsh_1 r322 ( .A(ALUinA), .DATA_TC(1'b0), .SH({ALUinB[31:6], n123, 
        n121, n6, n117, n115, n113}), .B({N408, N407, N406, N405, N404, N403, 
        N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, 
        N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, 
        N378, N377}) );
  NOR4X4 U8 ( .A(n308), .B(n307), .C(n306), .D(n305), .Y(n311) );
  OAI2BB2X2 U9 ( .B0(n1), .B1(n129), .A0N(N269), .A1N(n84), .Y(n396) );
  INVX1 U10 ( .A(N397), .Y(n1) );
  AO22X1 U11 ( .A0(N384), .A1(n88), .B0(N256), .B1(n85), .Y(n249) );
  NOR4X4 U12 ( .A(n489), .B(n488), .C(n487), .D(n486), .Y(n493) );
  AO22X2 U13 ( .A0(N290), .A1(n82), .B0(N354), .B1(n80), .Y(n274) );
  BUFX3 U14 ( .A(n523), .Y(n86) );
  NAND3BX2 U15 ( .AN(funct_regD[5]), .B(n141), .C(n142), .Y(n129) );
  NOR4X4 U16 ( .A(n214), .B(n213), .C(n215), .D(n212), .Y(n218) );
  AO22X2 U17 ( .A0(N285), .A1(n82), .B0(N349), .B1(n80), .Y(n214) );
  NAND2X2 U18 ( .A(n211), .B(n122), .Y(n216) );
  CLKINVX8 U19 ( .A(ALUinB[4]), .Y(n122) );
  NOR4BX2 U20 ( .AN(n2), .B(n341), .C(n342), .D(n340), .Y(n346) );
  CLKINVX20 U21 ( .A(n343), .Y(n2) );
  INVX1 U22 ( .A(N271), .Y(n424) );
  CLKINVX8 U23 ( .A(n120), .Y(n119) );
  NAND2X1 U24 ( .A(n201), .B(n120), .Y(n206) );
  NOR4BX2 U25 ( .AN(n3), .B(n262), .C(n261), .D(n260), .Y(n267) );
  CLKINVX20 U26 ( .A(n263), .Y(n3) );
  AO22X2 U27 ( .A0(N396), .A1(n87), .B0(N268), .B1(n84), .Y(n385) );
  AO22X1 U28 ( .A0(N381), .A1(n88), .B0(N253), .B1(n85), .Y(n213) );
  NOR4BX2 U29 ( .AN(n4), .B(n386), .C(n385), .D(n384), .Y(n390) );
  CLKINVX20 U30 ( .A(n387), .Y(n4) );
  NOR4X4 U31 ( .A(n224), .B(n225), .C(n226), .D(n223), .Y(n230) );
  AO22X2 U32 ( .A0(N286), .A1(n82), .B0(N350), .B1(n80), .Y(n225) );
  NOR4X2 U33 ( .A(n297), .B(n296), .C(n295), .D(n294), .Y(n300) );
  NOR4BX2 U34 ( .AN(n5), .B(n396), .C(n397), .D(n395), .Y(n401) );
  CLKINVX20 U35 ( .A(n398), .Y(n5) );
  NOR4X2 U36 ( .A(n239), .B(n238), .C(n237), .D(n236), .Y(n243) );
  NOR4X4 U37 ( .A(n332), .B(n331), .C(n330), .D(n329), .Y(n335) );
  AO22X2 U38 ( .A0(N391), .A1(n87), .B0(N263), .B1(n85), .Y(n330) );
  AO22X2 U39 ( .A0(N295), .A1(n82), .B0(N359), .B1(n80), .Y(n331) );
  NOR4X2 U40 ( .A(n319), .B(n320), .C(n318), .D(n317), .Y(n324) );
  INVX16 U41 ( .A(n122), .Y(n121) );
  AO22X1 U42 ( .A0(N294), .A1(n82), .B0(N358), .B1(n80), .Y(n319) );
  NOR4X2 U43 ( .A(n454), .B(n453), .C(n455), .D(n452), .Y(n458) );
  NOR4X4 U44 ( .A(n510), .B(n511), .C(n512), .D(n509), .Y(n515) );
  AO22X2 U45 ( .A0(N311), .A1(n83), .B0(N375), .B1(n81), .Y(n511) );
  AO22X1 U46 ( .A0(N392), .A1(n87), .B0(N264), .B1(n85), .Y(n341) );
  AO22X2 U47 ( .A0(N296), .A1(n82), .B0(N360), .B1(n80), .Y(n342) );
  AO22X2 U48 ( .A0(N297), .A1(n83), .B0(N361), .B1(n80), .Y(n353) );
  INVX20 U49 ( .A(n120), .Y(n6) );
  INVX20 U50 ( .A(n120), .Y(n7) );
  CLKINVX12 U51 ( .A(ALUinB[3]), .Y(n120) );
  OAI221X1 U52 ( .A0(n110), .A1(n448), .B0(n447), .B1(n103), .C0(n446), .Y(
        ALUout[24]) );
  NOR4X4 U53 ( .A(n443), .B(n442), .C(n441), .D(n440), .Y(n447) );
  OAI221X4 U54 ( .A0(n111), .A1(n325), .B0(n324), .B1(n103), .C0(n323), .Y(
        ALUout[13]) );
  OAI221X1 U55 ( .A0(n111), .A1(n347), .B0(n346), .B1(n103), .C0(n345), .Y(
        ALUout[15]) );
  NOR4X2 U56 ( .A(n354), .B(n353), .C(n352), .D(n351), .Y(n357) );
  XNOR2XL U57 ( .A(n176), .B(n115), .Y(n8) );
  AND2XL U58 ( .A(n115), .B(ALUinA[1]), .Y(n9) );
  AND2XL U59 ( .A(n6), .B(ALUinA[3]), .Y(n10) );
  XNOR2XL U60 ( .A(n201), .B(n7), .Y(n11) );
  AND2XL U61 ( .A(n123), .B(ALUinA[5]), .Y(n12) );
  INVX20 U62 ( .A(n124), .Y(n123) );
  XNOR2XL U63 ( .A(n247), .B(ALUinB[7]), .Y(n13) );
  AND2XL U64 ( .A(ALUinB[7]), .B(ALUinA[7]), .Y(n14) );
  AND2XL U65 ( .A(ALUinB[8]), .B(ALUinA[8]), .Y(n15) );
  AND2XL U66 ( .A(ALUinB[9]), .B(ALUinA[9]), .Y(n16) );
  XNOR2XL U67 ( .A(n271), .B(ALUinB[9]), .Y(n17) );
  XNOR2XL U68 ( .A(n293), .B(ALUinB[11]), .Y(n18) );
  AND2XL U69 ( .A(ALUinB[11]), .B(ALUinA[11]), .Y(n24) );
  AND2XL U70 ( .A(ALUinB[12]), .B(ALUinA[12]), .Y(n25) );
  XNOR2XL U71 ( .A(n304), .B(ALUinB[12]), .Y(n26) );
  AND2XL U72 ( .A(n117), .B(ALUinA[2]), .Y(n27) );
  CLKINVX12 U73 ( .A(n118), .Y(n117) );
  XNOR2XL U74 ( .A(n282), .B(ALUinB[10]), .Y(n28) );
  AND2XL U75 ( .A(ALUinB[10]), .B(ALUinA[10]), .Y(n29) );
  AND2XL U76 ( .A(n121), .B(ALUinA[4]), .Y(n30) );
  XNOR2XL U77 ( .A(n211), .B(n121), .Y(n31) );
  AND2XL U78 ( .A(ALUinB[6]), .B(ALUinA[6]), .Y(n32) );
  AND2XL U79 ( .A(ALUinB[13]), .B(ALUinA[13]), .Y(n33) );
  XNOR2XL U80 ( .A(n328), .B(ALUinB[14]), .Y(n34) );
  AND2XL U81 ( .A(ALUinB[14]), .B(ALUinA[14]), .Y(n35) );
  AND2XL U82 ( .A(ALUinB[15]), .B(ALUinA[15]), .Y(n36) );
  XNOR2XL U83 ( .A(n339), .B(ALUinB[15]), .Y(n37) );
  XNOR2XL U84 ( .A(n350), .B(ALUinB[16]), .Y(n38) );
  AND2XL U85 ( .A(ALUinB[16]), .B(ALUinA[16]), .Y(n39) );
  AND2XL U86 ( .A(ALUinB[17]), .B(ALUinA[17]), .Y(n40) );
  XNOR2XL U87 ( .A(n361), .B(ALUinB[17]), .Y(n41) );
  XNOR2XL U88 ( .A(n372), .B(ALUinB[18]), .Y(n42) );
  AND2XL U89 ( .A(ALUinB[18]), .B(ALUinA[18]), .Y(n43) );
  AND2XL U90 ( .A(ALUinB[19]), .B(ALUinA[19]), .Y(n44) );
  XNOR2XL U91 ( .A(n383), .B(ALUinB[19]), .Y(n45) );
  AND2XL U92 ( .A(ALUinB[20]), .B(ALUinA[20]), .Y(n46) );
  XNOR2XL U93 ( .A(n394), .B(ALUinB[20]), .Y(n47) );
  XNOR2XL U94 ( .A(n416), .B(ALUinB[22]), .Y(n48) );
  AND2XL U95 ( .A(ALUinB[22]), .B(ALUinA[22]), .Y(n49) );
  XNOR2XL U96 ( .A(n427), .B(ALUinB[23]), .Y(n50) );
  AND2XL U97 ( .A(ALUinB[23]), .B(ALUinA[23]), .Y(n51) );
  AND2XL U98 ( .A(ALUinB[24]), .B(ALUinA[24]), .Y(n52) );
  XNOR2XL U99 ( .A(n439), .B(ALUinB[24]), .Y(n53) );
  XNOR2XL U100 ( .A(n451), .B(ALUinB[25]), .Y(n54) );
  AND2XL U101 ( .A(ALUinB[25]), .B(ALUinA[25]), .Y(n55) );
  XNOR2XL U102 ( .A(n405), .B(ALUinB[21]), .Y(n56) );
  AND2XL U103 ( .A(ALUinB[21]), .B(ALUinA[21]), .Y(n57) );
  AND2XL U104 ( .A(ALUinB[26]), .B(ALUinA[26]), .Y(n58) );
  XNOR2XL U105 ( .A(n462), .B(ALUinB[26]), .Y(n59) );
  AND2XL U106 ( .A(ALUinB[27]), .B(ALUinA[27]), .Y(n60) );
  XNOR2XL U107 ( .A(n473), .B(ALUinB[27]), .Y(n61) );
  AND2XL U108 ( .A(ALUinB[30]), .B(ALUinA[30]), .Y(n62) );
  XNOR2XL U109 ( .A(n508), .B(ALUinB[30]), .Y(n63) );
  AND2XL U110 ( .A(ALUinB[28]), .B(ALUinA[28]), .Y(n64) );
  XNOR2XL U111 ( .A(n524), .B(ALUinB[31]), .Y(n65) );
  AND2XL U112 ( .A(ALUinB[31]), .B(ALUinA[31]), .Y(n66) );
  AND2XL U113 ( .A(ALUinB[29]), .B(ALUinA[29]), .Y(n67) );
  XNOR2XL U114 ( .A(n497), .B(ALUinB[29]), .Y(n68) );
  AO22X2 U115 ( .A0(N406), .A1(n86), .B0(N278), .B1(n84), .Y(n499) );
  AOI21X1 U116 ( .A0(n444), .A1(n132), .B0(funct_regD[1]), .Y(n522) );
  INVX1 U117 ( .A(n175), .Y(n526) );
  INVX1 U118 ( .A(n173), .Y(n519) );
  AO22X1 U119 ( .A0(n93), .A1(n65), .B0(n89), .B1(n66), .Y(n527) );
  INVX1 U120 ( .A(n485), .Y(n491) );
  CLKINVX4 U121 ( .A(ALUinB[1]), .Y(n116) );
  AO22XL U122 ( .A0(n93), .A1(n491), .B0(n64), .B1(n89), .Y(n486) );
  NOR4X4 U123 ( .A(n407), .B(n408), .C(n409), .D(n406), .Y(n412) );
  CLKINVX12 U124 ( .A(n116), .Y(n115) );
  CLKAND2X12 U125 ( .A(n540), .B(n157), .Y(n69) );
  INVX3 U126 ( .A(n182), .Y(n533) );
  BUFX2 U127 ( .A(n533), .Y(n97) );
  BUFX2 U128 ( .A(n533), .Y(n98) );
  CLKAND2X8 U129 ( .A(funct_regD[2]), .B(funct_regD[5]), .Y(n70) );
  AND2X1 U130 ( .A(n143), .B(n114), .Y(n71) );
  CLKAND2X3 U131 ( .A(ALUOp_regD[2]), .B(ALUOp_regD[3]), .Y(n72) );
  CLKAND2X3 U132 ( .A(n141), .B(n140), .Y(n73) );
  OAI221X2 U133 ( .A0(n112), .A1(n199), .B0(n198), .B1(n102), .C0(n197), .Y(
        ALUout[2]) );
  AO22X4 U134 ( .A0(N380), .A1(n88), .B0(N252), .B1(n85), .Y(n203) );
  OAI221X2 U135 ( .A0(n112), .A1(n209), .B0(n208), .B1(n102), .C0(n207), .Y(
        ALUout[3]) );
  OAI221X2 U136 ( .A0(n112), .A1(n187), .B0(n186), .B1(n102), .C0(n185), .Y(
        ALUout[1]) );
  OAI221X2 U137 ( .A0(n110), .A1(n494), .B0(n493), .B1(n104), .C0(n492), .Y(
        ALUout[28]) );
  AO22X2 U138 ( .A0(N386), .A1(n87), .B0(N258), .B1(n85), .Y(n273) );
  AO22X2 U139 ( .A0(N291), .A1(n82), .B0(N355), .B1(n80), .Y(n285) );
  AO22X4 U140 ( .A0(N387), .A1(n87), .B0(N259), .B1(n85), .Y(n284) );
  OAI221X1 U141 ( .A0(n111), .A1(n312), .B0(n311), .B1(n102), .C0(n310), .Y(
        ALUout[12]) );
  AO22X2 U142 ( .A0(N304), .A1(n83), .B0(N368), .B1(n81), .Y(n431) );
  AO22X2 U143 ( .A0(N400), .A1(n86), .B0(N272), .B1(n84), .Y(n430) );
  AO22X2 U144 ( .A0(N302), .A1(n83), .B0(N366), .B1(n81), .Y(n408) );
  AO22X2 U145 ( .A0(N388), .A1(n87), .B0(N260), .B1(n85), .Y(n295) );
  AO22X4 U146 ( .A0(N283), .A1(n82), .B0(N347), .B1(n80), .Y(n193) );
  AO22X4 U147 ( .A0(N379), .A1(n88), .B0(N251), .B1(n85), .Y(n192) );
  NAND4X1 U148 ( .A(n69), .B(n125), .C(n150), .D(n164), .Y(n152) );
  AO22X4 U149 ( .A0(N389), .A1(n87), .B0(N261), .B1(n85), .Y(n306) );
  MXI2X6 U150 ( .A(n153), .B(n152), .S0(ALUOp_regD[2]), .Y(n154) );
  NAND4BX4 U151 ( .AN(n151), .B(n164), .C(ALUOp_regD[1]), .D(n69), .Y(n153) );
  OAI221X2 U152 ( .A0(n110), .A1(n538), .B0(n537), .B1(n104), .C0(n535), .Y(
        ALUout[31]) );
  OAI221X2 U153 ( .A0(n111), .A1(n358), .B0(n357), .B1(n103), .C0(n356), .Y(
        ALUout[16]) );
  NAND4X4 U154 ( .A(n149), .B(n148), .C(n147), .D(n146), .Y(n155) );
  AOI21X4 U155 ( .A0(n135), .A1(funct_regD[3]), .B0(n134), .Y(n149) );
  OAI221X2 U156 ( .A0(n112), .A1(n219), .B0(n218), .B1(n102), .C0(n217), .Y(
        ALUout[4]) );
  OAI221X2 U157 ( .A0(n110), .A1(n481), .B0(n480), .B1(n104), .C0(n479), .Y(
        ALUout[27]) );
  OAI221X2 U158 ( .A0(n112), .A1(n231), .B0(n230), .B1(n102), .C0(n229), .Y(
        ALUout[5]) );
  NOR4X4 U159 ( .A(n249), .B(n250), .C(n251), .D(n248), .Y(n254) );
  AO22X2 U160 ( .A0(N284), .A1(n82), .B0(N348), .B1(n80), .Y(n204) );
  OAI221X2 U161 ( .A0(n110), .A1(n436), .B0(n435), .B1(n103), .C0(n434), .Y(
        ALUout[23]) );
  NOR4X2 U162 ( .A(n376), .B(n375), .C(n374), .D(n373), .Y(n379) );
  OAI221X2 U163 ( .A0(n110), .A1(n516), .B0(n515), .B1(n104), .C0(n514), .Y(
        ALUout[30]) );
  OAI221X2 U164 ( .A0(n111), .A1(n391), .B0(n390), .B1(n103), .C0(n389), .Y(
        ALUout[19]) );
  OAI221X2 U165 ( .A0(n110), .A1(n413), .B0(n412), .B1(n103), .C0(n411), .Y(
        ALUout[21]) );
  OAI221X1 U166 ( .A0(n111), .A1(n336), .B0(n335), .B1(n103), .C0(n334), .Y(
        ALUout[14]) );
  OAI221X4 U167 ( .A0(n111), .A1(n301), .B0(n300), .B1(n102), .C0(n299), .Y(
        ALUout[11]) );
  AO22X2 U168 ( .A0(N293), .A1(n82), .B0(N357), .B1(n80), .Y(n307) );
  OAI221X2 U169 ( .A0(n111), .A1(n369), .B0(n368), .B1(n103), .C0(n367), .Y(
        ALUout[17]) );
  OAI221X2 U170 ( .A0(n110), .A1(n470), .B0(n469), .B1(n104), .C0(n468), .Y(
        ALUout[26]) );
  NOR4X2 U171 ( .A(n274), .B(n273), .C(n275), .D(n272), .Y(n278) );
  OAI2BB1X4 U172 ( .A0N(N377), .A1N(n88), .B0(n133), .Y(n134) );
  OAI31X4 U173 ( .A0(n127), .A1(funct_regD[0]), .A2(n128), .B0(n138), .Y(n135)
         );
  NOR4X4 U174 ( .A(n530), .B(n529), .C(n528), .D(n527), .Y(n537) );
  NOR4X4 U175 ( .A(n286), .B(n285), .C(n284), .D(n283), .Y(n289) );
  OAI221X2 U176 ( .A0(n112), .A1(n255), .B0(n254), .B1(n102), .C0(n253), .Y(
        ALUout[7]) );
  OAI221X2 U177 ( .A0(n110), .A1(n424), .B0(n423), .B1(n103), .C0(n422), .Y(
        ALUout[22]) );
  NOR4X4 U178 ( .A(n465), .B(n466), .C(n464), .D(n463), .Y(n469) );
  CLKINVX8 U179 ( .A(ALUinB[2]), .Y(n118) );
  NOR4X4 U180 ( .A(n363), .B(n364), .C(n365), .D(n362), .Y(n368) );
  NOR4X4 U181 ( .A(n194), .B(n193), .C(n192), .D(n191), .Y(n198) );
  OAI221X2 U182 ( .A0(n111), .A1(n380), .B0(n379), .B1(n103), .C0(n378), .Y(
        ALUout[18]) );
  NAND4X4 U183 ( .A(n171), .B(n170), .C(n169), .D(n168), .Y(ALUout[0]) );
  AOI21X4 U184 ( .A0(n105), .A1(n155), .B0(n154), .Y(n171) );
  NOR4X4 U185 ( .A(n180), .B(n179), .C(n178), .D(n177), .Y(n186) );
  AO22X2 U186 ( .A0(N378), .A1(n88), .B0(N250), .B1(n84), .Y(n178) );
  NOR4X4 U187 ( .A(n477), .B(n476), .C(n475), .D(n474), .Y(n480) );
  INVX12 U188 ( .A(ALUinB[5]), .Y(n124) );
  INVX16 U189 ( .A(n114), .Y(n113) );
  OAI221X2 U190 ( .A0(n112), .A1(n244), .B0(n243), .B1(n102), .C0(n242), .Y(
        ALUout[6]) );
  OAI221X4 U191 ( .A0(n111), .A1(n279), .B0(n278), .B1(n102), .C0(n277), .Y(
        ALUout[9]) );
  NOR4X4 U192 ( .A(n432), .B(n431), .C(n430), .D(n428), .Y(n435) );
  NOR4X4 U193 ( .A(n420), .B(n419), .C(n418), .D(n417), .Y(n423) );
  NOR4X2 U194 ( .A(n500), .B(n501), .C(n499), .D(n498), .Y(n504) );
  AO22X2 U195 ( .A0(N289), .A1(n82), .B0(N353), .B1(n80), .Y(n262) );
  OAI221X1 U196 ( .A0(n111), .A1(n268), .B0(n267), .B1(n102), .C0(n266), .Y(
        ALUout[8]) );
  OAI221X4 U197 ( .A0(n111), .A1(n290), .B0(n289), .B1(n102), .C0(n288), .Y(
        ALUout[10]) );
  AO22X2 U198 ( .A0(N292), .A1(n82), .B0(N356), .B1(n80), .Y(n296) );
  NOR4X4 U199 ( .A(n205), .B(n204), .C(n203), .D(n202), .Y(n208) );
  AO22X4 U200 ( .A0(N301), .A1(n83), .B0(N365), .B1(n81), .Y(n397) );
  BUFX4 U201 ( .A(n109), .Y(n110) );
  CLKBUFX2 U202 ( .A(n539), .Y(n111) );
  MX2X1 U203 ( .A(n159), .B(n158), .S0(ALUOp_regD[1]), .Y(n161) );
  NAND2XL U204 ( .A(n157), .B(n156), .Y(n159) );
  INVX1 U205 ( .A(n433), .Y(n426) );
  NAND2BX1 U206 ( .AN(n138), .B(n142), .Y(n139) );
  INVX1 U207 ( .A(funct_regD[5]), .Y(n541) );
  NAND2X1 U208 ( .A(funct_regD[1]), .B(n542), .Y(n128) );
  CLKBUFX4 U209 ( .A(n521), .Y(n81) );
  INVX3 U210 ( .A(funct_regD[0]), .Y(n130) );
  NAND2X1 U211 ( .A(ALUOp_regD[3]), .B(n540), .Y(n429) );
  INVX1 U212 ( .A(funct_regD[2]), .Y(n542) );
  CLKMX2X2 U213 ( .A(n78), .B(n75), .S0(n349), .Y(n354) );
  CLKMX2X2 U214 ( .A(n78), .B(n75), .S0(n393), .Y(n398) );
  AO22X2 U215 ( .A0(N298), .A1(n83), .B0(N362), .B1(n80), .Y(n364) );
  CLKMX2X2 U216 ( .A(n78), .B(n75), .S0(n404), .Y(n409) );
  INVX1 U217 ( .A(n490), .Y(n483) );
  INVX1 U218 ( .A(n421), .Y(n415) );
  INVX1 U219 ( .A(n513), .Y(n507) );
  INVX1 U220 ( .A(n502), .Y(n496) );
  INVX1 U221 ( .A(n456), .Y(n450) );
  BUFX2 U222 ( .A(n523), .Y(n87) );
  CLKINVX8 U223 ( .A(ALUinB[0]), .Y(n114) );
  NAND4XL U224 ( .A(funct_regD[3]), .B(funct_regD[0]), .C(n542), .D(n541), .Y(
        n444) );
  INVX4 U225 ( .A(funct_regD[1]), .Y(n136) );
  INVX3 U226 ( .A(n131), .Y(n140) );
  NAND3BX2 U227 ( .AN(funct_regD[3]), .B(funct_regD[5]), .C(n130), .Y(n131) );
  INVXL U228 ( .A(N264), .Y(n347) );
  INVXL U229 ( .A(N263), .Y(n336) );
  INVXL U230 ( .A(N256), .Y(n255) );
  AO22X2 U231 ( .A0(N402), .A1(n86), .B0(N274), .B1(n84), .Y(n453) );
  AO22X2 U232 ( .A0(N398), .A1(n86), .B0(N270), .B1(n84), .Y(n407) );
  CLKMX2X2 U233 ( .A(n78), .B(n75), .S0(n415), .Y(n420) );
  AO22X2 U234 ( .A0(N399), .A1(n86), .B0(N271), .B1(n84), .Y(n418) );
  CLKMX2X2 U235 ( .A(n78), .B(n75), .S0(n360), .Y(n365) );
  AO22X2 U236 ( .A0(N408), .A1(n86), .B0(n84), .B1(N280), .Y(n528) );
  CLKINVX1 U237 ( .A(n399), .Y(n393) );
  CLKINVX1 U238 ( .A(n355), .Y(n349) );
  CLKINVX1 U239 ( .A(n410), .Y(n404) );
  CLKBUFX3 U240 ( .A(n534), .Y(n100) );
  NAND2XL U241 ( .A(n383), .B(n381), .Y(n388) );
  NAND2XL U242 ( .A(n234), .B(n232), .Y(n240) );
  NAND2XL U243 ( .A(n315), .B(n313), .Y(n321) );
  NAND2XL U244 ( .A(n339), .B(n337), .Y(n344) );
  NAND2X2 U245 ( .A(N441), .B(funct_regD[5]), .Y(n127) );
  OAI221X1 U246 ( .A0(n110), .A1(n505), .B0(n504), .B1(n104), .C0(n503), .Y(
        ALUout[29]) );
  NAND2X1 U247 ( .A(n140), .B(n542), .Y(n132) );
  NAND3BX2 U248 ( .AN(n161), .B(n164), .C(n160), .Y(n539) );
  AO22X4 U249 ( .A0(N309), .A1(n83), .B0(N373), .B1(n81), .Y(n488) );
  INVXL U250 ( .A(N255), .Y(n244) );
  INVXL U251 ( .A(N261), .Y(n312) );
  INVXL U252 ( .A(N260), .Y(n301) );
  INVXL U253 ( .A(N258), .Y(n279) );
  INVXL U254 ( .A(N252), .Y(n209) );
  MX2X1 U255 ( .A(n78), .B(n75), .S0(n426), .Y(n432) );
  MX2X1 U256 ( .A(n78), .B(n76), .S0(n450), .Y(n455) );
  INVX1 U257 ( .A(n190), .Y(n196) );
  NAND2BXL U258 ( .AN(n112), .B(N249), .Y(n170) );
  INVX1 U259 ( .A(n478), .Y(n472) );
  INVX1 U260 ( .A(n366), .Y(n360) );
  INVX1 U261 ( .A(n531), .Y(n518) );
  CLKBUFX2 U262 ( .A(n520), .Y(n79) );
  CLKBUFX2 U263 ( .A(n526), .Y(n93) );
  CLKINVX3 U264 ( .A(n105), .Y(n104) );
  CLKBUFX2 U265 ( .A(n519), .Y(n76) );
  CLKBUFX2 U266 ( .A(n534), .Y(n101) );
  CLKBUFX2 U267 ( .A(n532), .Y(n96) );
  NAND2XL U268 ( .A(n189), .B(n118), .Y(n195) );
  INVXL U269 ( .A(ALUinA[1]), .Y(n176) );
  INVXL U270 ( .A(ALUinA[3]), .Y(n201) );
  INVXL U271 ( .A(ALUinA[20]), .Y(n394) );
  INVXL U272 ( .A(ALUinA[16]), .Y(n350) );
  INVXL U273 ( .A(ALUinA[18]), .Y(n372) );
  NAND2BX2 U274 ( .AN(n163), .B(n164), .Y(n182) );
  AOI222XL U275 ( .A0(n101), .A1(n491), .B0(n64), .B1(n533), .C0(n96), .C1(
        n490), .Y(n492) );
  AOI222XL U276 ( .A0(n101), .A1(n59), .B0(n58), .B1(n98), .C0(n96), .C1(n467), 
        .Y(n468) );
  AOI222XL U277 ( .A0(n100), .A1(n42), .B0(n43), .B1(n98), .C0(n95), .C1(n377), 
        .Y(n378) );
  AOI222XL U278 ( .A0(n100), .A1(n45), .B0(n44), .B1(n98), .C0(n95), .C1(n388), 
        .Y(n389) );
  NAND3BXL U279 ( .AN(n542), .B(funct_regD[1]), .C(n140), .Y(n175) );
  NAND2X6 U280 ( .A(funct_regD[0]), .B(n89), .Y(n172) );
  INVX3 U281 ( .A(n137), .Y(n525) );
  NAND3BX2 U282 ( .AN(funct_regD[3]), .B(n136), .C(n70), .Y(n137) );
  INVX4 U283 ( .A(ALUOp_regD[4]), .Y(n164) );
  INVXL U284 ( .A(funct_regD[3]), .Y(n142) );
  NAND3BX2 U285 ( .AN(n163), .B(ALUOp_regD[0]), .C(n164), .Y(n183) );
  NAND4XL U286 ( .A(funct_regD[1]), .B(n70), .C(funct_regD[0]), .D(n142), .Y(
        n173) );
  NAND4X2 U287 ( .A(ALUOp_regD[1]), .B(n72), .C(n69), .D(n164), .Y(n181) );
  INVXL U288 ( .A(ALUOp_regD[1]), .Y(n125) );
  INVX3 U289 ( .A(ALUOp_regD[5]), .Y(n540) );
  INVX3 U290 ( .A(ALUOp_regD[0]), .Y(n157) );
  INVX3 U291 ( .A(n536), .Y(n108) );
  NAND3BX2 U292 ( .AN(funct_regD[4]), .B(n160), .C(n126), .Y(n536) );
  INVX3 U293 ( .A(n152), .Y(n126) );
  INVXL U294 ( .A(ALUOp_regD[3]), .Y(n150) );
  INVXL U295 ( .A(ALUOp_regD[2]), .Y(n160) );
  CLKINVX1 U296 ( .A(N253), .Y(n219) );
  CLKINVX1 U297 ( .A(N250), .Y(n187) );
  CLKINVX1 U298 ( .A(N251), .Y(n199) );
  CLKMX2X2 U299 ( .A(n79), .B(n76), .S0(n483), .Y(n489) );
  CLKMX2X2 U300 ( .A(n79), .B(n76), .S0(n518), .Y(n530) );
  CLKMX2X2 U301 ( .A(n79), .B(n76), .S0(n507), .Y(n512) );
  AO22X1 U302 ( .A0(n93), .A1(n63), .B0(n62), .B1(n89), .Y(n509) );
  AO22X1 U303 ( .A0(N407), .A1(n86), .B0(N279), .B1(n84), .Y(n510) );
  CLKMX2X2 U304 ( .A(n77), .B(n74), .S0(n200), .Y(n205) );
  AO22X1 U305 ( .A0(n91), .A1(n11), .B0(n10), .B1(n90), .Y(n202) );
  CLKMX2X2 U306 ( .A(n77), .B(n74), .S0(n174), .Y(n180) );
  AO22X1 U307 ( .A0(n91), .A1(n8), .B0(n9), .B1(n89), .Y(n177) );
  AO22X1 U308 ( .A0(N282), .A1(n82), .B0(N346), .B1(n80), .Y(n179) );
  CLKMX2X2 U309 ( .A(n78), .B(n75), .S0(n382), .Y(n387) );
  AO22X1 U310 ( .A0(n92), .A1(n45), .B0(n44), .B1(n89), .Y(n384) );
  AO22X1 U311 ( .A0(N300), .A1(n83), .B0(N364), .B1(n81), .Y(n386) );
  CLKMX2X2 U312 ( .A(n77), .B(n74), .S0(n210), .Y(n215) );
  AO22X1 U313 ( .A0(n91), .A1(n31), .B0(n30), .B1(n90), .Y(n212) );
  AO22X1 U314 ( .A0(n92), .A1(n41), .B0(n40), .B1(n89), .Y(n362) );
  AO22X1 U315 ( .A0(n92), .A1(n38), .B0(n39), .B1(n90), .Y(n351) );
  CLKMX2X2 U316 ( .A(n77), .B(n74), .S0(n188), .Y(n194) );
  AO22X1 U317 ( .A0(n91), .A1(n196), .B0(n27), .B1(n90), .Y(n191) );
  AO22X1 U318 ( .A0(n92), .A1(n47), .B0(n46), .B1(n89), .Y(n395) );
  CLKMX2X2 U319 ( .A(n78), .B(n75), .S0(n371), .Y(n376) );
  AO22X1 U320 ( .A0(n92), .A1(n42), .B0(n43), .B1(n89), .Y(n373) );
  AO22X1 U321 ( .A0(N299), .A1(n83), .B0(N363), .B1(n81), .Y(n375) );
  CLKMX2X2 U322 ( .A(n79), .B(n76), .S0(n496), .Y(n501) );
  AO22X1 U323 ( .A0(n93), .A1(n68), .B0(n67), .B1(n89), .Y(n498) );
  CLKMX2X2 U324 ( .A(n78), .B(n75), .S0(n338), .Y(n343) );
  AO22X1 U325 ( .A0(n92), .A1(n37), .B0(n36), .B1(n90), .Y(n340) );
  CLKMX2X2 U326 ( .A(n77), .B(n75), .S0(n314), .Y(n320) );
  AO22X1 U327 ( .A0(n92), .A1(n322), .B0(n33), .B1(n90), .Y(n317) );
  CLKMX2X2 U328 ( .A(n78), .B(n75), .S0(n327), .Y(n332) );
  AO22X1 U329 ( .A0(n92), .A1(n34), .B0(n35), .B1(n90), .Y(n329) );
  CLKMX2X2 U330 ( .A(n78), .B(n76), .S0(n461), .Y(n466) );
  AO22X1 U331 ( .A0(n93), .A1(n59), .B0(n58), .B1(n89), .Y(n463) );
  AO22X1 U332 ( .A0(N403), .A1(n86), .B0(N275), .B1(n84), .Y(n464) );
  CLKMX2X2 U333 ( .A(n79), .B(n76), .S0(n472), .Y(n477) );
  AO22X1 U334 ( .A0(n93), .A1(n61), .B0(n60), .B1(n89), .Y(n474) );
  AO22X1 U335 ( .A0(N404), .A1(n86), .B0(N276), .B1(n84), .Y(n475) );
  AO22X1 U336 ( .A0(n92), .A1(n48), .B0(n49), .B1(n89), .Y(n417) );
  AO22X1 U337 ( .A0(n92), .A1(n56), .B0(n57), .B1(n89), .Y(n406) );
  AO22X1 U338 ( .A0(n93), .A1(n54), .B0(n55), .B1(n89), .Y(n452) );
  AO22X1 U339 ( .A0(n92), .A1(n50), .B0(n51), .B1(n90), .Y(n428) );
  CLKMX2X2 U340 ( .A(n77), .B(n74), .S0(n257), .Y(n263) );
  AO22X1 U341 ( .A0(n91), .A1(n265), .B0(n15), .B1(n90), .Y(n260) );
  CLKMX2X2 U342 ( .A(n77), .B(n74), .S0(n246), .Y(n251) );
  AO22X1 U343 ( .A0(n91), .A1(n13), .B0(n14), .B1(n90), .Y(n248) );
  AO22X1 U344 ( .A0(N288), .A1(n82), .B0(N352), .B1(n80), .Y(n250) );
  CLKMX2X2 U345 ( .A(n77), .B(n74), .S0(n292), .Y(n297) );
  AO22X1 U346 ( .A0(n91), .A1(n18), .B0(n24), .B1(n90), .Y(n294) );
  CLKMX2X2 U347 ( .A(n77), .B(n74), .S0(n220), .Y(n226) );
  AO22X1 U348 ( .A0(n91), .A1(n228), .B0(n12), .B1(n90), .Y(n223) );
  CLKMX2X2 U349 ( .A(n77), .B(n74), .S0(n270), .Y(n275) );
  AO22X1 U350 ( .A0(n91), .A1(n17), .B0(n16), .B1(n90), .Y(n272) );
  CLKMX2X2 U351 ( .A(n77), .B(n74), .S0(n233), .Y(n239) );
  AO22X1 U352 ( .A0(n91), .A1(n241), .B0(n32), .B1(n90), .Y(n236) );
  AO22X1 U353 ( .A0(N287), .A1(n82), .B0(N351), .B1(n80), .Y(n238) );
  CLKMX2X2 U354 ( .A(n77), .B(n74), .S0(n281), .Y(n286) );
  AO22X1 U355 ( .A0(n91), .A1(n28), .B0(n29), .B1(n90), .Y(n283) );
  CLKMX2X2 U356 ( .A(n78), .B(n75), .S0(n438), .Y(n443) );
  AO22X1 U357 ( .A0(n92), .A1(n53), .B0(n52), .B1(n89), .Y(n440) );
  AO22X1 U358 ( .A0(N305), .A1(n83), .B0(N369), .B1(n81), .Y(n442) );
  CLKMX2X2 U359 ( .A(n77), .B(n74), .S0(n303), .Y(n308) );
  AO22X1 U360 ( .A0(n91), .A1(n26), .B0(n25), .B1(n90), .Y(n305) );
  AO22X1 U361 ( .A0(N312), .A1(n83), .B0(N376), .B1(n81), .Y(n529) );
  AO22X1 U362 ( .A0(N390), .A1(n87), .B0(N262), .B1(n85), .Y(n318) );
  AO22X1 U363 ( .A0(N385), .A1(n87), .B0(N257), .B1(n85), .Y(n261) );
  AO22X1 U364 ( .A0(N382), .A1(n88), .B0(N254), .B1(n85), .Y(n224) );
  AO22X1 U365 ( .A0(N383), .A1(n88), .B0(N255), .B1(n85), .Y(n237) );
  AO22X1 U366 ( .A0(N310), .A1(n83), .B0(N374), .B1(n81), .Y(n500) );
  AO22X1 U367 ( .A0(N307), .A1(n83), .B0(N371), .B1(n81), .Y(n465) );
  AO22X1 U368 ( .A0(N308), .A1(n83), .B0(N372), .B1(n81), .Y(n476) );
  AO22X1 U369 ( .A0(N303), .A1(n83), .B0(N367), .B1(n81), .Y(n419) );
  AO22X1 U370 ( .A0(N306), .A1(n83), .B0(N370), .B1(n81), .Y(n454) );
  AO22X1 U371 ( .A0(N401), .A1(n86), .B0(N273), .B1(n84), .Y(n441) );
  AO22X1 U372 ( .A0(N394), .A1(n87), .B0(N266), .B1(n84), .Y(n363) );
  AO22X1 U373 ( .A0(N395), .A1(n87), .B0(N267), .B1(n84), .Y(n374) );
  AO22X1 U374 ( .A0(N393), .A1(n87), .B0(N265), .B1(n85), .Y(n352) );
  XOR2X1 U375 ( .A(n143), .B(n113), .Y(n162) );
  INVX1 U376 ( .A(n222), .Y(n228) );
  XOR2X1 U377 ( .A(n221), .B(n123), .Y(n222) );
  XOR2X1 U378 ( .A(n189), .B(n117), .Y(n190) );
  NAND2BX1 U379 ( .AN(n165), .B(n89), .Y(n148) );
  CLKINVX1 U380 ( .A(n467), .Y(n461) );
  CLKINVX1 U381 ( .A(n388), .Y(n382) );
  CLKINVX1 U382 ( .A(n344), .Y(n338) );
  CLKINVX1 U383 ( .A(n240), .Y(n233) );
  CLKINVX1 U384 ( .A(n227), .Y(n220) );
  CLKINVX1 U385 ( .A(n309), .Y(n303) );
  CLKINVX1 U386 ( .A(n321), .Y(n314) );
  CLKINVX1 U387 ( .A(n377), .Y(n371) );
  CLKINVX1 U388 ( .A(n264), .Y(n257) );
  CLKINVX1 U389 ( .A(n445), .Y(n438) );
  CLKINVX1 U390 ( .A(n252), .Y(n246) );
  CLKINVX1 U391 ( .A(n276), .Y(n270) );
  CLKINVX1 U392 ( .A(n298), .Y(n292) );
  CLKINVX1 U393 ( .A(n287), .Y(n281) );
  CLKINVX1 U394 ( .A(n333), .Y(n327) );
  CLKINVX1 U395 ( .A(n195), .Y(n188) );
  CLKINVX1 U396 ( .A(n216), .Y(n210) );
  CLKINVX1 U397 ( .A(n184), .Y(n174) );
  CLKINVX1 U398 ( .A(n206), .Y(n200) );
  NAND2X1 U399 ( .A(N249), .B(n84), .Y(n133) );
  BUFX4 U400 ( .A(n521), .Y(n80) );
  CLKBUFX3 U401 ( .A(n73), .Y(n82) );
  CLKBUFX3 U402 ( .A(n73), .Y(n83) );
  CLKBUFX3 U403 ( .A(n534), .Y(n99) );
  CLKBUFX3 U404 ( .A(n532), .Y(n95) );
  CLKBUFX3 U405 ( .A(n532), .Y(n94) );
  CLKBUFX3 U406 ( .A(n520), .Y(n78) );
  CLKBUFX3 U407 ( .A(n520), .Y(n77) );
  CLKBUFX3 U408 ( .A(n526), .Y(n91) );
  CLKBUFX3 U409 ( .A(n526), .Y(n92) );
  CLKBUFX3 U410 ( .A(n519), .Y(n75) );
  CLKBUFX3 U411 ( .A(n519), .Y(n74) );
  XOR2XL U412 ( .A(n484), .B(ALUinB[28]), .Y(n485) );
  AOI2BB2X1 U413 ( .B0(N345), .B1(n80), .A0N(n175), .A1N(n162), .Y(n147) );
  INVXL U414 ( .A(ALUinA[28]), .Y(n484) );
  NOR2X1 U415 ( .A(n150), .B(N441), .Y(n151) );
  AOI222XL U416 ( .A0(n100), .A1(n322), .B0(n33), .B1(n98), .C0(n95), .C1(n321), .Y(n323) );
  INVXL U417 ( .A(N262), .Y(n325) );
  AOI222XL U418 ( .A0(n99), .A1(n28), .B0(n29), .B1(n97), .C0(n94), .C1(n287), 
        .Y(n288) );
  INVXL U419 ( .A(N259), .Y(n290) );
  NAND2X1 U420 ( .A(n484), .B(n482), .Y(n490) );
  INVXL U421 ( .A(ALUinB[28]), .Y(n482) );
  INVX1 U422 ( .A(n259), .Y(n265) );
  XOR2XL U423 ( .A(n258), .B(ALUinB[8]), .Y(n259) );
  INVX1 U424 ( .A(n235), .Y(n241) );
  XOR2XL U425 ( .A(n234), .B(ALUinB[6]), .Y(n235) );
  INVX1 U426 ( .A(n316), .Y(n322) );
  XOR2XL U427 ( .A(n315), .B(ALUinB[13]), .Y(n316) );
  INVXL U428 ( .A(ALUinA[9]), .Y(n271) );
  INVXL U429 ( .A(ALUinA[30]), .Y(n508) );
  NAND2XL U430 ( .A(n221), .B(n124), .Y(n227) );
  NAND2X1 U431 ( .A(n304), .B(n302), .Y(n309) );
  INVXL U432 ( .A(ALUinB[12]), .Y(n302) );
  INVXL U433 ( .A(ALUinB[13]), .Y(n313) );
  INVXL U434 ( .A(ALUinA[4]), .Y(n211) );
  NAND2X1 U435 ( .A(n293), .B(n291), .Y(n298) );
  INVXL U436 ( .A(ALUinB[11]), .Y(n291) );
  NAND2X1 U437 ( .A(n524), .B(n517), .Y(n531) );
  INVXL U438 ( .A(ALUinB[31]), .Y(n517) );
  NAND2X1 U439 ( .A(n176), .B(n116), .Y(n184) );
  INVXL U440 ( .A(ALUinA[22]), .Y(n416) );
  INVXL U441 ( .A(ALUinA[11]), .Y(n293) );
  INVXL U442 ( .A(ALUinA[21]), .Y(n405) );
  INVXL U443 ( .A(ALUinA[10]), .Y(n282) );
  INVXL U444 ( .A(ALUinA[23]), .Y(n427) );
  INVXL U445 ( .A(ALUinA[14]), .Y(n328) );
  INVXL U446 ( .A(ALUinA[25]), .Y(n451) );
  INVXL U447 ( .A(ALUinA[31]), .Y(n524) );
  INVXL U448 ( .A(ALUinA[27]), .Y(n473) );
  INVXL U449 ( .A(ALUinA[7]), .Y(n247) );
  INVXL U450 ( .A(ALUinA[2]), .Y(n189) );
  NAND2X1 U451 ( .A(n497), .B(n495), .Y(n502) );
  INVXL U452 ( .A(ALUinB[29]), .Y(n495) );
  NAND2X1 U453 ( .A(n361), .B(n359), .Y(n366) );
  INVXL U454 ( .A(ALUinB[17]), .Y(n359) );
  NAND2X1 U455 ( .A(n258), .B(n256), .Y(n264) );
  INVXL U456 ( .A(ALUinB[8]), .Y(n256) );
  NAND2X1 U457 ( .A(n439), .B(n437), .Y(n445) );
  INVXL U458 ( .A(ALUinB[24]), .Y(n437) );
  NAND2X1 U459 ( .A(n394), .B(n392), .Y(n399) );
  INVXL U460 ( .A(ALUinB[20]), .Y(n392) );
  NAND2X1 U461 ( .A(n350), .B(n348), .Y(n355) );
  INVXL U462 ( .A(ALUinB[16]), .Y(n348) );
  NAND2X1 U463 ( .A(n372), .B(n370), .Y(n377) );
  INVXL U464 ( .A(ALUinB[18]), .Y(n370) );
  NAND2X1 U465 ( .A(n416), .B(n414), .Y(n421) );
  INVXL U466 ( .A(ALUinB[22]), .Y(n414) );
  NAND2X1 U467 ( .A(n247), .B(n245), .Y(n252) );
  INVXL U468 ( .A(ALUinB[7]), .Y(n245) );
  NAND2X1 U469 ( .A(n508), .B(n506), .Y(n513) );
  INVXL U470 ( .A(ALUinB[30]), .Y(n506) );
  NAND2X1 U471 ( .A(n271), .B(n269), .Y(n276) );
  INVXL U472 ( .A(ALUinB[9]), .Y(n269) );
  INVXL U473 ( .A(ALUinB[6]), .Y(n232) );
  NAND2X1 U474 ( .A(n427), .B(n425), .Y(n433) );
  INVXL U475 ( .A(ALUinB[23]), .Y(n425) );
  NAND2X1 U476 ( .A(n451), .B(n449), .Y(n456) );
  INVXL U477 ( .A(ALUinB[25]), .Y(n449) );
  NAND2X1 U478 ( .A(n328), .B(n326), .Y(n333) );
  INVXL U479 ( .A(ALUinB[14]), .Y(n326) );
  NAND2X1 U480 ( .A(n405), .B(n403), .Y(n410) );
  INVXL U481 ( .A(ALUinB[21]), .Y(n403) );
  NAND2X1 U482 ( .A(n282), .B(n280), .Y(n287) );
  INVXL U483 ( .A(ALUinB[10]), .Y(n280) );
  NAND2X1 U484 ( .A(n473), .B(n471), .Y(n478) );
  INVXL U485 ( .A(ALUinB[27]), .Y(n471) );
  NAND2X1 U486 ( .A(n462), .B(n460), .Y(n467) );
  INVXL U487 ( .A(ALUinB[26]), .Y(n460) );
  INVXL U488 ( .A(ALUinB[19]), .Y(n381) );
  INVXL U489 ( .A(ALUinB[15]), .Y(n337) );
  NOR2BX1 U490 ( .AN(n145), .B(n144), .Y(n146) );
  NAND2X1 U491 ( .A(N281), .B(n82), .Y(n145) );
  MXI2X1 U492 ( .A(n172), .B(n173), .S0(n71), .Y(n144) );
  INVXL U493 ( .A(ALUinA[29]), .Y(n497) );
  CLKINVX1 U494 ( .A(ALUinA[17]), .Y(n361) );
  CLKINVX1 U495 ( .A(ALUinA[8]), .Y(n258) );
  INVXL U496 ( .A(ALUinA[24]), .Y(n439) );
  NOR2X1 U497 ( .A(n167), .B(n166), .Y(n168) );
  NOR2XL U498 ( .A(n183), .B(n71), .Y(n167) );
  NOR2XL U499 ( .A(n165), .B(n182), .Y(n166) );
  NAND4X1 U500 ( .A(n541), .B(n542), .C(n136), .D(n130), .Y(n138) );
  CLKINVX1 U501 ( .A(n128), .Y(n141) );
  CLKBUFX3 U502 ( .A(n525), .Y(n89) );
  CLKBUFX3 U503 ( .A(n522), .Y(n84) );
  CLKBUFX3 U504 ( .A(n525), .Y(n90) );
  CLKBUFX3 U505 ( .A(n522), .Y(n85) );
  CLKBUFX3 U506 ( .A(n108), .Y(n105) );
  CLKINVX1 U507 ( .A(n429), .Y(n156) );
  INVX3 U508 ( .A(n107), .Y(n102) );
  CLKBUFX3 U509 ( .A(n108), .Y(n107) );
  INVX3 U510 ( .A(n106), .Y(n103) );
  CLKBUFX3 U511 ( .A(n108), .Y(n106) );
  BUFX2 U512 ( .A(n523), .Y(n88) );
  CLKBUFX3 U513 ( .A(n109), .Y(n112) );
  CLKBUFX3 U514 ( .A(n539), .Y(n109) );
  INVXL U515 ( .A(N277), .Y(n494) );
  AOI222XL U516 ( .A0(n100), .A1(n53), .B0(n52), .B1(n98), .C0(n95), .C1(n445), 
        .Y(n446) );
  INVXL U517 ( .A(N273), .Y(n448) );
  AOI222XL U518 ( .A0(n99), .A1(n265), .B0(n15), .B1(n97), .C0(n94), .C1(n264), 
        .Y(n266) );
  INVXL U519 ( .A(N257), .Y(n268) );
  AOI222XL U520 ( .A0(n99), .A1(n228), .B0(n12), .B1(n97), .C0(n94), .C1(n227), 
        .Y(n229) );
  INVXL U521 ( .A(N254), .Y(n231) );
  AOI222XL U522 ( .A0(n99), .A1(n8), .B0(n9), .B1(n97), .C0(n94), .C1(n184), 
        .Y(n185) );
  AOI222XL U523 ( .A0(n99), .A1(n196), .B0(n27), .B1(n97), .C0(n94), .C1(n195), 
        .Y(n197) );
  AOI222XL U524 ( .A0(n99), .A1(n11), .B0(n10), .B1(n97), .C0(n94), .C1(n206), 
        .Y(n207) );
  AOI222XL U525 ( .A0(n99), .A1(n31), .B0(n30), .B1(n97), .C0(n94), .C1(n216), 
        .Y(n217) );
  AOI222XL U526 ( .A0(n99), .A1(n241), .B0(n32), .B1(n97), .C0(n94), .C1(n240), 
        .Y(n242) );
  AOI222XL U527 ( .A0(n99), .A1(n13), .B0(n14), .B1(n97), .C0(n94), .C1(n252), 
        .Y(n253) );
  AOI222XL U528 ( .A0(n99), .A1(n17), .B0(n16), .B1(n97), .C0(n94), .C1(n276), 
        .Y(n277) );
  AOI222XL U529 ( .A0(n99), .A1(n18), .B0(n24), .B1(n97), .C0(n94), .C1(n298), 
        .Y(n299) );
  AOI222XL U530 ( .A0(n99), .A1(n26), .B0(n25), .B1(n97), .C0(n94), .C1(n309), 
        .Y(n310) );
  AOI222XL U531 ( .A0(n100), .A1(n34), .B0(n35), .B1(n98), .C0(n95), .C1(n333), 
        .Y(n334) );
  AOI222XL U532 ( .A0(n100), .A1(n37), .B0(n36), .B1(n98), .C0(n95), .C1(n344), 
        .Y(n345) );
  OR2XL U533 ( .A(n162), .B(n181), .Y(n169) );
  OAI221X1 U534 ( .A0(n110), .A1(n402), .B0(n401), .B1(n103), .C0(n400), .Y(
        ALUout[20]) );
  AOI222XL U535 ( .A0(n100), .A1(n47), .B0(n46), .B1(n98), .C0(n95), .C1(n399), 
        .Y(n400) );
  INVXL U536 ( .A(N269), .Y(n402) );
  INVXL U537 ( .A(N268), .Y(n391) );
  AOI222XL U538 ( .A0(n101), .A1(n68), .B0(n67), .B1(n533), .C0(n96), .C1(n502), .Y(n503) );
  INVXL U539 ( .A(N278), .Y(n505) );
  AOI222XL U540 ( .A0(n101), .A1(n63), .B0(n62), .B1(n533), .C0(n96), .C1(n513), .Y(n514) );
  INVXL U541 ( .A(N279), .Y(n516) );
  AOI222XL U542 ( .A0(n101), .A1(n65), .B0(n66), .B1(n533), .C0(n96), .C1(n531), .Y(n535) );
  INVXL U543 ( .A(N280), .Y(n538) );
  AOI222XL U544 ( .A0(n100), .A1(n41), .B0(n40), .B1(n98), .C0(n95), .C1(n366), 
        .Y(n367) );
  INVXL U545 ( .A(N266), .Y(n369) );
  INVXL U546 ( .A(N275), .Y(n470) );
  AOI222XL U547 ( .A0(n101), .A1(n61), .B0(n60), .B1(n533), .C0(n96), .C1(n478), .Y(n479) );
  INVXL U548 ( .A(N276), .Y(n481) );
  AOI222XL U549 ( .A0(n100), .A1(n48), .B0(n49), .B1(n98), .C0(n95), .C1(n421), 
        .Y(n422) );
  AOI222XL U550 ( .A0(n100), .A1(n56), .B0(n57), .B1(n98), .C0(n95), .C1(n410), 
        .Y(n411) );
  INVXL U551 ( .A(N270), .Y(n413) );
  OAI221X1 U552 ( .A0(n110), .A1(n459), .B0(n458), .B1(n104), .C0(n457), .Y(
        ALUout[25]) );
  AOI222XL U553 ( .A0(n101), .A1(n54), .B0(n55), .B1(n97), .C0(n96), .C1(n456), 
        .Y(n457) );
  INVXL U554 ( .A(N274), .Y(n459) );
  AOI222XL U555 ( .A0(n100), .A1(n50), .B0(n51), .B1(n98), .C0(n95), .C1(n433), 
        .Y(n434) );
  INVXL U556 ( .A(N272), .Y(n436) );
  INVXL U557 ( .A(N267), .Y(n380) );
  AOI222XL U558 ( .A0(n100), .A1(n38), .B0(n39), .B1(n98), .C0(n95), .C1(n355), 
        .Y(n356) );
  INVXL U559 ( .A(N265), .Y(n358) );
  NAND2XL U560 ( .A(n429), .B(ALUOp_regD[0]), .Y(n158) );
  INVXL U561 ( .A(ALUinA[13]), .Y(n315) );
  INVXL U562 ( .A(ALUinA[26]), .Y(n462) );
  INVXL U563 ( .A(ALUinA[12]), .Y(n304) );
  INVXL U564 ( .A(ALUinA[19]), .Y(n383) );
  INVXL U565 ( .A(ALUinA[6]), .Y(n234) );
  NAND2XL U566 ( .A(n113), .B(ALUinA[0]), .Y(n165) );
  INVXL U567 ( .A(ALUinA[0]), .Y(n143) );
  INVXL U568 ( .A(ALUinA[5]), .Y(n221) );
  INVXL U569 ( .A(ALUinA[15]), .Y(n339) );
  CLKINVX3 U570 ( .A(n129), .Y(n523) );
  CLKINVX3 U571 ( .A(n139), .Y(n521) );
  NAND3BX2 U572 ( .AN(ALUOp_regD[1]), .B(n540), .C(n72), .Y(n163) );
  CLKINVX3 U573 ( .A(n172), .Y(n520) );
  CLKINVX3 U574 ( .A(n181), .Y(n534) );
  CLKINVX3 U575 ( .A(n183), .Y(n532) );
  AO22X4 U576 ( .A0(N405), .A1(n86), .B0(N277), .B1(n84), .Y(n487) );
endmodule


module MIPS_Pipeline_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n28, n29, n31, n32, n33,
         n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n50, n51, n52, n53, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65,
         n67, n68, n69, n70, n71, n74, n75, n76, n77, n78, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98,
         n99, n100, n102, n103, n104, n106, n107, n108, n109, n110, n112, n113,
         n114, n115, n116, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n138,
         n139, n140, n142, n144, n145, n146, n147, n149, n150, n152, n153,
         n154, n155, n156, n260, n261, n262;
  assign n7 = A[30];
  assign n14 = A[29];
  assign n19 = A[28];
  assign n26 = A[27];
  assign n31 = A[26];
  assign n38 = A[25];
  assign n43 = A[24];
  assign n50 = A[23];
  assign n55 = A[22];
  assign n62 = A[21];
  assign n67 = A[20];
  assign n74 = A[19];
  assign n77 = A[18];
  assign n83 = A[17];
  assign n88 = A[16];
  assign n95 = A[15];
  assign n100 = A[14];
  assign n107 = A[13];
  assign n112 = A[12];
  assign n119 = A[11];
  assign n122 = A[10];
  assign n128 = A[9];
  assign n132 = A[8];
  assign n138 = A[7];
  assign n142 = A[6];
  assign n147 = A[5];
  assign n150 = A[4];
  assign n154 = A[3];
  assign n156 = A[2];

  XNOR2X4 U146 ( .A(n130), .B(n129), .Y(SUM[9]) );
  XNOR2X4 U158 ( .A(n140), .B(n139), .Y(SUM[7]) );
  NOR2X8 U172 ( .A(n146), .B(n153), .Y(n145) );
  NOR2X2 U191 ( .A(n116), .B(n106), .Y(n103) );
  NOR2X1 U192 ( .A(n71), .B(n61), .Y(n58) );
  XOR2X1 U193 ( .A(n114), .B(n113), .Y(SUM[12]) );
  XNOR2X2 U194 ( .A(n134), .B(n133), .Y(SUM[8]) );
  XNOR2X2 U195 ( .A(n124), .B(n123), .Y(SUM[10]) );
  XOR2X2 U196 ( .A(n144), .B(n262), .Y(SUM[6]) );
  INVX1 U197 ( .A(n156), .Y(SUM[2]) );
  XNOR2X2 U198 ( .A(n155), .B(n156), .Y(SUM[3]) );
  INVXL U199 ( .A(n147), .Y(n261) );
  NAND2X4 U200 ( .A(n77), .B(n74), .Y(n71) );
  NAND2X4 U201 ( .A(n154), .B(n156), .Y(n153) );
  NOR2X6 U202 ( .A(n125), .B(n80), .Y(n1) );
  CLKINVX2 U203 ( .A(n125), .Y(n124) );
  NAND2X4 U204 ( .A(n103), .B(n81), .Y(n80) );
  INVXL U205 ( .A(n116), .Y(n115) );
  NAND2X1 U206 ( .A(n124), .B(n115), .Y(n114) );
  NAND2XL U207 ( .A(n150), .B(n152), .Y(n149) );
  INVXL U208 ( .A(n150), .Y(n260) );
  INVXL U209 ( .A(n135), .Y(n136) );
  INVXL U210 ( .A(n58), .Y(n59) );
  NOR2XL U211 ( .A(n104), .B(n87), .Y(n86) );
  NOR2XL U212 ( .A(n104), .B(n99), .Y(n98) );
  INVXL U213 ( .A(n47), .Y(n48) );
  INVX1 U214 ( .A(n145), .Y(n144) );
  XOR2X4 U215 ( .A(n149), .B(n261), .Y(SUM[5]) );
  NOR2X2 U216 ( .A(n92), .B(n82), .Y(n81) );
  NAND2X4 U217 ( .A(n150), .B(n147), .Y(n146) );
  INVXL U218 ( .A(n103), .Y(n104) );
  INVXL U219 ( .A(n153), .Y(n152) );
  NAND2XL U220 ( .A(n124), .B(n103), .Y(n102) );
  INVX1 U221 ( .A(n12), .Y(n11) );
  INVXL U222 ( .A(n142), .Y(n262) );
  NOR2XL U223 ( .A(n59), .B(n56), .Y(n53) );
  NAND2X1 U224 ( .A(n58), .B(n36), .Y(n2) );
  NOR2XL U225 ( .A(n59), .B(n47), .Y(n46) );
  NOR2X4 U226 ( .A(n135), .B(n127), .Y(n126) );
  NOR2XL U227 ( .A(n2), .B(n6), .Y(n5) );
  NOR2XL U228 ( .A(n144), .B(n135), .Y(n134) );
  NOR2X1 U229 ( .A(n144), .B(n262), .Y(n140) );
  NAND2XL U230 ( .A(n124), .B(n91), .Y(n90) );
  NOR2XL U231 ( .A(n104), .B(n92), .Y(n91) );
  NOR2X1 U232 ( .A(n144), .B(n131), .Y(n130) );
  XNOR2X1 U233 ( .A(n260), .B(n152), .Y(SUM[4]) );
  XOR2X1 U234 ( .A(n69), .B(n68), .Y(SUM[20]) );
  NAND2X1 U235 ( .A(n1), .B(n70), .Y(n69) );
  INVXL U236 ( .A(n71), .Y(n70) );
  XOR2X1 U237 ( .A(n57), .B(n56), .Y(SUM[22]) );
  NAND2XL U238 ( .A(n1), .B(n58), .Y(n57) );
  XOR2X1 U239 ( .A(n33), .B(n32), .Y(SUM[26]) );
  NAND2XL U240 ( .A(n1), .B(n34), .Y(n33) );
  CLKINVX1 U241 ( .A(n2), .Y(n34) );
  XOR2X4 U242 ( .A(n102), .B(n99), .Y(SUM[14]) );
  NAND2X1 U243 ( .A(n122), .B(n119), .Y(n116) );
  INVXL U244 ( .A(n122), .Y(n123) );
  NAND2XL U245 ( .A(n112), .B(n107), .Y(n106) );
  NAND2X6 U246 ( .A(n145), .B(n126), .Y(n125) );
  NAND2XL U247 ( .A(n132), .B(n128), .Y(n127) );
  XOR2X4 U248 ( .A(n109), .B(n108), .Y(SUM[13]) );
  INVXL U249 ( .A(n107), .Y(n108) );
  NAND2X1 U250 ( .A(n124), .B(n110), .Y(n109) );
  NOR2X1 U251 ( .A(n116), .B(n113), .Y(n110) );
  XOR2X4 U252 ( .A(n90), .B(n89), .Y(SUM[16]) );
  INVXL U253 ( .A(n88), .Y(n89) );
  XOR2X4 U254 ( .A(n121), .B(n120), .Y(SUM[11]) );
  INVXL U255 ( .A(n119), .Y(n120) );
  NAND2XL U256 ( .A(n124), .B(n122), .Y(n121) );
  XOR2X4 U257 ( .A(n97), .B(n96), .Y(SUM[15]) );
  INVXL U258 ( .A(n95), .Y(n96) );
  NAND2XL U259 ( .A(n124), .B(n98), .Y(n97) );
  INVXL U260 ( .A(n154), .Y(n155) );
  INVXL U261 ( .A(n67), .Y(n68) );
  INVXL U262 ( .A(n55), .Y(n56) );
  INVXL U263 ( .A(n31), .Y(n32) );
  INVXL U264 ( .A(n112), .Y(n113) );
  NAND2XL U265 ( .A(n55), .B(n50), .Y(n47) );
  NAND2XL U266 ( .A(n31), .B(n26), .Y(n23) );
  INVXL U267 ( .A(n100), .Y(n99) );
  INVXL U268 ( .A(n132), .Y(n133) );
  XNOR2X1 U269 ( .A(n1), .B(n78), .Y(SUM[18]) );
  INVXL U270 ( .A(n77), .Y(n78) );
  NAND2XL U271 ( .A(n100), .B(n95), .Y(n92) );
  INVXL U272 ( .A(n128), .Y(n129) );
  NAND2XL U273 ( .A(n136), .B(n132), .Y(n131) );
  INVXL U274 ( .A(n138), .Y(n139) );
  NOR2X1 U275 ( .A(n47), .B(n37), .Y(n36) );
  NAND2XL U276 ( .A(n43), .B(n38), .Y(n37) );
  NAND2X1 U277 ( .A(n142), .B(n138), .Y(n135) );
  NAND2XL U278 ( .A(n88), .B(n83), .Y(n82) );
  NAND2BXL U279 ( .AN(n23), .B(n19), .Y(n18) );
  NAND2XL U280 ( .A(n48), .B(n43), .Y(n42) );
  NAND2XL U281 ( .A(n67), .B(n62), .Y(n61) );
  NAND2XL U282 ( .A(n12), .B(n7), .Y(n6) );
  NOR2X1 U283 ( .A(n23), .B(n13), .Y(n12) );
  NAND2XL U284 ( .A(n19), .B(n14), .Y(n13) );
  NAND2XL U285 ( .A(n93), .B(n88), .Y(n87) );
  INVXL U286 ( .A(n92), .Y(n93) );
  XOR2X1 U287 ( .A(n21), .B(n20), .Y(SUM[28]) );
  INVXL U288 ( .A(n19), .Y(n20) );
  NAND2XL U289 ( .A(n1), .B(n22), .Y(n21) );
  NOR2X1 U290 ( .A(n2), .B(n23), .Y(n22) );
  XOR2X1 U291 ( .A(n16), .B(n15), .Y(SUM[29]) );
  INVXL U292 ( .A(n14), .Y(n15) );
  NAND2XL U293 ( .A(n1), .B(n17), .Y(n16) );
  NOR2X1 U294 ( .A(n2), .B(n18), .Y(n17) );
  XOR2X1 U295 ( .A(n9), .B(n8), .Y(SUM[30]) );
  INVXL U296 ( .A(n7), .Y(n8) );
  NAND2XL U297 ( .A(n1), .B(n10), .Y(n9) );
  NOR2X1 U298 ( .A(n2), .B(n11), .Y(n10) );
  XOR2X4 U299 ( .A(n45), .B(n44), .Y(SUM[24]) );
  INVXL U300 ( .A(n43), .Y(n44) );
  NAND2XL U301 ( .A(n1), .B(n46), .Y(n45) );
  XOR2X1 U302 ( .A(n28), .B(n27), .Y(SUM[27]) );
  INVXL U303 ( .A(n26), .Y(n27) );
  NAND2XL U304 ( .A(n1), .B(n29), .Y(n28) );
  NOR2X1 U305 ( .A(n2), .B(n32), .Y(n29) );
  XOR2X4 U306 ( .A(n85), .B(n84), .Y(SUM[17]) );
  INVXL U307 ( .A(n83), .Y(n84) );
  NAND2XL U308 ( .A(n124), .B(n86), .Y(n85) );
  XOR2X4 U309 ( .A(n52), .B(n51), .Y(SUM[23]) );
  INVXL U310 ( .A(n50), .Y(n51) );
  NAND2XL U311 ( .A(n1), .B(n53), .Y(n52) );
  XOR2X4 U312 ( .A(n64), .B(n63), .Y(SUM[21]) );
  INVXL U313 ( .A(n62), .Y(n63) );
  NAND2XL U314 ( .A(n1), .B(n65), .Y(n64) );
  NOR2XL U315 ( .A(n71), .B(n68), .Y(n65) );
  XOR2X1 U316 ( .A(n40), .B(n39), .Y(SUM[25]) );
  INVXL U317 ( .A(n38), .Y(n39) );
  NAND2X1 U318 ( .A(n1), .B(n41), .Y(n40) );
  NOR2X1 U319 ( .A(n59), .B(n42), .Y(n41) );
  XOR2X1 U320 ( .A(n76), .B(n75), .Y(SUM[19]) );
  INVXL U321 ( .A(n74), .Y(n75) );
  NAND2XL U322 ( .A(n1), .B(n77), .Y(n76) );
  XOR2X1 U323 ( .A(n4), .B(n3), .Y(SUM[31]) );
  INVXL U324 ( .A(A[31]), .Y(n3) );
  NAND2XL U325 ( .A(n1), .B(n5), .Y(n4) );
  CLKBUFX3 U326 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U327 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, flush, stallcache, stall_lw_use, JumpReg_m,
         MemRead_m, MemWrite_m, ALUsrc, RegWrite_m, Branch_DEC_m, MemRead_regD,
         MemWrite_regD, ALUsrc_regD, RegWrite_regD, JumpReg_regD, Branch_regD,
         RegWrite_regE, RegWrite_regM, Branch_DEC, MemRead, MemWrite, RegWrite,
         JumpReg, ExtOp, pred_cond, Jump_IF, Branch_IF, n52, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n103, n104, n105, n106, n107, n108, n109, n111, n112,
         n113, n114, n115, n116, n117, n119, n120, n122, n123, n126, n127,
         n128, n144, n145, n146, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241;
  wire   [31:0] PCplus4;
  wire   [15:0] branchOffset_D;
  wire   [5:0] opcode;
  wire   [4:0] Rs;
  wire   [4:0] Rt;
  wire   [4:0] Rd;
  wire   [4:0] shamt;
  wire   [5:0] funct;
  wire   [15:0] immediate;
  wire   [31:0] PCplus4_regI;
  wire   [1:0] MemtoReg;
  wire   [5:0] ALUOp;
  wire   [31:0] A_f;
  wire   [31:0] B_f;
  wire   [31:0] ExtOut;
  wire   [4:0] wsel;
  wire   [1:0] MemtoReg_regD;
  wire   [5:0] ALUOp_regD;
  wire   [5:0] funct_regD;
  wire   [31:0] A_regD;
  wire   [31:0] B_regD;
  wire   [31:0] ExtOut_regD;
  wire   [4:0] Rs_regD;
  wire   [4:0] Rt_regD;
  wire   [4:0] wsel_regD;
  wire   [31:0] PCplus4_regD;
  wire   [15:0] branchOffset_regD;
  wire   [31:0] tempALUinB;
  wire   [31:0] ALUout;
  wire   [1:0] MemtoReg_regE;
  wire   [4:0] wsel_regE;
  wire   [1:0] ALUout_regE;
  wire   [1:0] MemtoReg_regM;
  wire   [31:0] ALUout_regM;
  wire   [4:0] wsel_regM;
  wire   [31:0] dataOut_regM;
  wire   [1:0] RegDst;
  wire   [31:0] WriteData;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [1:0] FU_Asel;
  wire   [31:0] ALUinA;
  wire   [1:0] FU_Bsel;
  wire   [1:0] PCcur;
  wire   [2:0] PCsrc;
  wire   [31:0] PCnext;
  wire   [31:0] ALUinB;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;

  DFFRX4 \PCreg_reg[3]  ( .D(PCnext[3]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[1]) );
  DFFRX4 \PCreg_reg[4]  ( .D(PCnext[4]), .CK(clk), .RN(ICACHE_ren), .Q(n39), 
        .QN(n60) );
  DFFRX4 \PCreg_reg[5]  ( .D(PCnext[5]), .CK(clk), .RN(ICACHE_ren), .Q(n242), 
        .QN(n101) );
  IF_DEC_regFile i_IF_DEC_regFile ( .clk(clk), .rst_n(n186), .flush(n72), 
        .stallcache(n181), .stall_lw_use(stall_lw_use), .instruction_next({n78, 
        n76, n144, n126, n71, ICACHE_rdata[26:10], n35, ICACHE_rdata[8:6], n48, 
        ICACHE_rdata[4:0]}), .PCplus4(PCplus4), .branchOffset(branchOffset_D), 
        .opcode(opcode), .Rs(Rs), .Rt(Rt), .Rd(Rd), .shamt(shamt), .funct(
        funct), .immediate(immediate), .PCplus4_regI(PCplus4_regI) );
  DEC_EX_regFile i_DEC_EX_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(n181), .MemtoReg(MemtoReg), .ALUOp(ALUOp), .JumpReg(
        JumpReg_m), .MemRead(MemRead_m), .MemWrite(MemWrite_m), .ALUsrc(ALUsrc), .RegWrite(RegWrite_m), .Branch(Branch_DEC_m), .PCplus4_regI(PCplus4_regI), 
        .funct(funct), .branchOffset_D(branchOffset_D), .A(A_f), .B(B_f), 
        .ExtOut(ExtOut), .Rs({n180, n179, n178, n177, n176}), .Rt({n175, n174, 
        n173, n172, n171}), .wsel(wsel), .MemtoReg_regD(MemtoReg_regD), 
        .ALUOp_regD(ALUOp_regD), .MemRead_regD(MemRead_regD), .MemWrite_regD(
        MemWrite_regD), .ALUsrc_regD(ALUsrc_regD), .RegWrite_regD(
        RegWrite_regD), .funct_regD(funct_regD), .A_regD(A_regD), .B_regD(
        B_regD), .ExtOut_regD(ExtOut_regD), .Rs_regD(Rs_regD), .Rt_regD(
        Rt_regD), .wsel_regD(wsel_regD), .JumpReg_regD(JumpReg_regD), 
        .Branch_regD(Branch_regD), .PCplus4_regD(PCplus4_regD), 
        .branchOffset_regD(branchOffset_regD) );
  EX_MEM_regFile i_EX_MEM_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(n181), .MemtoReg_regD(MemtoReg_regD), .MemRead_regD(
        MemRead_regD), .MemWrite_regD(MemWrite_regD), .RegWrite_regD(
        RegWrite_regD), .B_regD({tempALUinB[31:30], n53, tempALUinB[28:13], 
        n51, tempALUinB[11:7], n62, tempALUinB[5:0]}), .wsel_regD(wsel_regD), 
        .ALUout(ALUout), .MemtoReg_regE(MemtoReg_regE), .MemRead_regE(
        DCACHE_ren), .MemWrite_regE(DCACHE_wen), .RegWrite_regE(RegWrite_regE), 
        .B_regE(DCACHE_wdata), .wsel_regE(wsel_regE), .ALUout_regE({n243, n244, 
        n245, DCACHE_addr[26], n246, n247, n248, DCACHE_addr[22], n249, n250, 
        n251, n252, n253, n254, n255, n256, n257, n258, DCACHE_addr[11], n259, 
        n260, DCACHE_addr[8], n261, n262, n263, n264, n265, n266, n267, 
        DCACHE_addr[0], ALUout_regE}) );
  MEM_WB_regFile i_MEM_WB_regFile ( .clk(clk), .rst_n(n186), .stallcache(n181), 
        .MemtoReg_regE(MemtoReg_regE), .RegWrite_regE(RegWrite_regE), 
        .ALUout_regE({DCACHE_addr, ALUout_regE}), .wsel_regE(wsel_regE), 
        .dataOut(DCACHE_rdata), .MemtoReg_regM(MemtoReg_regM), .RegWrite_regM(
        RegWrite_regM), .ALUout_regM(ALUout_regM), .wsel_regM(wsel_regM), 
        .dataOut_regM(dataOut_regM) );
  maincontrol i_maincontrol ( .opcode(opcode), .funct(funct), .RegDst(RegDst), 
        .MemtoReg(MemtoReg), .ALUOp(ALUOp), .Branch(Branch_DEC), .MemRead(
        MemRead), .MemWrite(MemWrite), .ALUsrc(ALUsrc), .RegWrite(RegWrite), 
        .JumpReg(JumpReg), .ExtOp(ExtOp) );
  registerFile i_registrefFile ( .clk(clk), .rst_n(n186), .rsel1({n180, n179, 
        n178, n177, n176}), .rsel2({n175, n174, n173, n172, n171}), .wsel({n47, 
        n59, n88, n94, n82}), .wen(RegWrite_regM), .wdata({WriteData[31:4], 
        n42, WriteData[2:0]}), .rdata1(A), .rdata2(B) );
  extender i_extender ( .shamt_i(shamt), .immed_i(immediate), .ExtOp_i(ExtOp), 
        .ExtOut_o(ExtOut) );
  MUX_5_3to1 MUX_wsel ( .data0_i({n175, n174, n173, n172, n171}), .data1_i(Rd), 
        .data2_i({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .select_i(RegDst), .data_o(
        wsel) );
  MUX_32_3to1_0 MUX_WriteData ( .data0_i(dataOut_regM), .data1_i(ALUout_regM), 
        .data2_i(ALUout_regM), .select_i(MemtoReg_regM), .data_o(WriteData) );
  MUX_32_3to1_2 MUX_ALUinA ( .data0_i(A_regD), .data1_i(WriteData), .data2_i({
        DCACHE_addr[29:28], n245, DCACHE_addr[26:19], n252, n253, 
        DCACHE_addr[16:14], n257, DCACHE_addr[12:11], n259, DCACHE_addr[9:7], 
        n262, DCACHE_addr[5:0], ALUout_regE}), .select_i(FU_Asel), .data_o(
        ALUinA) );
  MUX_32_3to1_1 MUX_ALUinB ( .data0_i(B_regD), .data1_i(WriteData), .data2_i({
        DCACHE_addr[29:14], n257, DCACHE_addr[12:0], ALUout_regE}), .select_i(
        FU_Bsel), .data_o(tempALUinB) );
  forwarding i_forwarding ( .Rs_regD(Rs_regD), .Rt_regD(Rt_regD), 
        .RegWrite_regE(RegWrite_regE), .wsel_regE(wsel_regE), .RegWrite_regM(
        RegWrite_regM), .wsel_regM(wsel_regM), .FU_Asel(FU_Asel), .FU_Bsel(
        FU_Bsel) );
  hazard_detection i_hazard_detection ( .Branch_EX(Branch_regD), .equal(n40), 
        .branchpred_his(1'b0), .JumpReg_regD(JumpReg_regD), .MemRead_regD(
        MemRead_regD), .Rt_regD({Rt_regD[4:1], n74}), .Rs({n180, n179, n178, 
        n177, n176}), .Rt({n175, n174, n173, n172, n171}), .ICACHE_stall(
        ICACHE_stall), .DCACHE_stall(DCACHE_stall), .stall_lw_use(stall_lw_use), .stallcache(stallcache), .flush(flush), .pred_cond(pred_cond) );
  branch_prediction i_branch_prediction ( .clk(clk), .rst_n(n186), .branch(
        Branch_regD), .equal(n241) );
  precontrolDec i_precontrolDec ( .instruction_next({ICACHE_rdata[31:30], n144, 
        n126, ICACHE_rdata[27:10], n35, ICACHE_rdata[8:6], n48, 
        ICACHE_rdata[4:0]}), .Jump_IF(Jump_IF), .Branch_IF(Branch_IF) );
  nextPCcalculator i_nextPCcalculator ( .PCcur({ICACHE_addr[29:17], n58, 
        ICACHE_addr[15:4], n242, n39, ICACHE_addr[1:0], PCcur}), .PCplus4(
        PCplus4), .PCplus4_regD(PCplus4_regD), .targetAddr({ICACHE_rdata[25:6], 
        n48, ICACHE_rdata[4:0]}), .branchOffset_I({ICACHE_rdata[15:6], n48, 
        ICACHE_rdata[4:0]}), .branchOffset_regD(branchOffset_regD), 
        .JumpRegAddr({n69, n93, n113, n145, n83, n50, n98, n87, n92, n97, n95, 
        n123, n90, n67, n115, n86, n65, n63, n56, n99, n109, n84, n104, n117, 
        n111, n64, n100, n54, n120, n89, n128, n96}), .PCsrc(PCsrc), .PCnext(
        PCnext) );
  PCsrcLogic i_PCsrcLogic ( .pred_cond(pred_cond), .Branch_EX(Branch_regD), 
        .Branch_IF(Branch_IF), .equal(n241), .Jump(Jump_IF), .JumpReg(
        JumpReg_regD), .predict(1'b0), .stallcache(n181), .stall_lw_use(
        stall_lw_use), .PCsrc(PCsrc) );
  ALU i_ALU ( .ALUOp_regD(ALUOp_regD), .funct_regD(funct_regD), .ALUinA({
        ALUinA[31], n93, n113, n145, ALUinA[27], n50, n98, n146, n92, n97, n95, 
        n123, n90, n67, n115, n86, n65, n63, n56, n99, n109, n84, n104, n117, 
        n111, n64, n100, n45, n120, ALUinA[2], n128, n96}), .ALUinB(ALUinB), 
        .ALUout(ALUout) );
  MIPS_Pipeline_DW01_add_1 add_403 ( .A({ICACHE_addr[29:17], n58, 
        ICACHE_addr[15:4], n242, n39, ICACHE_addr[1:0], PCcur}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(PCplus4)
         );
  DFFRX4 \PCreg_reg[2]  ( .D(PCnext[2]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[0]) );
  DFFRX2 \PCreg_reg[18]  ( .D(PCnext[18]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[16]), .QN(n57) );
  DFFRX4 \PCreg_reg[6]  ( .D(PCnext[6]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[4]) );
  DFFRX2 \PCreg_reg[26]  ( .D(PCnext[26]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[24]) );
  DFFRX4 \PCreg_reg[27]  ( .D(PCnext[27]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[25]) );
  DFFRX4 \PCreg_reg[28]  ( .D(PCnext[28]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[26]) );
  DFFRX4 \PCreg_reg[29]  ( .D(PCnext[29]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[27]) );
  DFFRX4 \PCreg_reg[23]  ( .D(PCnext[23]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[21]) );
  DFFRX4 \PCreg_reg[9]  ( .D(PCnext[9]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[7]) );
  DFFRX4 \PCreg_reg[19]  ( .D(PCnext[19]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[17]) );
  DFFRX4 \PCreg_reg[30]  ( .D(PCnext[30]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[28]) );
  DFFRX4 \PCreg_reg[7]  ( .D(PCnext[7]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[5]) );
  DFFRX2 \PCreg_reg[11]  ( .D(PCnext[11]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[9]) );
  DFFRX2 \PCreg_reg[12]  ( .D(PCnext[12]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[10]) );
  DFFRX4 \PCreg_reg[25]  ( .D(PCnext[25]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[23]) );
  DFFRX4 \PCreg_reg[21]  ( .D(PCnext[21]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[19]) );
  DFFRHQX2 \PCreg_reg[15]  ( .D(PCnext[15]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[13]) );
  DFFRHQX2 \PCreg_reg[14]  ( .D(PCnext[14]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[12]) );
  DFFRX4 \PCreg_reg[22]  ( .D(PCnext[22]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[20]) );
  DFFRX4 \PCreg_reg[20]  ( .D(PCnext[20]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[18]) );
  DFFRX4 \PCreg_reg[24]  ( .D(PCnext[24]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[22]) );
  DFFRX4 \PCreg_reg[8]  ( .D(PCnext[8]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[6]) );
  DFFRX4 \PCreg_reg[31]  ( .D(PCnext[31]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[29]) );
  DFFRX4 \PCreg_reg[16]  ( .D(PCnext[16]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[14]) );
  DFFRX2 \PCreg_reg[13]  ( .D(PCnext[13]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[11]) );
  DFFRHQX2 \PCreg_reg[17]  ( .D(PCnext[17]), .CK(clk), .RN(rst_n), .Q(
        ICACHE_addr[15]) );
  DFFRX4 \PCreg_reg[0]  ( .D(PCnext[0]), .CK(clk), .RN(n186), .Q(PCcur[0]) );
  DFFRX4 \PCreg_reg[1]  ( .D(PCnext[1]), .CK(clk), .RN(n186), .Q(PCcur[1]) );
  DFFRX4 \PCreg_reg[10]  ( .D(PCnext[10]), .CK(clk), .RN(n186), .Q(
        ICACHE_addr[8]) );
  NOR2X6 U37 ( .A(n201), .B(n202), .Y(n209) );
  NOR2X6 U38 ( .A(n213), .B(n214), .Y(n224) );
  BUFX3 U39 ( .A(ICACHE_rdata[9]), .Y(n35) );
  CLKBUFX2 U40 ( .A(ALUinA[23]), .Y(n36) );
  INVXL U41 ( .A(ALUinA[22]), .Y(n37) );
  INVX3 U42 ( .A(n37), .Y(n38) );
  NAND4X8 U43 ( .A(n207), .B(n209), .C(n210), .D(n208), .Y(n211) );
  BUFX12 U44 ( .A(ICACHE_rdata[29]), .Y(n144) );
  BUFX20 U45 ( .A(ALUinA[12]), .Y(n99) );
  NAND4X8 U46 ( .A(n197), .B(n195), .C(n196), .D(n198), .Y(n212) );
  BUFX20 U47 ( .A(ALUinA[28]), .Y(n145) );
  INVX6 U48 ( .A(n85), .Y(n86) );
  CLKBUFX20 U49 ( .A(stallcache), .Y(n181) );
  CLKAND2X2 U50 ( .A(n238), .B(n108), .Y(n241) );
  CLKBUFX12 U51 ( .A(ALUinA[19]), .Y(n90) );
  XNOR2X4 U52 ( .A(tempALUinB[3]), .B(n119), .Y(n227) );
  INVX16 U53 ( .A(n119), .Y(n120) );
  NOR2X8 U54 ( .A(n228), .B(n227), .Y(n234) );
  NOR2X6 U55 ( .A(n191), .B(n192), .Y(n196) );
  NOR2X6 U56 ( .A(n190), .B(n189), .Y(n197) );
  NOR2X6 U57 ( .A(n199), .B(n200), .Y(n210) );
  BUFX8 U58 ( .A(wsel_regM[1]), .Y(n94) );
  NOR2X6 U59 ( .A(n187), .B(n188), .Y(n198) );
  NOR2X6 U60 ( .A(n194), .B(n193), .Y(n195) );
  AND2X8 U61 ( .A(n238), .B(n108), .Y(n40) );
  CLKBUFX4 U62 ( .A(ALUinA[30]), .Y(n93) );
  BUFX8 U63 ( .A(ICACHE_rdata[28]), .Y(n126) );
  MX2X6 U64 ( .A(ExtOut_regD[10]), .B(tempALUinB[10]), .S0(n169), .Y(
        ALUinB[10]) );
  BUFX20 U65 ( .A(n256), .Y(DCACHE_addr[14]) );
  NOR2X6 U66 ( .A(n219), .B(n220), .Y(n221) );
  NOR2X6 U67 ( .A(n216), .B(n215), .Y(n223) );
  INVX3 U68 ( .A(wsel_regM[4]), .Y(n46) );
  INVX12 U69 ( .A(n112), .Y(n113) );
  CLKINVX6 U70 ( .A(ALUinA[6]), .Y(n105) );
  BUFX12 U71 ( .A(tempALUinB[6]), .Y(n62) );
  INVX6 U72 ( .A(n60), .Y(ICACHE_addr[2]) );
  MX2X2 U73 ( .A(ExtOut_regD[0]), .B(tempALUinB[0]), .S0(n169), .Y(ALUinB[0])
         );
  MX2X2 U74 ( .A(ExtOut_regD[5]), .B(tempALUinB[5]), .S0(n169), .Y(ALUinB[5])
         );
  AND2X2 U75 ( .A(n240), .B(n239), .Y(n41) );
  CLKMX2X4 U76 ( .A(ExtOut_regD[4]), .B(tempALUinB[4]), .S0(n169), .Y(
        ALUinB[4]) );
  BUFX20 U77 ( .A(n261), .Y(DCACHE_addr[7]) );
  BUFX20 U78 ( .A(n244), .Y(DCACHE_addr[28]) );
  BUFX20 U79 ( .A(n260), .Y(DCACHE_addr[9]) );
  BUFX20 U80 ( .A(n246), .Y(DCACHE_addr[25]) );
  AO22X2 U81 ( .A0(B[30]), .A1(n150), .B0(PCplus4_regI[30]), .B1(n162), .Y(
        B_f[30]) );
  MX2X8 U82 ( .A(ExtOut_regD[27]), .B(tempALUinB[27]), .S0(n169), .Y(
        ALUinB[27]) );
  MX2X8 U83 ( .A(ExtOut_regD[26]), .B(tempALUinB[26]), .S0(n169), .Y(
        ALUinB[26]) );
  CLKMX2X6 U84 ( .A(ExtOut_regD[3]), .B(tempALUinB[3]), .S0(n169), .Y(
        ALUinB[3]) );
  CLKBUFX2 U85 ( .A(WriteData[3]), .Y(n42) );
  XOR2X4 U86 ( .A(tempALUinB[5]), .B(ALUinA[5]), .Y(n43) );
  BUFX12 U87 ( .A(n38), .Y(n97) );
  CLKINVX3 U88 ( .A(ALUinA[9]), .Y(n103) );
  INVX4 U89 ( .A(ALUinA[8]), .Y(n116) );
  BUFX16 U90 ( .A(ALUinA[0]), .Y(n96) );
  INVX1 U91 ( .A(ALUinA[4]), .Y(n44) );
  INVX6 U92 ( .A(n44), .Y(n45) );
  INVX6 U93 ( .A(n46), .Y(n47) );
  CLKINVX4 U94 ( .A(ALUinA[1]), .Y(n127) );
  CLKINVX4 U95 ( .A(ALUinA[20]), .Y(n122) );
  CLKINVX12 U96 ( .A(n114), .Y(n115) );
  NAND4X8 U97 ( .A(n223), .B(n222), .C(n221), .D(n224), .Y(n237) );
  BUFX6 U98 ( .A(ICACHE_rdata[5]), .Y(n48) );
  CLKINVX2 U99 ( .A(ALUinA[26]), .Y(n49) );
  INVX8 U100 ( .A(n49), .Y(n50) );
  BUFX3 U101 ( .A(tempALUinB[12]), .Y(n51) );
  NOR2X6 U102 ( .A(n203), .B(n204), .Y(n208) );
  CLKMX2X8 U103 ( .A(ExtOut_regD[29]), .B(tempALUinB[29]), .S0(n169), .Y(
        ALUinB[29]) );
  CLKINVX4 U104 ( .A(ALUinA[29]), .Y(n112) );
  CLKBUFX2 U105 ( .A(tempALUinB[29]), .Y(n53) );
  CLKBUFX2 U106 ( .A(n45), .Y(n54) );
  CLKBUFX8 U107 ( .A(rst_n), .Y(n186) );
  CLKBUFX20 U108 ( .A(rst_n), .Y(ICACHE_ren) );
  XOR2X4 U109 ( .A(tempALUinB[0]), .B(ALUinA[0]), .Y(n220) );
  XOR2X4 U110 ( .A(tempALUinB[11]), .B(ALUinA[11]), .Y(n202) );
  XOR2X4 U111 ( .A(tempALUinB[20]), .B(ALUinA[20]), .Y(n191) );
  NOR2X6 U112 ( .A(n218), .B(n217), .Y(n222) );
  CLKINVX2 U113 ( .A(ALUinA[13]), .Y(n55) );
  INVX12 U114 ( .A(n55), .Y(n56) );
  INVX4 U115 ( .A(n57), .Y(n58) );
  BUFX8 U116 ( .A(wsel_regM[3]), .Y(n59) );
  XOR2X4 U117 ( .A(tempALUinB[23]), .B(ALUinA[23]), .Y(n194) );
  CLKMX2X12 U118 ( .A(ExtOut_regD[23]), .B(tempALUinB[23]), .S0(n170), .Y(
        ALUinB[23]) );
  BUFX20 U119 ( .A(ALUinA[14]), .Y(n63) );
  XOR2X4 U120 ( .A(tempALUinB[21]), .B(n95), .Y(n192) );
  MX2X8 U121 ( .A(ExtOut_regD[21]), .B(tempALUinB[21]), .S0(n170), .Y(
        ALUinB[21]) );
  CLKMX2X12 U122 ( .A(ExtOut_regD[30]), .B(tempALUinB[30]), .S0(n169), .Y(
        ALUinB[30]) );
  XOR2X4 U123 ( .A(tempALUinB[10]), .B(ALUinA[10]), .Y(n201) );
  XOR2X4 U124 ( .A(tempALUinB[9]), .B(ALUinA[9]), .Y(n200) );
  INVX8 U125 ( .A(n105), .Y(n64) );
  XOR2X4 U126 ( .A(tempALUinB[8]), .B(ALUinA[8]), .Y(n199) );
  XOR2X4 U127 ( .A(tempALUinB[29]), .B(ALUinA[29]), .Y(n217) );
  XOR2X4 U128 ( .A(tempALUinB[17]), .B(ALUinA[17]), .Y(n188) );
  INVX6 U129 ( .A(ALUinA[17]), .Y(n114) );
  BUFX20 U130 ( .A(ALUinA[15]), .Y(n65) );
  NAND4X8 U131 ( .A(n234), .B(n235), .C(n233), .D(n232), .Y(n236) );
  CLKINVX2 U132 ( .A(ALUinA[18]), .Y(n66) );
  INVX8 U133 ( .A(n66), .Y(n67) );
  XOR2X4 U134 ( .A(tempALUinB[14]), .B(ALUinA[14]), .Y(n205) );
  XOR2X4 U135 ( .A(tempALUinB[1]), .B(ALUinA[1]), .Y(n225) );
  INVX6 U136 ( .A(n122), .Y(n123) );
  INVXL U137 ( .A(ALUinA[31]), .Y(n68) );
  INVX1 U138 ( .A(n68), .Y(n69) );
  NOR2X8 U139 ( .A(n229), .B(n43), .Y(n233) );
  INVXL U140 ( .A(ICACHE_rdata[27]), .Y(n70) );
  CLKINVX2 U141 ( .A(n70), .Y(n71) );
  BUFX4 U142 ( .A(flush), .Y(n72) );
  INVXL U143 ( .A(Rt_regD[0]), .Y(n73) );
  INVX3 U144 ( .A(n73), .Y(n74) );
  INVX8 U145 ( .A(n101), .Y(ICACHE_addr[3]) );
  MX2X2 U146 ( .A(ExtOut_regD[2]), .B(tempALUinB[2]), .S0(n169), .Y(ALUinB[2])
         );
  XOR2X4 U147 ( .A(tempALUinB[30]), .B(ALUinA[30]), .Y(n218) );
  INVXL U148 ( .A(ICACHE_rdata[30]), .Y(n75) );
  INVX1 U149 ( .A(n75), .Y(n76) );
  INVXL U150 ( .A(ICACHE_rdata[31]), .Y(n77) );
  INVX2 U151 ( .A(n77), .Y(n78) );
  INVX16 U152 ( .A(n116), .Y(n117) );
  CLKBUFX2 U153 ( .A(wsel_regM[0]), .Y(n82) );
  CLKBUFX2 U154 ( .A(ALUinA[27]), .Y(n83) );
  BUFX20 U155 ( .A(ALUinA[10]), .Y(n84) );
  INVX1 U156 ( .A(ALUinA[16]), .Y(n85) );
  CLKBUFX2 U157 ( .A(n146), .Y(n87) );
  CLKBUFX2 U158 ( .A(wsel_regM[2]), .Y(n88) );
  NAND2X8 U159 ( .A(n106), .B(n107), .Y(n229) );
  CLKBUFX2 U160 ( .A(ALUinA[2]), .Y(n89) );
  MX2X2 U161 ( .A(ExtOut_regD[1]), .B(tempALUinB[1]), .S0(n169), .Y(ALUinB[1])
         );
  CLKMX2X12 U162 ( .A(ExtOut_regD[8]), .B(tempALUinB[8]), .S0(n169), .Y(
        ALUinB[8]) );
  INVX16 U163 ( .A(n127), .Y(n128) );
  MX2X8 U164 ( .A(ExtOut_regD[9]), .B(tempALUinB[9]), .S0(n169), .Y(ALUinB[9])
         );
  XOR2X4 U165 ( .A(tempALUinB[22]), .B(ALUinA[22]), .Y(n193) );
  XOR2X4 U166 ( .A(tempALUinB[27]), .B(ALUinA[27]), .Y(n215) );
  XOR2X4 U167 ( .A(tempALUinB[26]), .B(ALUinA[26]), .Y(n214) );
  XOR2X4 U168 ( .A(ALUinA[12]), .B(tempALUinB[12]), .Y(n203) );
  CLKINVX8 U169 ( .A(n36), .Y(n91) );
  INVX16 U170 ( .A(n91), .Y(n92) );
  XOR2X4 U171 ( .A(tempALUinB[25]), .B(ALUinA[25]), .Y(n213) );
  XOR2X4 U172 ( .A(ALUinA[31]), .B(tempALUinB[31]), .Y(n219) );
  BUFX20 U173 ( .A(ALUinA[21]), .Y(n95) );
  XOR2X4 U174 ( .A(tempALUinB[13]), .B(ALUinA[13]), .Y(n204) );
  NAND2BX4 U175 ( .AN(tempALUinB[6]), .B(ALUinA[6]), .Y(n107) );
  BUFX20 U176 ( .A(n264), .Y(DCACHE_addr[4]) );
  BUFX20 U177 ( .A(ALUinA[25]), .Y(n98) );
  MX2X8 U178 ( .A(ExtOut_regD[22]), .B(tempALUinB[22]), .S0(n170), .Y(
        ALUinB[22]) );
  MX2X8 U179 ( .A(ExtOut_regD[19]), .B(tempALUinB[19]), .S0(n170), .Y(
        ALUinB[19]) );
  XOR2X4 U180 ( .A(tempALUinB[4]), .B(ALUinA[4]), .Y(n228) );
  BUFX20 U181 ( .A(ALUinA[5]), .Y(n100) );
  XOR2X4 U182 ( .A(tempALUinB[19]), .B(ALUinA[19]), .Y(n190) );
  MX2X8 U183 ( .A(ExtOut_regD[12]), .B(n51), .S0(n169), .Y(ALUinB[12]) );
  MX2X8 U184 ( .A(ExtOut_regD[11]), .B(tempALUinB[11]), .S0(n169), .Y(
        ALUinB[11]) );
  NOR2X8 U185 ( .A(n236), .B(n237), .Y(n108) );
  INVX16 U186 ( .A(n103), .Y(n104) );
  MX2X8 U187 ( .A(ExtOut_regD[24]), .B(tempALUinB[24]), .S0(n170), .Y(
        ALUinB[24]) );
  MX2X8 U188 ( .A(ExtOut_regD[7]), .B(tempALUinB[7]), .S0(n169), .Y(ALUinB[7])
         );
  NAND2X6 U189 ( .A(n62), .B(n105), .Y(n106) );
  MX2X8 U190 ( .A(ExtOut_regD[14]), .B(tempALUinB[14]), .S0(n170), .Y(
        ALUinB[14]) );
  MX2X8 U191 ( .A(ExtOut_regD[15]), .B(tempALUinB[15]), .S0(n170), .Y(
        ALUinB[15]) );
  BUFX20 U192 ( .A(ALUinA[11]), .Y(n109) );
  MX2X8 U193 ( .A(ExtOut_regD[17]), .B(tempALUinB[17]), .S0(n170), .Y(
        ALUinB[17]) );
  MX2X8 U194 ( .A(ExtOut_regD[13]), .B(tempALUinB[13]), .S0(n170), .Y(
        ALUinB[13]) );
  NOR2X8 U195 ( .A(n211), .B(n212), .Y(n238) );
  MX2X8 U196 ( .A(ExtOut_regD[20]), .B(tempALUinB[20]), .S0(n170), .Y(
        ALUinB[20]) );
  MX2X8 U197 ( .A(ExtOut_regD[6]), .B(n62), .S0(n169), .Y(ALUinB[6]) );
  MX2X8 U198 ( .A(ExtOut_regD[28]), .B(tempALUinB[28]), .S0(n169), .Y(
        ALUinB[28]) );
  XOR2X4 U199 ( .A(tempALUinB[15]), .B(ALUinA[15]), .Y(n206) );
  MX2X8 U200 ( .A(ExtOut_regD[16]), .B(tempALUinB[16]), .S0(n170), .Y(
        ALUinB[16]) );
  NOR2X8 U201 ( .A(n205), .B(n206), .Y(n207) );
  MX2X8 U202 ( .A(ExtOut_regD[18]), .B(tempALUinB[18]), .S0(n170), .Y(
        ALUinB[18]) );
  BUFX20 U203 ( .A(n265), .Y(DCACHE_addr[3]) );
  BUFX20 U204 ( .A(ALUinA[24]), .Y(n146) );
  NOR2X6 U205 ( .A(n230), .B(n231), .Y(n232) );
  BUFX20 U206 ( .A(n266), .Y(DCACHE_addr[2]) );
  CLKBUFX20 U207 ( .A(n255), .Y(DCACHE_addr[15]) );
  CLKINVX1 U208 ( .A(n149), .Y(n166) );
  INVX8 U209 ( .A(n157), .Y(n154) );
  INVX8 U210 ( .A(n158), .Y(n153) );
  INVX8 U211 ( .A(n158), .Y(n152) );
  AND2X2 U212 ( .A(A[2]), .B(n153), .Y(A_f[2]) );
  AND2X2 U213 ( .A(A[3]), .B(n153), .Y(A_f[3]) );
  AND2X2 U214 ( .A(A[4]), .B(n153), .Y(A_f[4]) );
  AND2X2 U215 ( .A(A[18]), .B(n154), .Y(A_f[18]) );
  AND2X2 U216 ( .A(A[19]), .B(n154), .Y(A_f[19]) );
  AND2X2 U217 ( .A(A[24]), .B(n153), .Y(A_f[24]) );
  AND2X2 U218 ( .A(A[25]), .B(n153), .Y(A_f[25]) );
  AND2X2 U219 ( .A(A[26]), .B(n153), .Y(A_f[26]) );
  AND2X2 U220 ( .A(A[27]), .B(n153), .Y(A_f[27]) );
  AND2X2 U221 ( .A(A[28]), .B(n153), .Y(A_f[28]) );
  AND2X2 U222 ( .A(A[29]), .B(n153), .Y(A_f[29]) );
  AND2X2 U223 ( .A(A[30]), .B(n153), .Y(A_f[30]) );
  AND2X2 U224 ( .A(A[31]), .B(n153), .Y(A_f[31]) );
  BUFX12 U225 ( .A(Rt[1]), .Y(n172) );
  BUFX8 U226 ( .A(Rt[0]), .Y(n171) );
  BUFX8 U227 ( .A(Rs[0]), .Y(n176) );
  INVX6 U228 ( .A(n159), .Y(n151) );
  INVX1 U229 ( .A(n156), .Y(n155) );
  INVX1 U230 ( .A(n149), .Y(n164) );
  INVX1 U231 ( .A(n149), .Y(n167) );
  BUFX20 U232 ( .A(n168), .Y(n169) );
  AND2XL U233 ( .A(A[5]), .B(n152), .Y(A_f[5]) );
  AND2XL U234 ( .A(A[6]), .B(n152), .Y(A_f[6]) );
  AND2XL U235 ( .A(A[7]), .B(n152), .Y(A_f[7]) );
  AND2XL U236 ( .A(A[8]), .B(n152), .Y(A_f[8]) );
  AND2XL U237 ( .A(A[9]), .B(n152), .Y(A_f[9]) );
  AND2XL U238 ( .A(MemWrite), .B(n41), .Y(MemWrite_m) );
  AND2XL U239 ( .A(A[1]), .B(n154), .Y(A_f[1]) );
  AND2XL U240 ( .A(A[14]), .B(n154), .Y(A_f[14]) );
  CLKBUFX20 U241 ( .A(n251), .Y(DCACHE_addr[19]) );
  BUFX6 U242 ( .A(Rt[3]), .Y(n174) );
  BUFX6 U243 ( .A(Rt[2]), .Y(n173) );
  BUFX6 U244 ( .A(Rs[3]), .Y(n179) );
  BUFX6 U245 ( .A(Rs[2]), .Y(n178) );
  BUFX8 U246 ( .A(Rs[4]), .Y(n180) );
  INVX3 U247 ( .A(n165), .Y(n150) );
  CLKBUFX3 U248 ( .A(n166), .Y(n158) );
  CLKBUFX3 U249 ( .A(n166), .Y(n159) );
  CLKBUFX3 U250 ( .A(n167), .Y(n157) );
  CLKBUFX3 U251 ( .A(n167), .Y(n156) );
  CLKBUFX3 U252 ( .A(n165), .Y(n160) );
  CLKBUFX3 U253 ( .A(n165), .Y(n161) );
  CLKBUFX3 U254 ( .A(n164), .Y(n162) );
  CLKBUFX3 U255 ( .A(n164), .Y(n163) );
  CLKINVX1 U256 ( .A(n149), .Y(n165) );
  XOR2X4 U257 ( .A(tempALUinB[28]), .B(n145), .Y(n216) );
  CLKINVX1 U258 ( .A(stall_lw_use), .Y(n239) );
  INVXL U259 ( .A(n72), .Y(n240) );
  XOR2X4 U260 ( .A(tempALUinB[24]), .B(n146), .Y(n231) );
  CLKBUFX3 U261 ( .A(n168), .Y(n170) );
  BUFX4 U262 ( .A(n52), .Y(n149) );
  NAND2BX1 U263 ( .AN(MemtoReg[0]), .B(MemtoReg[1]), .Y(n52) );
  AND2XL U264 ( .A(MemRead), .B(n41), .Y(MemRead_m) );
  AND2XL U265 ( .A(Branch_DEC), .B(n41), .Y(Branch_DEC_m) );
  AND2XL U266 ( .A(JumpReg), .B(n41), .Y(JumpReg_m) );
  AO22X1 U267 ( .A0(B[0]), .A1(n152), .B0(PCplus4_regI[0]), .B1(n156), .Y(
        B_f[0]) );
  AO22X1 U268 ( .A0(B[1]), .A1(n151), .B0(PCplus4_regI[1]), .B1(n160), .Y(
        B_f[1]) );
  AO22X1 U269 ( .A0(B[2]), .A1(n150), .B0(PCplus4_regI[2]), .B1(n162), .Y(
        B_f[2]) );
  AO22X1 U270 ( .A0(B[3]), .A1(n150), .B0(PCplus4_regI[3]), .B1(n163), .Y(
        B_f[3]) );
  AO22X1 U271 ( .A0(B[4]), .A1(n150), .B0(PCplus4_regI[4]), .B1(n163), .Y(
        B_f[4]) );
  AO22X1 U272 ( .A0(B[5]), .A1(n150), .B0(PCplus4_regI[5]), .B1(n163), .Y(
        B_f[5]) );
  AO22X1 U273 ( .A0(B[6]), .A1(n150), .B0(PCplus4_regI[6]), .B1(n163), .Y(
        B_f[6]) );
  AO22X1 U274 ( .A0(B[7]), .A1(n150), .B0(PCplus4_regI[7]), .B1(n163), .Y(
        B_f[7]) );
  AO22X1 U275 ( .A0(B[8]), .A1(n150), .B0(PCplus4_regI[8]), .B1(n156), .Y(
        B_f[8]) );
  AO22X1 U276 ( .A0(B[9]), .A1(n150), .B0(PCplus4_regI[9]), .B1(n156), .Y(
        B_f[9]) );
  AO22X1 U277 ( .A0(B[10]), .A1(n152), .B0(PCplus4_regI[10]), .B1(n157), .Y(
        B_f[10]) );
  AO22X1 U278 ( .A0(B[11]), .A1(n152), .B0(PCplus4_regI[11]), .B1(n158), .Y(
        B_f[11]) );
  AO22X1 U279 ( .A0(B[12]), .A1(n152), .B0(PCplus4_regI[12]), .B1(n156), .Y(
        B_f[12]) );
  AO22X1 U280 ( .A0(B[13]), .A1(n152), .B0(PCplus4_regI[13]), .B1(n159), .Y(
        B_f[13]) );
  AO22X1 U281 ( .A0(B[14]), .A1(n152), .B0(PCplus4_regI[14]), .B1(n156), .Y(
        B_f[14]) );
  AO22X1 U282 ( .A0(B[15]), .A1(n152), .B0(PCplus4_regI[15]), .B1(n160), .Y(
        B_f[15]) );
  AO22X1 U283 ( .A0(B[16]), .A1(n152), .B0(PCplus4_regI[16]), .B1(n160), .Y(
        B_f[16]) );
  AO22X1 U284 ( .A0(B[17]), .A1(n151), .B0(PCplus4_regI[17]), .B1(n160), .Y(
        B_f[17]) );
  AO22X1 U285 ( .A0(B[18]), .A1(n151), .B0(PCplus4_regI[18]), .B1(n160), .Y(
        B_f[18]) );
  AO22X1 U286 ( .A0(B[19]), .A1(n151), .B0(PCplus4_regI[19]), .B1(n160), .Y(
        B_f[19]) );
  AO22X1 U287 ( .A0(B[20]), .A1(n151), .B0(PCplus4_regI[20]), .B1(n161), .Y(
        B_f[20]) );
  AO22X1 U288 ( .A0(B[21]), .A1(n151), .B0(PCplus4_regI[21]), .B1(n161), .Y(
        B_f[21]) );
  AO22X1 U289 ( .A0(B[22]), .A1(n151), .B0(PCplus4_regI[22]), .B1(n161), .Y(
        B_f[22]) );
  AO22X1 U290 ( .A0(B[23]), .A1(n151), .B0(PCplus4_regI[23]), .B1(n161), .Y(
        B_f[23]) );
  AO22X1 U291 ( .A0(B[24]), .A1(n151), .B0(PCplus4_regI[24]), .B1(n161), .Y(
        B_f[24]) );
  AO22X1 U292 ( .A0(B[25]), .A1(n151), .B0(PCplus4_regI[25]), .B1(n161), .Y(
        B_f[25]) );
  AO22X1 U293 ( .A0(B[26]), .A1(n151), .B0(PCplus4_regI[26]), .B1(n162), .Y(
        B_f[26]) );
  AO22X1 U294 ( .A0(B[27]), .A1(n151), .B0(PCplus4_regI[27]), .B1(n162), .Y(
        B_f[27]) );
  AO22X1 U295 ( .A0(B[28]), .A1(n150), .B0(PCplus4_regI[28]), .B1(n162), .Y(
        B_f[28]) );
  AO22X1 U296 ( .A0(B[29]), .A1(n150), .B0(PCplus4_regI[29]), .B1(n162), .Y(
        B_f[29]) );
  AO22X1 U297 ( .A0(B[31]), .A1(n150), .B0(PCplus4_regI[31]), .B1(n163), .Y(
        B_f[31]) );
  AND2X2 U298 ( .A(A[0]), .B(n155), .Y(A_f[0]) );
  AND2X2 U299 ( .A(A[10]), .B(n154), .Y(A_f[10]) );
  AND2X2 U300 ( .A(A[11]), .B(n154), .Y(A_f[11]) );
  AND2X2 U301 ( .A(A[12]), .B(n154), .Y(A_f[12]) );
  AND2X2 U302 ( .A(A[13]), .B(n154), .Y(A_f[13]) );
  AND2X2 U303 ( .A(A[15]), .B(n154), .Y(A_f[15]) );
  AND2X2 U304 ( .A(A[16]), .B(n154), .Y(A_f[16]) );
  AND2X2 U305 ( .A(A[17]), .B(n154), .Y(A_f[17]) );
  AND2X2 U306 ( .A(A[20]), .B(n154), .Y(A_f[20]) );
  AND2X2 U307 ( .A(A[21]), .B(n154), .Y(A_f[21]) );
  AND2X2 U308 ( .A(A[22]), .B(n153), .Y(A_f[22]) );
  AND2X2 U309 ( .A(A[23]), .B(n153), .Y(A_f[23]) );
  AND2XL U310 ( .A(RegWrite), .B(n41), .Y(RegWrite_m) );
  BUFX20 U311 ( .A(n263), .Y(DCACHE_addr[5]) );
  BUFX20 U312 ( .A(n267), .Y(DCACHE_addr[1]) );
  CLKBUFX16 U313 ( .A(n249), .Y(DCACHE_addr[21]) );
  BUFX8 U314 ( .A(ALUsrc_regD), .Y(n168) );
  BUFX8 U315 ( .A(Rt[4]), .Y(n175) );
  BUFX12 U316 ( .A(Rs[1]), .Y(n177) );
  BUFX20 U317 ( .A(ALUinA[7]), .Y(n111) );
  CLKINVX8 U318 ( .A(ALUinA[3]), .Y(n119) );
  CLKBUFX20 U319 ( .A(n248), .Y(DCACHE_addr[23]) );
  CLKBUFX20 U320 ( .A(n258), .Y(DCACHE_addr[12]) );
  CLKBUFX20 U321 ( .A(n250), .Y(DCACHE_addr[20]) );
  CLKBUFX20 U322 ( .A(n254), .Y(DCACHE_addr[16]) );
  CLKBUFX20 U323 ( .A(n243), .Y(DCACHE_addr[29]) );
  CLKBUFX20 U324 ( .A(n247), .Y(DCACHE_addr[24]) );
  BUFX20 U325 ( .A(n252), .Y(DCACHE_addr[18]) );
  BUFX20 U326 ( .A(n245), .Y(DCACHE_addr[27]) );
  BUFX20 U327 ( .A(n259), .Y(DCACHE_addr[10]) );
  BUFX20 U328 ( .A(n253), .Y(DCACHE_addr[17]) );
  BUFX20 U329 ( .A(n262), .Y(DCACHE_addr[6]) );
  XOR2X4 U330 ( .A(tempALUinB[18]), .B(ALUinA[18]), .Y(n189) );
  BUFX20 U331 ( .A(n257), .Y(DCACHE_addr[13]) );
  CLKMX2X4 U332 ( .A(ExtOut_regD[25]), .B(tempALUinB[25]), .S0(n170), .Y(
        ALUinB[25]) );
  CLKMX2X4 U333 ( .A(ExtOut_regD[31]), .B(tempALUinB[31]), .S0(n169), .Y(
        ALUinB[31]) );
  XOR2X4 U334 ( .A(tempALUinB[16]), .B(ALUinA[16]), .Y(n187) );
  XOR2X4 U335 ( .A(tempALUinB[2]), .B(ALUinA[2]), .Y(n226) );
  NOR2X6 U336 ( .A(n225), .B(n226), .Y(n235) );
  XOR2X4 U337 ( .A(tempALUinB[7]), .B(n111), .Y(n230) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, \blocktag[7][24] ,
         \blocktag[7][23] , \blocktag[7][22] , \blocktag[7][21] ,
         \blocktag[7][20] , \blocktag[7][19] , \blocktag[7][18] ,
         \blocktag[7][17] , \blocktag[7][16] , \blocktag[7][15] ,
         \blocktag[7][14] , \blocktag[7][13] , \blocktag[7][12] ,
         \blocktag[7][11] , \blocktag[7][10] , \blocktag[7][9] ,
         \blocktag[7][8] , \blocktag[7][7] , \blocktag[7][6] ,
         \blocktag[7][5] , \blocktag[7][4] , \blocktag[7][3] ,
         \blocktag[7][2] , \blocktag[7][1] , \blocktag[7][0] ,
         \blocktag[6][24] , \blocktag[6][23] , \blocktag[6][22] ,
         \blocktag[6][21] , \blocktag[6][20] , \blocktag[6][19] ,
         \blocktag[6][18] , \blocktag[6][17] , \blocktag[6][16] ,
         \blocktag[6][15] , \blocktag[6][14] , \blocktag[6][13] ,
         \blocktag[6][12] , \blocktag[6][11] , \blocktag[6][10] ,
         \blocktag[6][9] , \blocktag[6][8] , \blocktag[6][7] ,
         \blocktag[6][6] , \blocktag[6][5] , \blocktag[6][4] ,
         \blocktag[6][3] , \blocktag[6][2] , \blocktag[6][1] ,
         \blocktag[6][0] , \blocktag[5][24] , \blocktag[5][23] ,
         \blocktag[5][22] , \blocktag[5][21] , \blocktag[5][20] ,
         \blocktag[5][19] , \blocktag[5][18] , \blocktag[5][17] ,
         \blocktag[5][16] , \blocktag[5][15] , \blocktag[5][14] ,
         \blocktag[5][13] , \blocktag[5][12] , \blocktag[5][11] ,
         \blocktag[5][10] , \blocktag[5][9] , \blocktag[5][8] ,
         \blocktag[5][7] , \blocktag[5][6] , \blocktag[5][5] ,
         \blocktag[5][4] , \blocktag[5][3] , \blocktag[5][2] ,
         \blocktag[5][1] , \blocktag[5][0] , \blocktag[4][24] ,
         \blocktag[4][23] , \blocktag[4][22] , \blocktag[4][21] ,
         \blocktag[4][20] , \blocktag[4][19] , \blocktag[4][18] ,
         \blocktag[4][17] , \blocktag[4][16] , \blocktag[4][15] ,
         \blocktag[4][14] , \blocktag[4][13] , \blocktag[4][12] ,
         \blocktag[4][11] , \blocktag[4][10] , \blocktag[4][9] ,
         \blocktag[4][8] , \blocktag[4][7] , \blocktag[4][6] ,
         \blocktag[4][5] , \blocktag[4][4] , \blocktag[4][3] ,
         \blocktag[4][2] , \blocktag[4][1] , \blocktag[4][0] ,
         \blocktag[3][24] , \blocktag[3][23] , \blocktag[3][22] ,
         \blocktag[3][21] , \blocktag[3][20] , \blocktag[3][19] ,
         \blocktag[3][18] , \blocktag[3][17] , \blocktag[3][16] ,
         \blocktag[3][15] , \blocktag[3][14] , \blocktag[3][13] ,
         \blocktag[3][12] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][9] , \blocktag[3][8] , \blocktag[3][7] ,
         \blocktag[3][6] , \blocktag[3][5] , \blocktag[3][4] ,
         \blocktag[3][3] , \blocktag[3][2] , \blocktag[3][1] ,
         \blocktag[3][0] , \blocktag[2][24] , \blocktag[2][23] ,
         \blocktag[2][22] , \blocktag[2][21] , \blocktag[2][20] ,
         \blocktag[2][19] , \blocktag[2][18] , \blocktag[2][17] ,
         \blocktag[2][16] , \blocktag[2][15] , \blocktag[2][14] ,
         \blocktag[2][13] , \blocktag[2][12] , \blocktag[2][11] ,
         \blocktag[2][10] , \blocktag[2][9] , \blocktag[2][8] ,
         \blocktag[2][7] , \blocktag[2][6] , \blocktag[2][5] ,
         \blocktag[2][4] , \blocktag[2][3] , \blocktag[2][2] ,
         \blocktag[2][1] , \blocktag[2][0] , \blocktag[1][24] ,
         \blocktag[1][23] , \blocktag[1][22] , \blocktag[1][21] ,
         \blocktag[1][20] , \blocktag[1][19] , \blocktag[1][18] ,
         \blocktag[1][17] , \blocktag[1][16] , \blocktag[1][15] ,
         \blocktag[1][14] , \blocktag[1][13] , \blocktag[1][12] ,
         \blocktag[1][11] , \blocktag[1][10] , \blocktag[1][9] ,
         \blocktag[1][8] , \blocktag[1][7] , \blocktag[1][6] ,
         \blocktag[1][5] , \blocktag[1][4] , \blocktag[1][3] ,
         \blocktag[1][2] , \blocktag[1][1] , \blocktag[1][0] ,
         \blocktag[0][24] , \blocktag[0][23] , \blocktag[0][22] ,
         \blocktag[0][21] , \blocktag[0][20] , \blocktag[0][19] ,
         \blocktag[0][18] , \blocktag[0][17] , \blocktag[0][16] ,
         \blocktag[0][15] , \blocktag[0][14] , \blocktag[0][13] ,
         \blocktag[0][12] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][9] , \blocktag[0][8] , \blocktag[0][7] ,
         \blocktag[0][6] , \blocktag[0][5] , \blocktag[0][4] ,
         \blocktag[0][3] , \blocktag[0][2] , \blocktag[0][1] ,
         \blocktag[0][0] , valid, dirty, \block[7][127] , \block[7][126] ,
         \block[7][125] , \block[7][124] , \block[7][123] , \block[7][122] ,
         \block[7][121] , \block[7][120] , \block[7][119] , \block[7][118] ,
         \block[7][117] , \block[7][116] , \block[7][115] , \block[7][114] ,
         \block[7][113] , \block[7][112] , \block[7][111] , \block[7][110] ,
         \block[7][109] , \block[7][108] , \block[7][107] , \block[7][106] ,
         \block[7][105] , \block[7][104] , \block[7][103] , \block[7][102] ,
         \block[7][101] , \block[7][100] , \block[7][99] , \block[7][98] ,
         \block[7][97] , \block[7][96] , \block[7][95] , \block[7][94] ,
         \block[7][93] , \block[7][92] , \block[7][91] , \block[7][90] ,
         \block[7][89] , \block[7][88] , \block[7][87] , \block[7][86] ,
         \block[7][85] , \block[7][84] , \block[7][83] , \block[7][82] ,
         \block[7][81] , \block[7][80] , \block[7][79] , \block[7][78] ,
         \block[7][77] , \block[7][76] , \block[7][75] , \block[7][74] ,
         \block[7][73] , \block[7][72] , \block[7][71] , \block[7][70] ,
         \block[7][69] , \block[7][68] , \block[7][67] , \block[7][66] ,
         \block[7][65] , \block[7][64] , \block[7][63] , \block[7][62] ,
         \block[7][61] , \block[7][60] , \block[7][59] , \block[7][58] ,
         \block[7][57] , \block[7][56] , \block[7][55] , \block[7][54] ,
         \block[7][53] , \block[7][52] , \block[7][51] , \block[7][50] ,
         \block[7][49] , \block[7][48] , \block[7][47] , \block[7][46] ,
         \block[7][45] , \block[7][44] , \block[7][43] , \block[7][42] ,
         \block[7][41] , \block[7][40] , \block[7][39] , \block[7][38] ,
         \block[7][37] , \block[7][36] , \block[7][35] , \block[7][34] ,
         \block[7][33] , \block[7][32] , \block[7][31] , \block[7][30] ,
         \block[7][29] , \block[7][28] , \block[7][27] , \block[7][26] ,
         \block[7][25] , \block[7][24] , \block[7][23] , \block[7][22] ,
         \block[7][21] , \block[7][20] , \block[7][19] , \block[7][18] ,
         \block[7][17] , \block[7][16] , \block[7][15] , \block[7][14] ,
         \block[7][13] , \block[7][12] , \block[7][11] , \block[7][10] ,
         \block[7][9] , \block[7][8] , \block[7][7] , \block[7][6] ,
         \block[7][5] , \block[7][4] , \block[7][3] , \block[7][2] ,
         \block[7][1] , \block[7][0] , \block[6][127] , \block[6][126] ,
         \block[6][125] , \block[6][124] , \block[6][123] , \block[6][122] ,
         \block[6][121] , \block[6][120] , \block[6][119] , \block[6][118] ,
         \block[6][117] , \block[6][116] , \block[6][115] , \block[6][114] ,
         \block[6][113] , \block[6][112] , \block[6][111] , \block[6][110] ,
         \block[6][109] , \block[6][108] , \block[6][107] , \block[6][106] ,
         \block[6][105] , \block[6][104] , \block[6][103] , \block[6][102] ,
         \block[6][101] , \block[6][100] , \block[6][99] , \block[6][98] ,
         \block[6][97] , \block[6][96] , \block[6][95] , \block[6][94] ,
         \block[6][93] , \block[6][92] , \block[6][91] , \block[6][90] ,
         \block[6][89] , \block[6][88] , \block[6][87] , \block[6][86] ,
         \block[6][85] , \block[6][84] , \block[6][83] , \block[6][82] ,
         \block[6][81] , \block[6][80] , \block[6][79] , \block[6][78] ,
         \block[6][77] , \block[6][76] , \block[6][75] , \block[6][74] ,
         \block[6][73] , \block[6][72] , \block[6][71] , \block[6][70] ,
         \block[6][69] , \block[6][68] , \block[6][67] , \block[6][66] ,
         \block[6][65] , \block[6][64] , \block[6][63] , \block[6][62] ,
         \block[6][61] , \block[6][60] , \block[6][59] , \block[6][58] ,
         \block[6][57] , \block[6][56] , \block[6][55] , \block[6][54] ,
         \block[6][53] , \block[6][52] , \block[6][51] , \block[6][50] ,
         \block[6][49] , \block[6][48] , \block[6][47] , \block[6][46] ,
         \block[6][45] , \block[6][44] , \block[6][43] , \block[6][42] ,
         \block[6][41] , \block[6][40] , \block[6][39] , \block[6][38] ,
         \block[6][37] , \block[6][36] , \block[6][35] , \block[6][34] ,
         \block[6][33] , \block[6][32] , \block[6][31] , \block[6][30] ,
         \block[6][29] , \block[6][28] , \block[6][27] , \block[6][26] ,
         \block[6][25] , \block[6][24] , \block[6][23] , \block[6][22] ,
         \block[6][21] , \block[6][20] , \block[6][19] , \block[6][18] ,
         \block[6][17] , \block[6][16] , \block[6][15] , \block[6][14] ,
         \block[6][13] , \block[6][12] , \block[6][11] , \block[6][10] ,
         \block[6][9] , \block[6][8] , \block[6][7] , \block[6][6] ,
         \block[6][5] , \block[6][4] , \block[6][3] , \block[6][2] ,
         \block[6][1] , \block[6][0] , \block[5][127] , \block[5][126] ,
         \block[5][125] , \block[5][124] , \block[5][123] , \block[5][122] ,
         \block[5][121] , \block[5][120] , \block[5][119] , \block[5][118] ,
         \block[5][117] , \block[5][116] , \block[5][115] , \block[5][114] ,
         \block[5][113] , \block[5][112] , \block[5][111] , \block[5][110] ,
         \block[5][109] , \block[5][108] , \block[5][107] , \block[5][106] ,
         \block[5][105] , \block[5][104] , \block[5][103] , \block[5][102] ,
         \block[5][101] , \block[5][100] , \block[5][99] , \block[5][98] ,
         \block[5][97] , \block[5][96] , \block[5][95] , \block[5][94] ,
         \block[5][93] , \block[5][92] , \block[5][91] , \block[5][90] ,
         \block[5][89] , \block[5][88] , \block[5][87] , \block[5][86] ,
         \block[5][85] , \block[5][84] , \block[5][83] , \block[5][82] ,
         \block[5][81] , \block[5][80] , \block[5][79] , \block[5][78] ,
         \block[5][77] , \block[5][76] , \block[5][75] , \block[5][74] ,
         \block[5][73] , \block[5][72] , \block[5][71] , \block[5][70] ,
         \block[5][69] , \block[5][68] , \block[5][67] , \block[5][66] ,
         \block[5][65] , \block[5][64] , \block[5][63] , \block[5][62] ,
         \block[5][61] , \block[5][60] , \block[5][59] , \block[5][58] ,
         \block[5][57] , \block[5][56] , \block[5][55] , \block[5][54] ,
         \block[5][53] , \block[5][52] , \block[5][51] , \block[5][50] ,
         \block[5][49] , \block[5][48] , \block[5][47] , \block[5][46] ,
         \block[5][45] , \block[5][44] , \block[5][43] , \block[5][42] ,
         \block[5][41] , \block[5][40] , \block[5][39] , \block[5][38] ,
         \block[5][37] , \block[5][36] , \block[5][35] , \block[5][34] ,
         \block[5][33] , \block[5][32] , \block[5][31] , \block[5][30] ,
         \block[5][29] , \block[5][28] , \block[5][27] , \block[5][26] ,
         \block[5][25] , \block[5][24] , \block[5][23] , \block[5][22] ,
         \block[5][21] , \block[5][20] , \block[5][19] , \block[5][18] ,
         \block[5][17] , \block[5][16] , \block[5][15] , \block[5][14] ,
         \block[5][13] , \block[5][12] , \block[5][11] , \block[5][10] ,
         \block[5][9] , \block[5][8] , \block[5][7] , \block[5][6] ,
         \block[5][5] , \block[5][4] , \block[5][3] , \block[5][2] ,
         \block[5][1] , \block[5][0] , \block[4][127] , \block[4][126] ,
         \block[4][125] , \block[4][124] , \block[4][123] , \block[4][122] ,
         \block[4][121] , \block[4][120] , \block[4][119] , \block[4][118] ,
         \block[4][117] , \block[4][116] , \block[4][115] , \block[4][114] ,
         \block[4][113] , \block[4][112] , \block[4][111] , \block[4][110] ,
         \block[4][109] , \block[4][108] , \block[4][107] , \block[4][106] ,
         \block[4][105] , \block[4][104] , \block[4][103] , \block[4][102] ,
         \block[4][101] , \block[4][100] , \block[4][99] , \block[4][98] ,
         \block[4][97] , \block[4][96] , \block[4][95] , \block[4][94] ,
         \block[4][93] , \block[4][92] , \block[4][91] , \block[4][90] ,
         \block[4][89] , \block[4][88] , \block[4][87] , \block[4][86] ,
         \block[4][85] , \block[4][84] , \block[4][83] , \block[4][82] ,
         \block[4][81] , \block[4][80] , \block[4][79] , \block[4][78] ,
         \block[4][77] , \block[4][76] , \block[4][75] , \block[4][74] ,
         \block[4][73] , \block[4][72] , \block[4][71] , \block[4][70] ,
         \block[4][69] , \block[4][68] , \block[4][67] , \block[4][66] ,
         \block[4][65] , \block[4][64] , \block[4][63] , \block[4][62] ,
         \block[4][61] , \block[4][60] , \block[4][59] , \block[4][58] ,
         \block[4][57] , \block[4][56] , \block[4][55] , \block[4][54] ,
         \block[4][53] , \block[4][52] , \block[4][51] , \block[4][50] ,
         \block[4][49] , \block[4][48] , \block[4][47] , \block[4][46] ,
         \block[4][45] , \block[4][44] , \block[4][43] , \block[4][42] ,
         \block[4][41] , \block[4][40] , \block[4][39] , \block[4][38] ,
         \block[4][37] , \block[4][36] , \block[4][35] , \block[4][34] ,
         \block[4][33] , \block[4][32] , \block[4][31] , \block[4][30] ,
         \block[4][29] , \block[4][28] , \block[4][27] , \block[4][26] ,
         \block[4][25] , \block[4][24] , \block[4][23] , \block[4][22] ,
         \block[4][21] , \block[4][20] , \block[4][19] , \block[4][18] ,
         \block[4][17] , \block[4][16] , \block[4][15] , \block[4][14] ,
         \block[4][13] , \block[4][12] , \block[4][11] , \block[4][10] ,
         \block[4][9] , \block[4][8] , \block[4][7] , \block[4][6] ,
         \block[4][5] , \block[4][4] , \block[4][3] , \block[4][2] ,
         \block[4][1] , \block[4][0] , \block[3][127] , \block[3][126] ,
         \block[3][125] , \block[3][124] , \block[3][123] , \block[3][122] ,
         \block[3][121] , \block[3][120] , \block[3][119] , \block[3][118] ,
         \block[3][117] , \block[3][116] , \block[3][115] , \block[3][114] ,
         \block[3][113] , \block[3][112] , \block[3][111] , \block[3][110] ,
         \block[3][109] , \block[3][108] , \block[3][107] , \block[3][106] ,
         \block[3][105] , \block[3][104] , \block[3][103] , \block[3][102] ,
         \block[3][101] , \block[3][100] , \block[3][99] , \block[3][98] ,
         \block[3][97] , \block[3][96] , \block[3][95] , \block[3][94] ,
         \block[3][93] , \block[3][92] , \block[3][91] , \block[3][90] ,
         \block[3][89] , \block[3][88] , \block[3][87] , \block[3][86] ,
         \block[3][85] , \block[3][84] , \block[3][83] , \block[3][82] ,
         \block[3][81] , \block[3][80] , \block[3][79] , \block[3][78] ,
         \block[3][77] , \block[3][76] , \block[3][75] , \block[3][74] ,
         \block[3][73] , \block[3][72] , \block[3][71] , \block[3][70] ,
         \block[3][69] , \block[3][68] , \block[3][67] , \block[3][66] ,
         \block[3][65] , \block[3][64] , \block[3][63] , \block[3][62] ,
         \block[3][61] , \block[3][60] , \block[3][59] , \block[3][58] ,
         \block[3][57] , \block[3][56] , \block[3][55] , \block[3][54] ,
         \block[3][53] , \block[3][52] , \block[3][51] , \block[3][50] ,
         \block[3][49] , \block[3][48] , \block[3][47] , \block[3][46] ,
         \block[3][45] , \block[3][44] , \block[3][43] , \block[3][42] ,
         \block[3][41] , \block[3][40] , \block[3][39] , \block[3][38] ,
         \block[3][37] , \block[3][36] , \block[3][35] , \block[3][34] ,
         \block[3][33] , \block[3][32] , \block[3][31] , \block[3][30] ,
         \block[3][29] , \block[3][28] , \block[3][27] , \block[3][26] ,
         \block[3][25] , \block[3][24] , \block[3][23] , \block[3][22] ,
         \block[3][21] , \block[3][20] , \block[3][19] , \block[3][18] ,
         \block[3][17] , \block[3][16] , \block[3][15] , \block[3][14] ,
         \block[3][13] , \block[3][12] , \block[3][11] , \block[3][10] ,
         \block[3][9] , \block[3][8] , \block[3][7] , \block[3][6] ,
         \block[3][5] , \block[3][4] , \block[3][3] , \block[3][2] ,
         \block[3][1] , \block[3][0] , \block[2][127] , \block[2][126] ,
         \block[2][125] , \block[2][124] , \block[2][123] , \block[2][122] ,
         \block[2][121] , \block[2][120] , \block[2][119] , \block[2][118] ,
         \block[2][117] , \block[2][116] , \block[2][115] , \block[2][114] ,
         \block[2][113] , \block[2][112] , \block[2][111] , \block[2][110] ,
         \block[2][109] , \block[2][108] , \block[2][107] , \block[2][106] ,
         \block[2][105] , \block[2][104] , \block[2][103] , \block[2][102] ,
         \block[2][101] , \block[2][100] , \block[2][99] , \block[2][98] ,
         \block[2][97] , \block[2][96] , \block[2][95] , \block[2][94] ,
         \block[2][93] , \block[2][92] , \block[2][91] , \block[2][90] ,
         \block[2][89] , \block[2][88] , \block[2][87] , \block[2][86] ,
         \block[2][85] , \block[2][84] , \block[2][83] , \block[2][82] ,
         \block[2][81] , \block[2][80] , \block[2][79] , \block[2][78] ,
         \block[2][77] , \block[2][76] , \block[2][75] , \block[2][74] ,
         \block[2][73] , \block[2][72] , \block[2][71] , \block[2][70] ,
         \block[2][69] , \block[2][68] , \block[2][67] , \block[2][66] ,
         \block[2][65] , \block[2][64] , \block[2][63] , \block[2][62] ,
         \block[2][61] , \block[2][60] , \block[2][59] , \block[2][58] ,
         \block[2][57] , \block[2][56] , \block[2][55] , \block[2][54] ,
         \block[2][53] , \block[2][52] , \block[2][51] , \block[2][50] ,
         \block[2][49] , \block[2][48] , \block[2][47] , \block[2][46] ,
         \block[2][45] , \block[2][44] , \block[2][43] , \block[2][42] ,
         \block[2][41] , \block[2][40] , \block[2][39] , \block[2][38] ,
         \block[2][37] , \block[2][36] , \block[2][35] , \block[2][34] ,
         \block[2][33] , \block[2][32] , \block[2][31] , \block[2][30] ,
         \block[2][29] , \block[2][28] , \block[2][27] , \block[2][26] ,
         \block[2][25] , \block[2][24] , \block[2][23] , \block[2][22] ,
         \block[2][21] , \block[2][20] , \block[2][19] , \block[2][18] ,
         \block[2][17] , \block[2][16] , \block[2][15] , \block[2][14] ,
         \block[2][13] , \block[2][12] , \block[2][11] , \block[2][10] ,
         \block[2][9] , \block[2][8] , \block[2][7] , \block[2][6] ,
         \block[2][5] , \block[2][4] , \block[2][3] , \block[2][2] ,
         \block[2][1] , \block[2][0] , \block[1][127] , \block[1][126] ,
         \block[1][125] , \block[1][124] , \block[1][123] , \block[1][122] ,
         \block[1][121] , \block[1][120] , \block[1][119] , \block[1][118] ,
         \block[1][117] , \block[1][116] , \block[1][115] , \block[1][114] ,
         \block[1][113] , \block[1][112] , \block[1][111] , \block[1][110] ,
         \block[1][109] , \block[1][108] , \block[1][107] , \block[1][106] ,
         \block[1][105] , \block[1][104] , \block[1][103] , \block[1][102] ,
         \block[1][101] , \block[1][100] , \block[1][99] , \block[1][98] ,
         \block[1][97] , \block[1][96] , \block[1][95] , \block[1][94] ,
         \block[1][93] , \block[1][92] , \block[1][91] , \block[1][90] ,
         \block[1][89] , \block[1][88] , \block[1][87] , \block[1][86] ,
         \block[1][85] , \block[1][84] , \block[1][83] , \block[1][82] ,
         \block[1][81] , \block[1][80] , \block[1][79] , \block[1][78] ,
         \block[1][77] , \block[1][76] , \block[1][75] , \block[1][74] ,
         \block[1][73] , \block[1][72] , \block[1][71] , \block[1][70] ,
         \block[1][69] , \block[1][68] , \block[1][67] , \block[1][66] ,
         \block[1][65] , \block[1][64] , \block[1][63] , \block[1][62] ,
         \block[1][61] , \block[1][60] , \block[1][59] , \block[1][58] ,
         \block[1][57] , \block[1][56] , \block[1][55] , \block[1][54] ,
         \block[1][53] , \block[1][52] , \block[1][51] , \block[1][50] ,
         \block[1][49] , \block[1][48] , \block[1][47] , \block[1][46] ,
         \block[1][45] , \block[1][44] , \block[1][43] , \block[1][42] ,
         \block[1][41] , \block[1][40] , \block[1][39] , \block[1][38] ,
         \block[1][37] , \block[1][36] , \block[1][35] , \block[1][34] ,
         \block[1][33] , \block[1][32] , \block[1][31] , \block[1][30] ,
         \block[1][29] , \block[1][28] , \block[1][27] , \block[1][26] ,
         \block[1][25] , \block[1][24] , \block[1][23] , \block[1][22] ,
         \block[1][21] , \block[1][20] , \block[1][19] , \block[1][18] ,
         \block[1][17] , \block[1][16] , \block[1][15] , \block[1][14] ,
         \block[1][13] , \block[1][12] , \block[1][11] , \block[1][10] ,
         \block[1][9] , \block[1][8] , \block[1][7] , \block[1][6] ,
         \block[1][5] , \block[1][4] , \block[1][3] , \block[1][2] ,
         \block[1][1] , \block[1][0] , \block[0][127] , \block[0][126] ,
         \block[0][125] , \block[0][124] , \block[0][123] , \block[0][122] ,
         \block[0][121] , \block[0][120] , \block[0][119] , \block[0][118] ,
         \block[0][117] , \block[0][116] , \block[0][115] , \block[0][114] ,
         \block[0][113] , \block[0][112] , \block[0][111] , \block[0][110] ,
         \block[0][109] , \block[0][108] , \block[0][107] , \block[0][106] ,
         \block[0][105] , \block[0][104] , \block[0][103] , \block[0][102] ,
         \block[0][101] , \block[0][100] , \block[0][99] , \block[0][98] ,
         \block[0][97] , \block[0][96] , \block[0][95] , \block[0][94] ,
         \block[0][93] , \block[0][92] , \block[0][91] , \block[0][90] ,
         \block[0][89] , \block[0][88] , \block[0][87] , \block[0][86] ,
         \block[0][85] , \block[0][84] , \block[0][83] , \block[0][82] ,
         \block[0][81] , \block[0][80] , \block[0][79] , \block[0][78] ,
         \block[0][77] , \block[0][76] , \block[0][75] , \block[0][74] ,
         \block[0][73] , \block[0][72] , \block[0][71] , \block[0][70] ,
         \block[0][69] , \block[0][68] , \block[0][67] , \block[0][66] ,
         \block[0][65] , \block[0][64] , \block[0][63] , \block[0][62] ,
         \block[0][61] , \block[0][60] , \block[0][59] , \block[0][58] ,
         \block[0][57] , \block[0][56] , \block[0][55] , \block[0][54] ,
         \block[0][53] , \block[0][52] , \block[0][51] , \block[0][50] ,
         \block[0][49] , \block[0][48] , \block[0][47] , \block[0][46] ,
         \block[0][45] , \block[0][44] , \block[0][43] , \block[0][42] ,
         \block[0][41] , \block[0][40] , \block[0][39] , \block[0][38] ,
         \block[0][37] , \block[0][36] , \block[0][35] , \block[0][34] ,
         \block[0][33] , \block[0][32] , \block[0][31] , \block[0][30] ,
         \block[0][29] , \block[0][28] , \block[0][27] , \block[0][26] ,
         \block[0][25] , \block[0][24] , \block[0][23] , \block[0][22] ,
         \block[0][21] , \block[0][20] , \block[0][19] , \block[0][18] ,
         \block[0][17] , \block[0][16] , \block[0][15] , \block[0][14] ,
         \block[0][13] , \block[0][12] , \block[0][11] , \block[0][10] ,
         \block[0][9] , \block[0][8] , \block[0][7] , \block[0][6] ,
         \block[0][5] , \block[0][4] , \block[0][3] , \block[0][2] ,
         \block[0][1] , \block[0][0] , n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n503, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n20, n22, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n93, n95, n97, n99, n100, n101, n102, n103, n104, n105, n107,
         n108, n109, n110, n111, n112, n114, n116, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n502, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1624, n1625, n1626, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  DFFRX4 \blockvalid_reg[7]  ( .D(n503), .CK(clk), .RN(n1628), .Q(
        blockvalid[7]), .QN(n486) );
  DFFRX4 \blockvalid_reg[5]  ( .D(n500), .CK(clk), .RN(n1628), .Q(
        blockvalid[5]), .QN(n484) );
  DFFRX4 \blockvalid_reg[4]  ( .D(n499), .CK(clk), .RN(n1628), .Q(
        blockvalid[4]), .QN(n483) );
  DFFRX4 \blockvalid_reg[3]  ( .D(n498), .CK(clk), .RN(n1628), .Q(
        blockvalid[3]), .QN(n482) );
  DFFQXL \block_reg[7][71]  ( .D(n1047), .CK(clk), .Q(\block[7][71] ) );
  CLKMX2X2 \block_reg[7][70]/U3  ( .A(\block[7][70] ), .B(block_next[70]), 
        .S0(n1503), .Y(n1046) );
  DFFQXL \block_reg[7][70]  ( .D(n1046), .CK(clk), .Q(\block[7][70] ) );
  CLKMX2X2 \block_reg[7][69]/U3  ( .A(\block[7][69] ), .B(block_next[69]), 
        .S0(n1503), .Y(n1045) );
  DFFQXL \block_reg[7][69]  ( .D(n1045), .CK(clk), .Q(\block[7][69] ) );
  CLKMX2X2 \block_reg[7][68]/U3  ( .A(\block[7][68] ), .B(block_next[68]), 
        .S0(n1503), .Y(n1044) );
  DFFQXL \block_reg[7][68]  ( .D(n1044), .CK(clk), .Q(\block[7][68] ) );
  DFFQXL \block_reg[7][67]  ( .D(n1043), .CK(clk), .Q(\block[7][67] ) );
  CLKMX2X2 \block_reg[7][66]/U3  ( .A(\block[7][66] ), .B(block_next[66]), 
        .S0(n1503), .Y(n1042) );
  DFFQXL \block_reg[7][66]  ( .D(n1042), .CK(clk), .Q(\block[7][66] ) );
  CLKMX2X2 \block_reg[7][65]/U3  ( .A(\block[7][65] ), .B(block_next[65]), 
        .S0(n1502), .Y(n1041) );
  DFFQXL \block_reg[7][65]  ( .D(n1041), .CK(clk), .Q(\block[7][65] ) );
  CLKMX2X2 \block_reg[7][64]/U3  ( .A(\block[7][64] ), .B(block_next[64]), 
        .S0(n1502), .Y(n1040) );
  DFFQXL \block_reg[7][64]  ( .D(n1040), .CK(clk), .Q(\block[7][64] ) );
  DFFQXL \block_reg[6][71]  ( .D(n1039), .CK(clk), .Q(\block[6][71] ) );
  CLKMX2X2 \block_reg[6][70]/U3  ( .A(\block[6][70] ), .B(block_next[70]), 
        .S0(n1518), .Y(n1038) );
  DFFQXL \block_reg[6][70]  ( .D(n1038), .CK(clk), .Q(\block[6][70] ) );
  CLKMX2X2 \block_reg[6][69]/U3  ( .A(\block[6][69] ), .B(block_next[69]), 
        .S0(n1518), .Y(n1037) );
  DFFQXL \block_reg[6][69]  ( .D(n1037), .CK(clk), .Q(\block[6][69] ) );
  CLKMX2X2 \block_reg[6][68]/U3  ( .A(\block[6][68] ), .B(block_next[68]), 
        .S0(n1518), .Y(n1036) );
  DFFQXL \block_reg[6][68]  ( .D(n1036), .CK(clk), .Q(\block[6][68] ) );
  DFFQXL \block_reg[6][67]  ( .D(n1035), .CK(clk), .Q(\block[6][67] ) );
  CLKMX2X2 \block_reg[6][66]/U3  ( .A(\block[6][66] ), .B(block_next[66]), 
        .S0(n1518), .Y(n1034) );
  DFFQXL \block_reg[6][66]  ( .D(n1034), .CK(clk), .Q(\block[6][66] ) );
  CLKMX2X2 \block_reg[6][65]/U3  ( .A(\block[6][65] ), .B(block_next[65]), 
        .S0(n1517), .Y(n1033) );
  DFFQXL \block_reg[6][65]  ( .D(n1033), .CK(clk), .Q(\block[6][65] ) );
  CLKMX2X2 \block_reg[6][64]/U3  ( .A(\block[6][64] ), .B(block_next[64]), 
        .S0(n1517), .Y(n1032) );
  DFFQXL \block_reg[6][64]  ( .D(n1032), .CK(clk), .Q(\block[6][64] ) );
  CLKMX2X2 \block_reg[5][70]/U3  ( .A(\block[5][70] ), .B(block_next[70]), 
        .S0(n1534), .Y(n1030) );
  DFFQXL \block_reg[5][70]  ( .D(n1030), .CK(clk), .Q(\block[5][70] ) );
  CLKMX2X2 \block_reg[5][69]/U3  ( .A(\block[5][69] ), .B(block_next[69]), 
        .S0(n1534), .Y(n1029) );
  DFFQXL \block_reg[5][69]  ( .D(n1029), .CK(clk), .Q(\block[5][69] ) );
  CLKMX2X2 \block_reg[5][68]/U3  ( .A(\block[5][68] ), .B(block_next[68]), 
        .S0(n1534), .Y(n1028) );
  DFFQXL \block_reg[5][68]  ( .D(n1028), .CK(clk), .Q(\block[5][68] ) );
  DFFQXL \block_reg[5][67]  ( .D(n1027), .CK(clk), .Q(\block[5][67] ) );
  CLKMX2X2 \block_reg[5][66]/U3  ( .A(\block[5][66] ), .B(block_next[66]), 
        .S0(n1534), .Y(n1026) );
  DFFQXL \block_reg[5][66]  ( .D(n1026), .CK(clk), .Q(\block[5][66] ) );
  CLKMX2X2 \block_reg[5][65]/U3  ( .A(\block[5][65] ), .B(block_next[65]), 
        .S0(n1533), .Y(n1025) );
  DFFQXL \block_reg[5][65]  ( .D(n1025), .CK(clk), .Q(\block[5][65] ) );
  CLKMX2X2 \block_reg[5][64]/U3  ( .A(\block[5][64] ), .B(block_next[64]), 
        .S0(n1533), .Y(n1024) );
  DFFQXL \block_reg[5][64]  ( .D(n1024), .CK(clk), .Q(\block[5][64] ) );
  DFFQXL \block_reg[4][71]  ( .D(n1023), .CK(clk), .Q(\block[4][71] ) );
  CLKMX2X2 \block_reg[4][70]/U3  ( .A(\block[4][70] ), .B(block_next[70]), 
        .S0(n1551), .Y(n1022) );
  DFFQXL \block_reg[4][70]  ( .D(n1022), .CK(clk), .Q(\block[4][70] ) );
  CLKMX2X2 \block_reg[4][69]/U3  ( .A(\block[4][69] ), .B(block_next[69]), 
        .S0(n1551), .Y(n1021) );
  DFFQXL \block_reg[4][69]  ( .D(n1021), .CK(clk), .Q(\block[4][69] ) );
  CLKMX2X2 \block_reg[4][68]/U3  ( .A(\block[4][68] ), .B(block_next[68]), 
        .S0(n1551), .Y(n1020) );
  DFFQXL \block_reg[4][68]  ( .D(n1020), .CK(clk), .Q(\block[4][68] ) );
  DFFQXL \block_reg[4][67]  ( .D(n1019), .CK(clk), .Q(\block[4][67] ) );
  CLKMX2X2 \block_reg[4][66]/U3  ( .A(\block[4][66] ), .B(block_next[66]), 
        .S0(n1551), .Y(n1018) );
  DFFQXL \block_reg[4][66]  ( .D(n1018), .CK(clk), .Q(\block[4][66] ) );
  CLKMX2X2 \block_reg[4][65]/U3  ( .A(\block[4][65] ), .B(block_next[65]), 
        .S0(n1550), .Y(n1017) );
  DFFQXL \block_reg[4][65]  ( .D(n1017), .CK(clk), .Q(\block[4][65] ) );
  CLKMX2X2 \block_reg[4][64]/U3  ( .A(\block[4][64] ), .B(block_next[64]), 
        .S0(n1550), .Y(n1016) );
  DFFQXL \block_reg[4][64]  ( .D(n1016), .CK(clk), .Q(\block[4][64] ) );
  DFFQXL \block_reg[3][71]  ( .D(n1015), .CK(clk), .Q(\block[3][71] ) );
  CLKMX2X2 \block_reg[3][70]/U3  ( .A(\block[3][70] ), .B(block_next[70]), 
        .S0(n1568), .Y(n1014) );
  DFFQXL \block_reg[3][70]  ( .D(n1014), .CK(clk), .Q(\block[3][70] ) );
  CLKMX2X2 \block_reg[3][69]/U3  ( .A(\block[3][69] ), .B(block_next[69]), 
        .S0(n1568), .Y(n1013) );
  DFFQXL \block_reg[3][69]  ( .D(n1013), .CK(clk), .Q(\block[3][69] ) );
  CLKMX2X2 \block_reg[3][68]/U3  ( .A(\block[3][68] ), .B(block_next[68]), 
        .S0(n1568), .Y(n1012) );
  DFFQXL \block_reg[3][68]  ( .D(n1012), .CK(clk), .Q(\block[3][68] ) );
  DFFQXL \block_reg[3][67]  ( .D(n1011), .CK(clk), .Q(\block[3][67] ) );
  CLKMX2X2 \block_reg[3][66]/U3  ( .A(\block[3][66] ), .B(block_next[66]), 
        .S0(n1568), .Y(n1010) );
  DFFQXL \block_reg[3][66]  ( .D(n1010), .CK(clk), .Q(\block[3][66] ) );
  CLKMX2X2 \block_reg[3][65]/U3  ( .A(\block[3][65] ), .B(block_next[65]), 
        .S0(n1567), .Y(n1009) );
  DFFQXL \block_reg[3][65]  ( .D(n1009), .CK(clk), .Q(\block[3][65] ) );
  CLKMX2X2 \block_reg[3][64]/U3  ( .A(\block[3][64] ), .B(block_next[64]), 
        .S0(n1567), .Y(n1008) );
  DFFQXL \block_reg[3][64]  ( .D(n1008), .CK(clk), .Q(\block[3][64] ) );
  DFFQXL \block_reg[2][71]  ( .D(n1007), .CK(clk), .Q(\block[2][71] ) );
  CLKMX2X2 \block_reg[2][70]/U3  ( .A(\block[2][70] ), .B(block_next[70]), 
        .S0(n1581), .Y(n1006) );
  DFFQXL \block_reg[2][70]  ( .D(n1006), .CK(clk), .Q(\block[2][70] ) );
  CLKMX2X2 \block_reg[2][69]/U3  ( .A(\block[2][69] ), .B(block_next[69]), 
        .S0(n1581), .Y(n1005) );
  DFFQXL \block_reg[2][69]  ( .D(n1005), .CK(clk), .Q(\block[2][69] ) );
  CLKMX2X2 \block_reg[2][68]/U3  ( .A(\block[2][68] ), .B(block_next[68]), 
        .S0(n1581), .Y(n1004) );
  DFFQXL \block_reg[2][68]  ( .D(n1004), .CK(clk), .Q(\block[2][68] ) );
  DFFQXL \block_reg[2][67]  ( .D(n1003), .CK(clk), .Q(\block[2][67] ) );
  CLKMX2X2 \block_reg[2][66]/U3  ( .A(\block[2][66] ), .B(block_next[66]), 
        .S0(n1581), .Y(n1002) );
  DFFQXL \block_reg[2][66]  ( .D(n1002), .CK(clk), .Q(\block[2][66] ) );
  CLKMX2X2 \block_reg[2][65]/U3  ( .A(\block[2][65] ), .B(block_next[65]), 
        .S0(n1580), .Y(n1001) );
  DFFQXL \block_reg[2][65]  ( .D(n1001), .CK(clk), .Q(\block[2][65] ) );
  CLKMX2X2 \block_reg[2][64]/U3  ( .A(\block[2][64] ), .B(block_next[64]), 
        .S0(n1580), .Y(n1000) );
  DFFQXL \block_reg[2][64]  ( .D(n1000), .CK(clk), .Q(\block[2][64] ) );
  DFFQXL \block_reg[1][71]  ( .D(n999), .CK(clk), .Q(\block[1][71] ) );
  CLKMX2X2 \block_reg[1][70]/U3  ( .A(\block[1][70] ), .B(block_next[70]), 
        .S0(n1595), .Y(n998) );
  DFFQXL \block_reg[1][70]  ( .D(n998), .CK(clk), .Q(\block[1][70] ) );
  CLKMX2X2 \block_reg[1][69]/U3  ( .A(\block[1][69] ), .B(block_next[69]), 
        .S0(n1595), .Y(n997) );
  DFFQXL \block_reg[1][69]  ( .D(n997), .CK(clk), .Q(\block[1][69] ) );
  CLKMX2X2 \block_reg[1][68]/U3  ( .A(\block[1][68] ), .B(block_next[68]), 
        .S0(n1595), .Y(n996) );
  DFFQXL \block_reg[1][68]  ( .D(n996), .CK(clk), .Q(\block[1][68] ) );
  DFFQXL \block_reg[1][67]  ( .D(n995), .CK(clk), .Q(\block[1][67] ) );
  CLKMX2X2 \block_reg[1][66]/U3  ( .A(\block[1][66] ), .B(block_next[66]), 
        .S0(n1595), .Y(n994) );
  DFFQXL \block_reg[1][66]  ( .D(n994), .CK(clk), .Q(\block[1][66] ) );
  CLKMX2X2 \block_reg[1][65]/U3  ( .A(\block[1][65] ), .B(block_next[65]), 
        .S0(n1594), .Y(n993) );
  DFFQXL \block_reg[1][65]  ( .D(n993), .CK(clk), .Q(\block[1][65] ) );
  CLKMX2X2 \block_reg[1][64]/U3  ( .A(\block[1][64] ), .B(block_next[64]), 
        .S0(n1594), .Y(n992) );
  DFFQXL \block_reg[1][64]  ( .D(n992), .CK(clk), .Q(\block[1][64] ) );
  DFFQXL \block_reg[0][71]  ( .D(n991), .CK(clk), .Q(\block[0][71] ) );
  CLKMX2X2 \block_reg[0][70]/U3  ( .A(\block[0][70] ), .B(block_next[70]), 
        .S0(n1610), .Y(n990) );
  DFFQXL \block_reg[0][70]  ( .D(n990), .CK(clk), .Q(\block[0][70] ) );
  CLKMX2X2 \block_reg[0][69]/U3  ( .A(\block[0][69] ), .B(block_next[69]), 
        .S0(n1610), .Y(n989) );
  DFFQXL \block_reg[0][69]  ( .D(n989), .CK(clk), .Q(\block[0][69] ) );
  CLKMX2X2 \block_reg[0][68]/U3  ( .A(\block[0][68] ), .B(block_next[68]), 
        .S0(n1610), .Y(n988) );
  DFFQXL \block_reg[0][68]  ( .D(n988), .CK(clk), .Q(\block[0][68] ) );
  CLKMX2X2 \block_reg[0][66]/U3  ( .A(\block[0][66] ), .B(block_next[66]), 
        .S0(n1610), .Y(n986) );
  DFFQXL \block_reg[0][66]  ( .D(n986), .CK(clk), .Q(\block[0][66] ) );
  CLKMX2X2 \block_reg[0][65]/U3  ( .A(\block[0][65] ), .B(block_next[65]), 
        .S0(n1609), .Y(n985) );
  DFFQXL \block_reg[0][65]  ( .D(n985), .CK(clk), .Q(\block[0][65] ) );
  CLKMX2X2 \block_reg[0][64]/U3  ( .A(\block[0][64] ), .B(block_next[64]), 
        .S0(n1609), .Y(n984) );
  DFFQXL \block_reg[0][64]  ( .D(n984), .CK(clk), .Q(\block[0][64] ) );
  CLKMX2X2 \block_reg[7][103]/U3  ( .A(\block[7][103] ), .B(block_next[103]), 
        .S0(n1505), .Y(n983) );
  DFFQXL \block_reg[7][103]  ( .D(n983), .CK(clk), .Q(\block[7][103] ) );
  CLKMX2X2 \block_reg[7][102]/U3  ( .A(\block[7][102] ), .B(block_next[102]), 
        .S0(n1505), .Y(n982) );
  DFFQXL \block_reg[7][102]  ( .D(n982), .CK(clk), .Q(\block[7][102] ) );
  CLKMX2X2 \block_reg[7][101]/U3  ( .A(\block[7][101] ), .B(block_next[101]), 
        .S0(n1505), .Y(n981) );
  DFFQXL \block_reg[7][101]  ( .D(n981), .CK(clk), .Q(\block[7][101] ) );
  CLKMX2X2 \block_reg[7][100]/U3  ( .A(\block[7][100] ), .B(block_next[100]), 
        .S0(n1505), .Y(n980) );
  DFFQXL \block_reg[7][100]  ( .D(n980), .CK(clk), .Q(\block[7][100] ) );
  DFFQXL \block_reg[7][99]  ( .D(n979), .CK(clk), .Q(\block[7][99] ) );
  CLKMX2X2 \block_reg[7][98]/U3  ( .A(\block[7][98] ), .B(block_next[98]), 
        .S0(n1505), .Y(n978) );
  DFFQXL \block_reg[7][98]  ( .D(n978), .CK(clk), .Q(\block[7][98] ) );
  CLKMX2X2 \block_reg[7][97]/U3  ( .A(\block[7][97] ), .B(block_next[97]), 
        .S0(n1505), .Y(n977) );
  DFFQXL \block_reg[7][97]  ( .D(n977), .CK(clk), .Q(\block[7][97] ) );
  CLKMX2X2 \block_reg[6][103]/U3  ( .A(\block[6][103] ), .B(block_next[103]), 
        .S0(n1520), .Y(n976) );
  DFFQXL \block_reg[6][103]  ( .D(n976), .CK(clk), .Q(\block[6][103] ) );
  CLKMX2X2 \block_reg[6][102]/U3  ( .A(\block[6][102] ), .B(block_next[102]), 
        .S0(n1520), .Y(n975) );
  DFFQXL \block_reg[6][102]  ( .D(n975), .CK(clk), .Q(\block[6][102] ) );
  CLKMX2X2 \block_reg[6][101]/U3  ( .A(\block[6][101] ), .B(block_next[101]), 
        .S0(n1520), .Y(n974) );
  DFFQXL \block_reg[6][101]  ( .D(n974), .CK(clk), .Q(\block[6][101] ) );
  CLKMX2X2 \block_reg[6][100]/U3  ( .A(\block[6][100] ), .B(block_next[100]), 
        .S0(n1520), .Y(n973) );
  DFFQXL \block_reg[6][100]  ( .D(n973), .CK(clk), .Q(\block[6][100] ) );
  DFFQXL \block_reg[6][99]  ( .D(n972), .CK(clk), .Q(\block[6][99] ) );
  CLKMX2X2 \block_reg[6][98]/U3  ( .A(\block[6][98] ), .B(block_next[98]), 
        .S0(n1520), .Y(n971) );
  DFFQXL \block_reg[6][98]  ( .D(n971), .CK(clk), .Q(\block[6][98] ) );
  CLKMX2X2 \block_reg[6][97]/U3  ( .A(\block[6][97] ), .B(block_next[97]), 
        .S0(n1520), .Y(n970) );
  DFFQXL \block_reg[6][97]  ( .D(n970), .CK(clk), .Q(\block[6][97] ) );
  CLKMX2X2 \block_reg[5][103]/U3  ( .A(\block[5][103] ), .B(block_next[103]), 
        .S0(n1536), .Y(n969) );
  DFFQXL \block_reg[5][103]  ( .D(n969), .CK(clk), .Q(\block[5][103] ) );
  CLKMX2X2 \block_reg[5][102]/U3  ( .A(\block[5][102] ), .B(block_next[102]), 
        .S0(n1536), .Y(n968) );
  DFFQXL \block_reg[5][102]  ( .D(n968), .CK(clk), .Q(\block[5][102] ) );
  CLKMX2X2 \block_reg[5][101]/U3  ( .A(\block[5][101] ), .B(block_next[101]), 
        .S0(n1536), .Y(n967) );
  DFFQXL \block_reg[5][101]  ( .D(n967), .CK(clk), .Q(\block[5][101] ) );
  CLKMX2X2 \block_reg[5][100]/U3  ( .A(\block[5][100] ), .B(block_next[100]), 
        .S0(n1536), .Y(n966) );
  DFFQXL \block_reg[5][100]  ( .D(n966), .CK(clk), .Q(\block[5][100] ) );
  DFFQXL \block_reg[5][99]  ( .D(n965), .CK(clk), .Q(\block[5][99] ) );
  DFFQXL \block_reg[5][96]  ( .D(n964), .CK(clk), .Q(\block[5][96] ) );
  CLKMX2X2 \block_reg[4][103]/U3  ( .A(\block[4][103] ), .B(block_next[103]), 
        .S0(n1553), .Y(n963) );
  DFFQXL \block_reg[4][103]  ( .D(n963), .CK(clk), .Q(\block[4][103] ) );
  CLKMX2X2 \block_reg[4][102]/U3  ( .A(\block[4][102] ), .B(block_next[102]), 
        .S0(n1553), .Y(n962) );
  DFFQXL \block_reg[4][102]  ( .D(n962), .CK(clk), .Q(\block[4][102] ) );
  CLKMX2X2 \block_reg[4][101]/U3  ( .A(\block[4][101] ), .B(block_next[101]), 
        .S0(n1553), .Y(n961) );
  DFFQXL \block_reg[4][101]  ( .D(n961), .CK(clk), .Q(\block[4][101] ) );
  CLKMX2X2 \block_reg[4][100]/U3  ( .A(\block[4][100] ), .B(block_next[100]), 
        .S0(n1553), .Y(n960) );
  DFFQXL \block_reg[4][100]  ( .D(n960), .CK(clk), .Q(\block[4][100] ) );
  DFFQXL \block_reg[4][99]  ( .D(n959), .CK(clk), .Q(\block[4][99] ) );
  DFFQXL \block_reg[4][96]  ( .D(n958), .CK(clk), .Q(\block[4][96] ) );
  CLKMX2X2 \block_reg[3][103]/U3  ( .A(\block[3][103] ), .B(block_next[103]), 
        .S0(n1570), .Y(n957) );
  DFFQXL \block_reg[3][103]  ( .D(n957), .CK(clk), .Q(\block[3][103] ) );
  CLKMX2X2 \block_reg[3][102]/U3  ( .A(\block[3][102] ), .B(block_next[102]), 
        .S0(n1570), .Y(n956) );
  DFFQXL \block_reg[3][102]  ( .D(n956), .CK(clk), .Q(\block[3][102] ) );
  CLKMX2X2 \block_reg[3][101]/U3  ( .A(\block[3][101] ), .B(block_next[101]), 
        .S0(n1570), .Y(n955) );
  DFFQXL \block_reg[3][101]  ( .D(n955), .CK(clk), .Q(\block[3][101] ) );
  CLKMX2X2 \block_reg[3][100]/U3  ( .A(\block[3][100] ), .B(block_next[100]), 
        .S0(n1570), .Y(n954) );
  DFFQXL \block_reg[3][100]  ( .D(n954), .CK(clk), .Q(\block[3][100] ) );
  DFFQXL \block_reg[3][99]  ( .D(n953), .CK(clk), .Q(\block[3][99] ) );
  CLKMX2X2 \block_reg[3][97]/U3  ( .A(\block[3][97] ), .B(block_next[97]), 
        .S0(n1570), .Y(n952) );
  DFFQXL \block_reg[3][97]  ( .D(n952), .CK(clk), .Q(\block[3][97] ) );
  DFFQXL \block_reg[3][96]  ( .D(n951), .CK(clk), .Q(\block[3][96] ) );
  CLKMX2X2 \block_reg[2][103]/U3  ( .A(\block[2][103] ), .B(block_next[103]), 
        .S0(n1583), .Y(n950) );
  DFFQXL \block_reg[2][103]  ( .D(n950), .CK(clk), .Q(\block[2][103] ) );
  CLKMX2X2 \block_reg[2][102]/U3  ( .A(\block[2][102] ), .B(block_next[102]), 
        .S0(n1583), .Y(n949) );
  DFFQXL \block_reg[2][102]  ( .D(n949), .CK(clk), .Q(\block[2][102] ) );
  CLKMX2X2 \block_reg[2][101]/U3  ( .A(\block[2][101] ), .B(block_next[101]), 
        .S0(n1583), .Y(n948) );
  DFFQXL \block_reg[2][101]  ( .D(n948), .CK(clk), .Q(\block[2][101] ) );
  CLKMX2X2 \block_reg[2][100]/U3  ( .A(\block[2][100] ), .B(block_next[100]), 
        .S0(n1583), .Y(n947) );
  DFFQXL \block_reg[2][100]  ( .D(n947), .CK(clk), .Q(\block[2][100] ) );
  DFFQXL \block_reg[2][99]  ( .D(n946), .CK(clk), .Q(\block[2][99] ) );
  CLKMX2X2 \block_reg[2][97]/U3  ( .A(\block[2][97] ), .B(block_next[97]), 
        .S0(n1583), .Y(n945) );
  DFFQXL \block_reg[2][97]  ( .D(n945), .CK(clk), .Q(\block[2][97] ) );
  DFFQXL \block_reg[2][96]  ( .D(n944), .CK(clk), .Q(\block[2][96] ) );
  CLKMX2X2 \block_reg[1][103]/U3  ( .A(\block[1][103] ), .B(block_next[103]), 
        .S0(n1597), .Y(n943) );
  DFFQXL \block_reg[1][103]  ( .D(n943), .CK(clk), .Q(\block[1][103] ) );
  CLKMX2X2 \block_reg[1][102]/U3  ( .A(\block[1][102] ), .B(block_next[102]), 
        .S0(n1597), .Y(n942) );
  DFFQXL \block_reg[1][102]  ( .D(n942), .CK(clk), .Q(\block[1][102] ) );
  CLKMX2X2 \block_reg[1][101]/U3  ( .A(\block[1][101] ), .B(block_next[101]), 
        .S0(n1597), .Y(n941) );
  DFFQXL \block_reg[1][101]  ( .D(n941), .CK(clk), .Q(\block[1][101] ) );
  CLKMX2X2 \block_reg[1][100]/U3  ( .A(\block[1][100] ), .B(block_next[100]), 
        .S0(n1597), .Y(n940) );
  DFFQXL \block_reg[1][100]  ( .D(n940), .CK(clk), .Q(\block[1][100] ) );
  DFFQXL \block_reg[1][99]  ( .D(n939), .CK(clk), .Q(\block[1][99] ) );
  CLKMX2X2 \block_reg[1][97]/U3  ( .A(\block[1][97] ), .B(block_next[97]), 
        .S0(n1597), .Y(n938) );
  DFFQXL \block_reg[1][97]  ( .D(n938), .CK(clk), .Q(\block[1][97] ) );
  DFFQXL \block_reg[1][96]  ( .D(n937), .CK(clk), .Q(\block[1][96] ) );
  CLKMX2X2 \block_reg[0][103]/U3  ( .A(\block[0][103] ), .B(block_next[103]), 
        .S0(n1612), .Y(n936) );
  DFFQXL \block_reg[0][103]  ( .D(n936), .CK(clk), .Q(\block[0][103] ) );
  CLKMX2X2 \block_reg[0][102]/U3  ( .A(\block[0][102] ), .B(block_next[102]), 
        .S0(n1612), .Y(n935) );
  DFFQXL \block_reg[0][102]  ( .D(n935), .CK(clk), .Q(\block[0][102] ) );
  CLKMX2X2 \block_reg[0][101]/U3  ( .A(\block[0][101] ), .B(block_next[101]), 
        .S0(n1612), .Y(n934) );
  DFFQXL \block_reg[0][101]  ( .D(n934), .CK(clk), .Q(\block[0][101] ) );
  DFFQXL \block_reg[0][100]  ( .D(n933), .CK(clk), .Q(\block[0][100] ) );
  CLKMX2X2 \block_reg[0][97]/U3  ( .A(\block[0][97] ), .B(block_next[97]), 
        .S0(n1612), .Y(n931) );
  DFFQXL \block_reg[0][97]  ( .D(n931), .CK(clk), .Q(\block[0][97] ) );
  DFFQXL \block_reg[0][96]  ( .D(n930), .CK(clk), .Q(\block[0][96] ) );
  CLKMX2X2 \block_reg[7][95]/U3  ( .A(\block[7][95] ), .B(block_next[95]), 
        .S0(n1505), .Y(n929) );
  DFFQXL \block_reg[7][95]  ( .D(n929), .CK(clk), .Q(\block[7][95] ) );
  CLKMX2X2 \block_reg[7][94]/U3  ( .A(\block[7][94] ), .B(block_next[94]), 
        .S0(n1505), .Y(n928) );
  DFFQXL \block_reg[7][94]  ( .D(n928), .CK(clk), .Q(\block[7][94] ) );
  CLKMX2X2 \block_reg[7][93]/U3  ( .A(\block[7][93] ), .B(block_next[93]), 
        .S0(n1505), .Y(n927) );
  DFFQXL \block_reg[7][93]  ( .D(n927), .CK(clk), .Q(\block[7][93] ) );
  CLKMX2X2 \block_reg[7][92]/U3  ( .A(\block[7][92] ), .B(block_next[92]), 
        .S0(n1505), .Y(n926) );
  DFFQXL \block_reg[7][92]  ( .D(n926), .CK(clk), .Q(\block[7][92] ) );
  CLKMX2X2 \block_reg[7][91]/U3  ( .A(\block[7][91] ), .B(block_next[91]), 
        .S0(n1504), .Y(n925) );
  DFFQXL \block_reg[7][91]  ( .D(n925), .CK(clk), .Q(\block[7][91] ) );
  CLKMX2X2 \block_reg[7][90]/U3  ( .A(\block[7][90] ), .B(block_next[90]), 
        .S0(n1504), .Y(n924) );
  DFFQXL \block_reg[7][90]  ( .D(n924), .CK(clk), .Q(\block[7][90] ) );
  CLKMX2X2 \block_reg[7][89]/U3  ( .A(\block[7][89] ), .B(block_next[89]), 
        .S0(n1504), .Y(n923) );
  DFFQXL \block_reg[7][89]  ( .D(n923), .CK(clk), .Q(\block[7][89] ) );
  CLKMX2X2 \block_reg[7][88]/U3  ( .A(\block[7][88] ), .B(block_next[88]), 
        .S0(n1504), .Y(n922) );
  DFFQXL \block_reg[7][88]  ( .D(n922), .CK(clk), .Q(\block[7][88] ) );
  DFFQXL \block_reg[7][86]  ( .D(n920), .CK(clk), .Q(\block[7][86] ) );
  CLKMX2X2 \block_reg[7][78]/U3  ( .A(\block[7][78] ), .B(block_next[78]), 
        .S0(n1503), .Y(n912) );
  DFFQXL \block_reg[7][78]  ( .D(n912), .CK(clk), .Q(\block[7][78] ) );
  DFFQXL \block_reg[7][76]  ( .D(n910), .CK(clk), .Q(\block[7][76] ) );
  CLKMX2X2 \block_reg[7][75]/U3  ( .A(\block[7][75] ), .B(block_next[75]), 
        .S0(n1503), .Y(n909) );
  DFFQXL \block_reg[7][75]  ( .D(n909), .CK(clk), .Q(\block[7][75] ) );
  DFFQXL \block_reg[7][74]  ( .D(n908), .CK(clk), .Q(\block[7][74] ) );
  DFFQXL \block_reg[7][73]  ( .D(n907), .CK(clk), .Q(\block[7][73] ) );
  DFFQXL \block_reg[7][72]  ( .D(n906), .CK(clk), .Q(\block[7][72] ) );
  CLKMX2X2 \block_reg[6][95]/U3  ( .A(\block[6][95] ), .B(block_next[95]), 
        .S0(n1520), .Y(n905) );
  DFFQXL \block_reg[6][95]  ( .D(n905), .CK(clk), .Q(\block[6][95] ) );
  CLKMX2X2 \block_reg[6][94]/U3  ( .A(\block[6][94] ), .B(block_next[94]), 
        .S0(n1520), .Y(n904) );
  DFFQXL \block_reg[6][94]  ( .D(n904), .CK(clk), .Q(\block[6][94] ) );
  CLKMX2X2 \block_reg[6][93]/U3  ( .A(\block[6][93] ), .B(block_next[93]), 
        .S0(n1520), .Y(n903) );
  DFFQXL \block_reg[6][93]  ( .D(n903), .CK(clk), .Q(\block[6][93] ) );
  CLKMX2X2 \block_reg[6][92]/U3  ( .A(\block[6][92] ), .B(block_next[92]), 
        .S0(n1520), .Y(n902) );
  DFFQXL \block_reg[6][92]  ( .D(n902), .CK(clk), .Q(\block[6][92] ) );
  CLKMX2X2 \block_reg[6][91]/U3  ( .A(\block[6][91] ), .B(block_next[91]), 
        .S0(n1519), .Y(n901) );
  DFFQXL \block_reg[6][91]  ( .D(n901), .CK(clk), .Q(\block[6][91] ) );
  CLKMX2X2 \block_reg[6][90]/U3  ( .A(\block[6][90] ), .B(block_next[90]), 
        .S0(n1519), .Y(n900) );
  DFFQXL \block_reg[6][90]  ( .D(n900), .CK(clk), .Q(\block[6][90] ) );
  CLKMX2X2 \block_reg[6][89]/U3  ( .A(\block[6][89] ), .B(block_next[89]), 
        .S0(n1519), .Y(n899) );
  DFFQXL \block_reg[6][89]  ( .D(n899), .CK(clk), .Q(\block[6][89] ) );
  CLKMX2X2 \block_reg[6][88]/U3  ( .A(\block[6][88] ), .B(block_next[88]), 
        .S0(n1519), .Y(n898) );
  DFFQXL \block_reg[6][88]  ( .D(n898), .CK(clk), .Q(\block[6][88] ) );
  DFFQXL \block_reg[6][87]  ( .D(n897), .CK(clk), .Q(\block[6][87] ) );
  CLKMX2X2 \block_reg[6][86]/U3  ( .A(\block[6][86] ), .B(block_next[86]), 
        .S0(n1519), .Y(n896) );
  DFFQXL \block_reg[6][86]  ( .D(n896), .CK(clk), .Q(\block[6][86] ) );
  DFFQXL \block_reg[6][85]  ( .D(n895), .CK(clk), .Q(\block[6][85] ) );
  DFFQXL \block_reg[6][84]  ( .D(n894), .CK(clk), .Q(\block[6][84] ) );
  DFFQXL \block_reg[6][83]  ( .D(n893), .CK(clk), .Q(\block[6][83] ) );
  DFFQXL \block_reg[6][82]  ( .D(n892), .CK(clk), .Q(\block[6][82] ) );
  DFFQXL \block_reg[6][81]  ( .D(n891), .CK(clk), .Q(\block[6][81] ) );
  DFFQXL \block_reg[6][80]  ( .D(n890), .CK(clk), .Q(\block[6][80] ) );
  DFFQXL \block_reg[6][79]  ( .D(n889), .CK(clk), .Q(\block[6][79] ) );
  CLKMX2X2 \block_reg[6][78]/U3  ( .A(\block[6][78] ), .B(block_next[78]), 
        .S0(n1518), .Y(n888) );
  DFFQXL \block_reg[6][78]  ( .D(n888), .CK(clk), .Q(\block[6][78] ) );
  DFFQXL \block_reg[6][77]  ( .D(n887), .CK(clk), .Q(\block[6][77] ) );
  DFFQXL \block_reg[6][76]  ( .D(n886), .CK(clk), .Q(\block[6][76] ) );
  CLKMX2X2 \block_reg[6][75]/U3  ( .A(\block[6][75] ), .B(block_next[75]), 
        .S0(n1518), .Y(n885) );
  DFFQXL \block_reg[6][75]  ( .D(n885), .CK(clk), .Q(\block[6][75] ) );
  DFFQXL \block_reg[6][74]  ( .D(n884), .CK(clk), .Q(\block[6][74] ) );
  DFFQXL \block_reg[6][73]  ( .D(n883), .CK(clk), .Q(\block[6][73] ) );
  DFFQXL \block_reg[6][72]  ( .D(n882), .CK(clk), .Q(\block[6][72] ) );
  CLKMX2X2 \block_reg[5][95]/U3  ( .A(\block[5][95] ), .B(block_next[95]), 
        .S0(n1536), .Y(n881) );
  DFFQXL \block_reg[5][95]  ( .D(n881), .CK(clk), .Q(\block[5][95] ) );
  CLKMX2X2 \block_reg[5][94]/U3  ( .A(\block[5][94] ), .B(block_next[94]), 
        .S0(n1536), .Y(n880) );
  DFFQXL \block_reg[5][94]  ( .D(n880), .CK(clk), .Q(\block[5][94] ) );
  CLKMX2X2 \block_reg[5][93]/U3  ( .A(\block[5][93] ), .B(block_next[93]), 
        .S0(n1536), .Y(n879) );
  DFFQXL \block_reg[5][93]  ( .D(n879), .CK(clk), .Q(\block[5][93] ) );
  CLKMX2X2 \block_reg[5][92]/U3  ( .A(\block[5][92] ), .B(block_next[92]), 
        .S0(n1536), .Y(n878) );
  DFFQXL \block_reg[5][92]  ( .D(n878), .CK(clk), .Q(\block[5][92] ) );
  CLKMX2X2 \block_reg[5][91]/U3  ( .A(\block[5][91] ), .B(block_next[91]), 
        .S0(n1535), .Y(n877) );
  DFFQXL \block_reg[5][91]  ( .D(n877), .CK(clk), .Q(\block[5][91] ) );
  CLKMX2X2 \block_reg[5][90]/U3  ( .A(\block[5][90] ), .B(block_next[90]), 
        .S0(n1535), .Y(n876) );
  DFFQXL \block_reg[5][90]  ( .D(n876), .CK(clk), .Q(\block[5][90] ) );
  CLKMX2X2 \block_reg[5][89]/U3  ( .A(\block[5][89] ), .B(block_next[89]), 
        .S0(n1535), .Y(n875) );
  DFFQXL \block_reg[5][89]  ( .D(n875), .CK(clk), .Q(\block[5][89] ) );
  CLKMX2X2 \block_reg[5][88]/U3  ( .A(\block[5][88] ), .B(block_next[88]), 
        .S0(n1535), .Y(n874) );
  DFFQXL \block_reg[5][88]  ( .D(n874), .CK(clk), .Q(\block[5][88] ) );
  DFFQXL \block_reg[5][87]  ( .D(n873), .CK(clk), .Q(\block[5][87] ) );
  CLKMX2X2 \block_reg[5][86]/U3  ( .A(\block[5][86] ), .B(block_next[86]), 
        .S0(n1535), .Y(n872) );
  DFFQXL \block_reg[5][86]  ( .D(n872), .CK(clk), .Q(\block[5][86] ) );
  DFFQXL \block_reg[5][85]  ( .D(n871), .CK(clk), .Q(\block[5][85] ) );
  DFFQXL \block_reg[5][84]  ( .D(n870), .CK(clk), .Q(\block[5][84] ) );
  DFFQXL \block_reg[5][83]  ( .D(n869), .CK(clk), .Q(\block[5][83] ) );
  DFFQXL \block_reg[5][82]  ( .D(n868), .CK(clk), .Q(\block[5][82] ) );
  DFFQXL \block_reg[5][81]  ( .D(n867), .CK(clk), .Q(\block[5][81] ) );
  DFFQXL \block_reg[5][80]  ( .D(n866), .CK(clk), .Q(\block[5][80] ) );
  DFFQXL \block_reg[5][79]  ( .D(n865), .CK(clk), .Q(\block[5][79] ) );
  CLKMX2X2 \block_reg[5][78]/U3  ( .A(\block[5][78] ), .B(block_next[78]), 
        .S0(n1534), .Y(n864) );
  DFFQXL \block_reg[5][78]  ( .D(n864), .CK(clk), .Q(\block[5][78] ) );
  DFFQXL \block_reg[5][77]  ( .D(n863), .CK(clk), .Q(\block[5][77] ) );
  DFFQXL \block_reg[5][76]  ( .D(n862), .CK(clk), .Q(\block[5][76] ) );
  CLKMX2X2 \block_reg[5][75]/U3  ( .A(\block[5][75] ), .B(block_next[75]), 
        .S0(n1534), .Y(n861) );
  DFFQXL \block_reg[5][75]  ( .D(n861), .CK(clk), .Q(\block[5][75] ) );
  DFFQXL \block_reg[5][74]  ( .D(n860), .CK(clk), .Q(\block[5][74] ) );
  DFFQXL \block_reg[5][73]  ( .D(n859), .CK(clk), .Q(\block[5][73] ) );
  DFFQXL \block_reg[5][72]  ( .D(n858), .CK(clk), .Q(\block[5][72] ) );
  CLKMX2X2 \block_reg[4][95]/U3  ( .A(\block[4][95] ), .B(block_next[95]), 
        .S0(n1553), .Y(n857) );
  DFFQXL \block_reg[4][95]  ( .D(n857), .CK(clk), .Q(\block[4][95] ) );
  CLKMX2X2 \block_reg[4][94]/U3  ( .A(\block[4][94] ), .B(block_next[94]), 
        .S0(n1553), .Y(n856) );
  DFFQXL \block_reg[4][94]  ( .D(n856), .CK(clk), .Q(\block[4][94] ) );
  CLKMX2X2 \block_reg[4][93]/U3  ( .A(\block[4][93] ), .B(block_next[93]), 
        .S0(n1553), .Y(n855) );
  DFFQXL \block_reg[4][93]  ( .D(n855), .CK(clk), .Q(\block[4][93] ) );
  CLKMX2X2 \block_reg[4][92]/U3  ( .A(\block[4][92] ), .B(block_next[92]), 
        .S0(n1553), .Y(n854) );
  DFFQXL \block_reg[4][92]  ( .D(n854), .CK(clk), .Q(\block[4][92] ) );
  CLKMX2X2 \block_reg[4][91]/U3  ( .A(\block[4][91] ), .B(block_next[91]), 
        .S0(n1552), .Y(n853) );
  DFFQXL \block_reg[4][91]  ( .D(n853), .CK(clk), .Q(\block[4][91] ) );
  CLKMX2X2 \block_reg[4][90]/U3  ( .A(\block[4][90] ), .B(block_next[90]), 
        .S0(n1552), .Y(n852) );
  DFFQXL \block_reg[4][90]  ( .D(n852), .CK(clk), .Q(\block[4][90] ) );
  CLKMX2X2 \block_reg[4][89]/U3  ( .A(\block[4][89] ), .B(block_next[89]), 
        .S0(n1552), .Y(n851) );
  DFFQXL \block_reg[4][89]  ( .D(n851), .CK(clk), .Q(\block[4][89] ) );
  CLKMX2X2 \block_reg[4][88]/U3  ( .A(\block[4][88] ), .B(block_next[88]), 
        .S0(n1552), .Y(n850) );
  DFFQXL \block_reg[4][88]  ( .D(n850), .CK(clk), .Q(\block[4][88] ) );
  DFFQXL \block_reg[4][87]  ( .D(n849), .CK(clk), .Q(\block[4][87] ) );
  CLKMX2X2 \block_reg[4][86]/U3  ( .A(\block[4][86] ), .B(block_next[86]), 
        .S0(n1552), .Y(n848) );
  DFFQXL \block_reg[4][86]  ( .D(n848), .CK(clk), .Q(\block[4][86] ) );
  DFFQXL \block_reg[4][85]  ( .D(n847), .CK(clk), .Q(\block[4][85] ) );
  DFFQXL \block_reg[4][84]  ( .D(n846), .CK(clk), .Q(\block[4][84] ) );
  DFFQXL \block_reg[4][83]  ( .D(n845), .CK(clk), .Q(\block[4][83] ) );
  DFFQXL \block_reg[4][82]  ( .D(n844), .CK(clk), .Q(\block[4][82] ) );
  DFFQXL \block_reg[4][81]  ( .D(n843), .CK(clk), .Q(\block[4][81] ) );
  DFFQXL \block_reg[4][80]  ( .D(n842), .CK(clk), .Q(\block[4][80] ) );
  DFFQXL \block_reg[4][79]  ( .D(n841), .CK(clk), .Q(\block[4][79] ) );
  CLKMX2X2 \block_reg[4][78]/U3  ( .A(\block[4][78] ), .B(block_next[78]), 
        .S0(n1551), .Y(n840) );
  DFFQXL \block_reg[4][78]  ( .D(n840), .CK(clk), .Q(\block[4][78] ) );
  DFFQXL \block_reg[4][77]  ( .D(n839), .CK(clk), .Q(\block[4][77] ) );
  DFFQXL \block_reg[4][76]  ( .D(n838), .CK(clk), .Q(\block[4][76] ) );
  CLKMX2X2 \block_reg[4][75]/U3  ( .A(\block[4][75] ), .B(block_next[75]), 
        .S0(n1551), .Y(n837) );
  DFFQXL \block_reg[4][75]  ( .D(n837), .CK(clk), .Q(\block[4][75] ) );
  DFFQXL \block_reg[4][74]  ( .D(n836), .CK(clk), .Q(\block[4][74] ) );
  DFFQXL \block_reg[4][73]  ( .D(n835), .CK(clk), .Q(\block[4][73] ) );
  DFFQXL \block_reg[4][72]  ( .D(n834), .CK(clk), .Q(\block[4][72] ) );
  CLKMX2X2 \block_reg[3][95]/U3  ( .A(\block[3][95] ), .B(block_next[95]), 
        .S0(n1570), .Y(n833) );
  DFFQXL \block_reg[3][95]  ( .D(n833), .CK(clk), .Q(\block[3][95] ) );
  CLKMX2X2 \block_reg[3][94]/U3  ( .A(\block[3][94] ), .B(block_next[94]), 
        .S0(n1570), .Y(n832) );
  DFFQXL \block_reg[3][94]  ( .D(n832), .CK(clk), .Q(\block[3][94] ) );
  CLKMX2X2 \block_reg[3][93]/U3  ( .A(\block[3][93] ), .B(block_next[93]), 
        .S0(n1570), .Y(n831) );
  DFFQXL \block_reg[3][93]  ( .D(n831), .CK(clk), .Q(\block[3][93] ) );
  CLKMX2X2 \block_reg[3][92]/U3  ( .A(\block[3][92] ), .B(block_next[92]), 
        .S0(n1570), .Y(n830) );
  DFFQXL \block_reg[3][92]  ( .D(n830), .CK(clk), .Q(\block[3][92] ) );
  CLKMX2X2 \block_reg[3][91]/U3  ( .A(\block[3][91] ), .B(block_next[91]), 
        .S0(n1569), .Y(n829) );
  DFFQXL \block_reg[3][91]  ( .D(n829), .CK(clk), .Q(\block[3][91] ) );
  CLKMX2X2 \block_reg[3][90]/U3  ( .A(\block[3][90] ), .B(block_next[90]), 
        .S0(n1569), .Y(n828) );
  DFFQXL \block_reg[3][90]  ( .D(n828), .CK(clk), .Q(\block[3][90] ) );
  CLKMX2X2 \block_reg[3][89]/U3  ( .A(\block[3][89] ), .B(block_next[89]), 
        .S0(n1569), .Y(n827) );
  DFFQXL \block_reg[3][89]  ( .D(n827), .CK(clk), .Q(\block[3][89] ) );
  CLKMX2X2 \block_reg[3][88]/U3  ( .A(\block[3][88] ), .B(block_next[88]), 
        .S0(n1569), .Y(n826) );
  DFFQXL \block_reg[3][88]  ( .D(n826), .CK(clk), .Q(\block[3][88] ) );
  DFFQXL \block_reg[3][87]  ( .D(n825), .CK(clk), .Q(\block[3][87] ) );
  CLKMX2X2 \block_reg[3][86]/U3  ( .A(\block[3][86] ), .B(block_next[86]), 
        .S0(n1569), .Y(n824) );
  DFFQXL \block_reg[3][86]  ( .D(n824), .CK(clk), .Q(\block[3][86] ) );
  DFFQXL \block_reg[3][85]  ( .D(n823), .CK(clk), .Q(\block[3][85] ) );
  DFFQXL \block_reg[3][84]  ( .D(n822), .CK(clk), .Q(\block[3][84] ) );
  DFFQXL \block_reg[3][83]  ( .D(n821), .CK(clk), .Q(\block[3][83] ) );
  DFFQXL \block_reg[3][82]  ( .D(n820), .CK(clk), .Q(\block[3][82] ) );
  DFFQXL \block_reg[3][81]  ( .D(n819), .CK(clk), .Q(\block[3][81] ) );
  DFFQXL \block_reg[3][80]  ( .D(n818), .CK(clk), .Q(\block[3][80] ) );
  DFFQXL \block_reg[3][79]  ( .D(n817), .CK(clk), .Q(\block[3][79] ) );
  CLKMX2X2 \block_reg[3][78]/U3  ( .A(\block[3][78] ), .B(block_next[78]), 
        .S0(n1568), .Y(n816) );
  DFFQXL \block_reg[3][78]  ( .D(n816), .CK(clk), .Q(\block[3][78] ) );
  DFFQXL \block_reg[3][77]  ( .D(n815), .CK(clk), .Q(\block[3][77] ) );
  DFFQXL \block_reg[3][76]  ( .D(n814), .CK(clk), .Q(\block[3][76] ) );
  CLKMX2X2 \block_reg[3][75]/U3  ( .A(\block[3][75] ), .B(block_next[75]), 
        .S0(n1568), .Y(n813) );
  DFFQXL \block_reg[3][75]  ( .D(n813), .CK(clk), .Q(\block[3][75] ) );
  DFFQXL \block_reg[3][74]  ( .D(n812), .CK(clk), .Q(\block[3][74] ) );
  DFFQXL \block_reg[3][73]  ( .D(n811), .CK(clk), .Q(\block[3][73] ) );
  DFFQXL \block_reg[3][72]  ( .D(n810), .CK(clk), .Q(\block[3][72] ) );
  CLKMX2X2 \block_reg[2][95]/U3  ( .A(\block[2][95] ), .B(block_next[95]), 
        .S0(n1583), .Y(n809) );
  DFFQXL \block_reg[2][95]  ( .D(n809), .CK(clk), .Q(\block[2][95] ) );
  CLKMX2X2 \block_reg[2][94]/U3  ( .A(\block[2][94] ), .B(block_next[94]), 
        .S0(n1583), .Y(n808) );
  DFFQXL \block_reg[2][94]  ( .D(n808), .CK(clk), .Q(\block[2][94] ) );
  CLKMX2X2 \block_reg[2][93]/U3  ( .A(\block[2][93] ), .B(block_next[93]), 
        .S0(n1583), .Y(n807) );
  DFFQXL \block_reg[2][93]  ( .D(n807), .CK(clk), .Q(\block[2][93] ) );
  CLKMX2X2 \block_reg[2][92]/U3  ( .A(\block[2][92] ), .B(block_next[92]), 
        .S0(n1583), .Y(n806) );
  DFFQXL \block_reg[2][92]  ( .D(n806), .CK(clk), .Q(\block[2][92] ) );
  CLKMX2X2 \block_reg[2][91]/U3  ( .A(\block[2][91] ), .B(block_next[91]), 
        .S0(n1582), .Y(n805) );
  DFFQXL \block_reg[2][91]  ( .D(n805), .CK(clk), .Q(\block[2][91] ) );
  CLKMX2X2 \block_reg[2][90]/U3  ( .A(\block[2][90] ), .B(block_next[90]), 
        .S0(n1582), .Y(n804) );
  DFFQXL \block_reg[2][90]  ( .D(n804), .CK(clk), .Q(\block[2][90] ) );
  CLKMX2X2 \block_reg[2][89]/U3  ( .A(\block[2][89] ), .B(block_next[89]), 
        .S0(n1582), .Y(n803) );
  DFFQXL \block_reg[2][89]  ( .D(n803), .CK(clk), .Q(\block[2][89] ) );
  CLKMX2X2 \block_reg[2][88]/U3  ( .A(\block[2][88] ), .B(block_next[88]), 
        .S0(n1582), .Y(n802) );
  DFFQXL \block_reg[2][88]  ( .D(n802), .CK(clk), .Q(\block[2][88] ) );
  DFFQXL \block_reg[2][87]  ( .D(n801), .CK(clk), .Q(\block[2][87] ) );
  CLKMX2X2 \block_reg[2][86]/U3  ( .A(\block[2][86] ), .B(block_next[86]), 
        .S0(n1582), .Y(n800) );
  DFFQXL \block_reg[2][86]  ( .D(n800), .CK(clk), .Q(\block[2][86] ) );
  DFFQXL \block_reg[2][85]  ( .D(n799), .CK(clk), .Q(\block[2][85] ) );
  DFFQXL \block_reg[2][84]  ( .D(n798), .CK(clk), .Q(\block[2][84] ) );
  DFFQXL \block_reg[2][83]  ( .D(n797), .CK(clk), .Q(\block[2][83] ) );
  DFFQXL \block_reg[2][82]  ( .D(n796), .CK(clk), .Q(\block[2][82] ) );
  DFFQXL \block_reg[2][81]  ( .D(n795), .CK(clk), .Q(\block[2][81] ) );
  DFFQXL \block_reg[2][80]  ( .D(n794), .CK(clk), .Q(\block[2][80] ) );
  DFFQXL \block_reg[2][79]  ( .D(n793), .CK(clk), .Q(\block[2][79] ) );
  CLKMX2X2 \block_reg[2][78]/U3  ( .A(\block[2][78] ), .B(block_next[78]), 
        .S0(n1581), .Y(n792) );
  DFFQXL \block_reg[2][78]  ( .D(n792), .CK(clk), .Q(\block[2][78] ) );
  DFFQXL \block_reg[2][77]  ( .D(n791), .CK(clk), .Q(\block[2][77] ) );
  CLKMX2X2 \block_reg[1][95]/U3  ( .A(\block[1][95] ), .B(block_next[95]), 
        .S0(n1597), .Y(n785) );
  DFFQXL \block_reg[1][95]  ( .D(n785), .CK(clk), .Q(\block[1][95] ) );
  CLKMX2X2 \block_reg[1][94]/U3  ( .A(\block[1][94] ), .B(block_next[94]), 
        .S0(n1597), .Y(n784) );
  DFFQXL \block_reg[1][94]  ( .D(n784), .CK(clk), .Q(\block[1][94] ) );
  CLKMX2X2 \block_reg[1][93]/U3  ( .A(\block[1][93] ), .B(block_next[93]), 
        .S0(n1597), .Y(n783) );
  DFFQXL \block_reg[1][93]  ( .D(n783), .CK(clk), .Q(\block[1][93] ) );
  CLKMX2X2 \block_reg[1][92]/U3  ( .A(\block[1][92] ), .B(block_next[92]), 
        .S0(n1597), .Y(n782) );
  DFFQXL \block_reg[1][92]  ( .D(n782), .CK(clk), .Q(\block[1][92] ) );
  CLKMX2X2 \block_reg[1][91]/U3  ( .A(\block[1][91] ), .B(block_next[91]), 
        .S0(n1596), .Y(n781) );
  DFFQXL \block_reg[1][91]  ( .D(n781), .CK(clk), .Q(\block[1][91] ) );
  CLKMX2X2 \block_reg[1][90]/U3  ( .A(\block[1][90] ), .B(block_next[90]), 
        .S0(n1596), .Y(n780) );
  DFFQXL \block_reg[1][90]  ( .D(n780), .CK(clk), .Q(\block[1][90] ) );
  CLKMX2X2 \block_reg[1][89]/U3  ( .A(\block[1][89] ), .B(block_next[89]), 
        .S0(n1596), .Y(n779) );
  DFFQXL \block_reg[1][89]  ( .D(n779), .CK(clk), .Q(\block[1][89] ) );
  CLKMX2X2 \block_reg[1][88]/U3  ( .A(\block[1][88] ), .B(block_next[88]), 
        .S0(n1596), .Y(n778) );
  DFFQXL \block_reg[1][88]  ( .D(n778), .CK(clk), .Q(\block[1][88] ) );
  DFFQXL \block_reg[1][87]  ( .D(n777), .CK(clk), .Q(\block[1][87] ) );
  CLKMX2X2 \block_reg[1][86]/U3  ( .A(\block[1][86] ), .B(block_next[86]), 
        .S0(n1596), .Y(n776) );
  DFFQXL \block_reg[1][86]  ( .D(n776), .CK(clk), .Q(\block[1][86] ) );
  DFFQXL \block_reg[1][85]  ( .D(n775), .CK(clk), .Q(\block[1][85] ) );
  DFFQXL \block_reg[1][84]  ( .D(n774), .CK(clk), .Q(\block[1][84] ) );
  DFFQXL \block_reg[1][83]  ( .D(n773), .CK(clk), .Q(\block[1][83] ) );
  DFFQXL \block_reg[1][82]  ( .D(n772), .CK(clk), .Q(\block[1][82] ) );
  DFFQXL \block_reg[1][81]  ( .D(n771), .CK(clk), .Q(\block[1][81] ) );
  DFFQXL \block_reg[1][80]  ( .D(n770), .CK(clk), .Q(\block[1][80] ) );
  DFFQXL \block_reg[1][79]  ( .D(n769), .CK(clk), .Q(\block[1][79] ) );
  CLKMX2X2 \block_reg[1][78]/U3  ( .A(\block[1][78] ), .B(block_next[78]), 
        .S0(n1595), .Y(n768) );
  DFFQXL \block_reg[1][78]  ( .D(n768), .CK(clk), .Q(\block[1][78] ) );
  DFFQXL \block_reg[1][77]  ( .D(n767), .CK(clk), .Q(\block[1][77] ) );
  DFFQXL \block_reg[1][76]  ( .D(n766), .CK(clk), .Q(\block[1][76] ) );
  CLKMX2X2 \block_reg[1][75]/U3  ( .A(\block[1][75] ), .B(block_next[75]), 
        .S0(n1595), .Y(n765) );
  DFFQXL \block_reg[1][75]  ( .D(n765), .CK(clk), .Q(\block[1][75] ) );
  DFFQXL \block_reg[1][74]  ( .D(n764), .CK(clk), .Q(\block[1][74] ) );
  DFFQXL \block_reg[1][73]  ( .D(n763), .CK(clk), .Q(\block[1][73] ) );
  DFFQXL \block_reg[1][72]  ( .D(n762), .CK(clk), .Q(\block[1][72] ) );
  CLKMX2X2 \block_reg[0][95]/U3  ( .A(\block[0][95] ), .B(block_next[95]), 
        .S0(n1612), .Y(n761) );
  DFFQXL \block_reg[0][95]  ( .D(n761), .CK(clk), .Q(\block[0][95] ) );
  CLKMX2X2 \block_reg[0][94]/U3  ( .A(\block[0][94] ), .B(block_next[94]), 
        .S0(n1612), .Y(n760) );
  DFFQXL \block_reg[0][94]  ( .D(n760), .CK(clk), .Q(\block[0][94] ) );
  CLKMX2X2 \block_reg[0][93]/U3  ( .A(\block[0][93] ), .B(block_next[93]), 
        .S0(n1612), .Y(n759) );
  DFFQXL \block_reg[0][93]  ( .D(n759), .CK(clk), .Q(\block[0][93] ) );
  CLKMX2X2 \block_reg[0][92]/U3  ( .A(\block[0][92] ), .B(block_next[92]), 
        .S0(n1612), .Y(n758) );
  DFFQXL \block_reg[0][92]  ( .D(n758), .CK(clk), .Q(\block[0][92] ) );
  CLKMX2X2 \block_reg[0][91]/U3  ( .A(\block[0][91] ), .B(block_next[91]), 
        .S0(n1611), .Y(n757) );
  DFFQXL \block_reg[0][91]  ( .D(n757), .CK(clk), .Q(\block[0][91] ) );
  CLKMX2X2 \block_reg[0][90]/U3  ( .A(\block[0][90] ), .B(block_next[90]), 
        .S0(n1611), .Y(n756) );
  DFFQXL \block_reg[0][90]  ( .D(n756), .CK(clk), .Q(\block[0][90] ) );
  CLKMX2X2 \block_reg[0][89]/U3  ( .A(\block[0][89] ), .B(block_next[89]), 
        .S0(n1611), .Y(n755) );
  DFFQXL \block_reg[0][89]  ( .D(n755), .CK(clk), .Q(\block[0][89] ) );
  CLKMX2X2 \block_reg[0][88]/U3  ( .A(\block[0][88] ), .B(block_next[88]), 
        .S0(n1611), .Y(n754) );
  DFFQXL \block_reg[0][88]  ( .D(n754), .CK(clk), .Q(\block[0][88] ) );
  DFFQXL \block_reg[0][87]  ( .D(n753), .CK(clk), .Q(\block[0][87] ) );
  CLKMX2X2 \block_reg[0][86]/U3  ( .A(\block[0][86] ), .B(block_next[86]), 
        .S0(n1611), .Y(n752) );
  DFFQXL \block_reg[0][86]  ( .D(n752), .CK(clk), .Q(\block[0][86] ) );
  DFFQXL \block_reg[0][85]  ( .D(n751), .CK(clk), .Q(\block[0][85] ) );
  DFFQXL \block_reg[0][84]  ( .D(n750), .CK(clk), .Q(\block[0][84] ) );
  DFFQXL \block_reg[0][83]  ( .D(n749), .CK(clk), .Q(\block[0][83] ) );
  DFFQXL \block_reg[0][82]  ( .D(n748), .CK(clk), .Q(\block[0][82] ) );
  DFFQXL \block_reg[0][81]  ( .D(n747), .CK(clk), .Q(\block[0][81] ) );
  DFFQXL \block_reg[0][80]  ( .D(n746), .CK(clk), .Q(\block[0][80] ) );
  DFFQXL \block_reg[0][79]  ( .D(n745), .CK(clk), .Q(\block[0][79] ) );
  CLKMX2X2 \block_reg[0][78]/U3  ( .A(\block[0][78] ), .B(block_next[78]), 
        .S0(n1610), .Y(n744) );
  DFFQXL \block_reg[0][78]  ( .D(n744), .CK(clk), .Q(\block[0][78] ) );
  DFFQXL \block_reg[0][77]  ( .D(n743), .CK(clk), .Q(\block[0][77] ) );
  DFFQXL \block_reg[0][76]  ( .D(n742), .CK(clk), .Q(\block[0][76] ) );
  CLKMX2X2 \block_reg[0][75]/U3  ( .A(\block[0][75] ), .B(block_next[75]), 
        .S0(n1610), .Y(n741) );
  DFFQXL \block_reg[0][75]  ( .D(n741), .CK(clk), .Q(\block[0][75] ) );
  DFFQXL \block_reg[0][74]  ( .D(n740), .CK(clk), .Q(\block[0][74] ) );
  DFFQXL \block_reg[0][73]  ( .D(n739), .CK(clk), .Q(\block[0][73] ) );
  DFFQXL \block_reg[0][72]  ( .D(n738), .CK(clk), .Q(\block[0][72] ) );
  CLKMX2X2 \block_reg[7][115]/U3  ( .A(\block[7][115] ), .B(block_next[115]), 
        .S0(n1506), .Y(n737) );
  DFFQXL \block_reg[7][115]  ( .D(n737), .CK(clk), .Q(\block[7][115] ) );
  CLKMX2X2 \block_reg[7][114]/U3  ( .A(\block[7][114] ), .B(block_next[114]), 
        .S0(n1506), .Y(n736) );
  DFFQXL \block_reg[7][114]  ( .D(n736), .CK(clk), .Q(\block[7][114] ) );
  CLKMX2X2 \block_reg[7][113]/U3  ( .A(\block[7][113] ), .B(block_next[113]), 
        .S0(n1506), .Y(n735) );
  DFFQXL \block_reg[7][113]  ( .D(n735), .CK(clk), .Q(\block[7][113] ) );
  CLKMX2X2 \block_reg[7][112]/U3  ( .A(\block[7][112] ), .B(block_next[112]), 
        .S0(n1506), .Y(n734) );
  DFFQXL \block_reg[7][112]  ( .D(n734), .CK(clk), .Q(\block[7][112] ) );
  CLKMX2X2 \block_reg[7][111]/U3  ( .A(\block[7][111] ), .B(block_next[111]), 
        .S0(n1506), .Y(n733) );
  DFFQXL \block_reg[7][111]  ( .D(n733), .CK(clk), .Q(\block[7][111] ) );
  CLKMX2X2 \block_reg[7][110]/U3  ( .A(\block[7][110] ), .B(block_next[110]), 
        .S0(n1506), .Y(n732) );
  DFFQXL \block_reg[7][110]  ( .D(n732), .CK(clk), .Q(\block[7][110] ) );
  CLKMX2X2 \block_reg[7][109]/U3  ( .A(\block[7][109] ), .B(block_next[109]), 
        .S0(n1506), .Y(n731) );
  DFFQXL \block_reg[7][109]  ( .D(n731), .CK(clk), .Q(\block[7][109] ) );
  CLKMX2X2 \block_reg[7][108]/U3  ( .A(\block[7][108] ), .B(block_next[108]), 
        .S0(n1506), .Y(n730) );
  DFFQXL \block_reg[7][108]  ( .D(n730), .CK(clk), .Q(\block[7][108] ) );
  CLKMX2X2 \block_reg[7][107]/U3  ( .A(\block[7][107] ), .B(block_next[107]), 
        .S0(n1506), .Y(n729) );
  DFFQXL \block_reg[7][107]  ( .D(n729), .CK(clk), .Q(\block[7][107] ) );
  CLKMX2X2 \block_reg[7][105]/U3  ( .A(\block[7][105] ), .B(block_next[105]), 
        .S0(n1506), .Y(n728) );
  DFFQXL \block_reg[7][105]  ( .D(n728), .CK(clk), .Q(\block[7][105] ) );
  CLKMX2X2 \block_reg[6][115]/U3  ( .A(\block[6][115] ), .B(block_next[115]), 
        .S0(n1521), .Y(n727) );
  DFFQXL \block_reg[6][115]  ( .D(n727), .CK(clk), .Q(\block[6][115] ) );
  CLKMX2X2 \block_reg[6][114]/U3  ( .A(\block[6][114] ), .B(block_next[114]), 
        .S0(n1521), .Y(n726) );
  DFFQXL \block_reg[6][114]  ( .D(n726), .CK(clk), .Q(\block[6][114] ) );
  CLKMX2X2 \block_reg[6][113]/U3  ( .A(\block[6][113] ), .B(block_next[113]), 
        .S0(n1521), .Y(n725) );
  DFFQXL \block_reg[6][113]  ( .D(n725), .CK(clk), .Q(\block[6][113] ) );
  CLKMX2X2 \block_reg[6][112]/U3  ( .A(\block[6][112] ), .B(block_next[112]), 
        .S0(n1521), .Y(n724) );
  DFFQXL \block_reg[6][112]  ( .D(n724), .CK(clk), .Q(\block[6][112] ) );
  CLKMX2X2 \block_reg[6][111]/U3  ( .A(\block[6][111] ), .B(block_next[111]), 
        .S0(n1521), .Y(n723) );
  DFFQXL \block_reg[6][111]  ( .D(n723), .CK(clk), .Q(\block[6][111] ) );
  CLKMX2X2 \block_reg[6][110]/U3  ( .A(\block[6][110] ), .B(block_next[110]), 
        .S0(n1521), .Y(n722) );
  DFFQXL \block_reg[6][110]  ( .D(n722), .CK(clk), .Q(\block[6][110] ) );
  CLKMX2X2 \block_reg[6][109]/U3  ( .A(\block[6][109] ), .B(block_next[109]), 
        .S0(n1521), .Y(n721) );
  DFFQXL \block_reg[6][109]  ( .D(n721), .CK(clk), .Q(\block[6][109] ) );
  CLKMX2X2 \block_reg[6][108]/U3  ( .A(\block[6][108] ), .B(block_next[108]), 
        .S0(n1521), .Y(n720) );
  DFFQXL \block_reg[6][108]  ( .D(n720), .CK(clk), .Q(\block[6][108] ) );
  CLKMX2X2 \block_reg[6][107]/U3  ( .A(\block[6][107] ), .B(block_next[107]), 
        .S0(n1521), .Y(n719) );
  DFFQXL \block_reg[6][107]  ( .D(n719), .CK(clk), .Q(\block[6][107] ) );
  CLKMX2X2 \block_reg[6][105]/U3  ( .A(\block[6][105] ), .B(block_next[105]), 
        .S0(n1521), .Y(n718) );
  DFFQXL \block_reg[6][105]  ( .D(n718), .CK(clk), .Q(\block[6][105] ) );
  CLKMX2X2 \block_reg[5][115]/U3  ( .A(\block[5][115] ), .B(block_next[115]), 
        .S0(n1537), .Y(n717) );
  DFFQXL \block_reg[5][115]  ( .D(n717), .CK(clk), .Q(\block[5][115] ) );
  CLKMX2X2 \block_reg[5][114]/U3  ( .A(\block[5][114] ), .B(block_next[114]), 
        .S0(n1537), .Y(n716) );
  DFFQXL \block_reg[5][114]  ( .D(n716), .CK(clk), .Q(\block[5][114] ) );
  CLKMX2X2 \block_reg[5][113]/U3  ( .A(\block[5][113] ), .B(block_next[113]), 
        .S0(n1537), .Y(n715) );
  DFFQXL \block_reg[5][113]  ( .D(n715), .CK(clk), .Q(\block[5][113] ) );
  CLKMX2X2 \block_reg[5][112]/U3  ( .A(\block[5][112] ), .B(block_next[112]), 
        .S0(n1537), .Y(n714) );
  DFFQXL \block_reg[5][112]  ( .D(n714), .CK(clk), .Q(\block[5][112] ) );
  CLKMX2X2 \block_reg[5][111]/U3  ( .A(\block[5][111] ), .B(block_next[111]), 
        .S0(n1537), .Y(n713) );
  DFFQXL \block_reg[5][111]  ( .D(n713), .CK(clk), .Q(\block[5][111] ) );
  CLKMX2X2 \block_reg[5][110]/U3  ( .A(\block[5][110] ), .B(block_next[110]), 
        .S0(n1537), .Y(n712) );
  DFFQXL \block_reg[5][110]  ( .D(n712), .CK(clk), .Q(\block[5][110] ) );
  CLKMX2X2 \block_reg[5][109]/U3  ( .A(\block[5][109] ), .B(block_next[109]), 
        .S0(n1537), .Y(n711) );
  DFFQXL \block_reg[5][109]  ( .D(n711), .CK(clk), .Q(\block[5][109] ) );
  CLKMX2X2 \block_reg[5][108]/U3  ( .A(\block[5][108] ), .B(block_next[108]), 
        .S0(n1537), .Y(n710) );
  DFFQXL \block_reg[5][108]  ( .D(n710), .CK(clk), .Q(\block[5][108] ) );
  CLKMX2X2 \block_reg[5][107]/U3  ( .A(\block[5][107] ), .B(block_next[107]), 
        .S0(n1537), .Y(n709) );
  DFFQXL \block_reg[5][107]  ( .D(n709), .CK(clk), .Q(\block[5][107] ) );
  CLKMX2X2 \block_reg[5][105]/U3  ( .A(\block[5][105] ), .B(block_next[105]), 
        .S0(n1537), .Y(n708) );
  DFFQXL \block_reg[5][105]  ( .D(n708), .CK(clk), .Q(\block[5][105] ) );
  CLKMX2X2 \block_reg[4][115]/U3  ( .A(\block[4][115] ), .B(block_next[115]), 
        .S0(n1554), .Y(n707) );
  DFFQXL \block_reg[4][115]  ( .D(n707), .CK(clk), .Q(\block[4][115] ) );
  CLKMX2X2 \block_reg[4][114]/U3  ( .A(\block[4][114] ), .B(block_next[114]), 
        .S0(n1554), .Y(n706) );
  DFFQXL \block_reg[4][114]  ( .D(n706), .CK(clk), .Q(\block[4][114] ) );
  CLKMX2X2 \block_reg[4][113]/U3  ( .A(\block[4][113] ), .B(block_next[113]), 
        .S0(n1554), .Y(n705) );
  DFFQXL \block_reg[4][113]  ( .D(n705), .CK(clk), .Q(\block[4][113] ) );
  CLKMX2X2 \block_reg[4][112]/U3  ( .A(\block[4][112] ), .B(block_next[112]), 
        .S0(n1554), .Y(n704) );
  DFFQXL \block_reg[4][112]  ( .D(n704), .CK(clk), .Q(\block[4][112] ) );
  CLKMX2X2 \block_reg[4][111]/U3  ( .A(\block[4][111] ), .B(block_next[111]), 
        .S0(n1554), .Y(n703) );
  DFFQXL \block_reg[4][111]  ( .D(n703), .CK(clk), .Q(\block[4][111] ) );
  CLKMX2X2 \block_reg[4][110]/U3  ( .A(\block[4][110] ), .B(block_next[110]), 
        .S0(n1554), .Y(n702) );
  DFFQXL \block_reg[4][110]  ( .D(n702), .CK(clk), .Q(\block[4][110] ) );
  CLKMX2X2 \block_reg[4][109]/U3  ( .A(\block[4][109] ), .B(block_next[109]), 
        .S0(n1554), .Y(n701) );
  DFFQXL \block_reg[4][109]  ( .D(n701), .CK(clk), .Q(\block[4][109] ) );
  CLKMX2X2 \block_reg[4][108]/U3  ( .A(\block[4][108] ), .B(block_next[108]), 
        .S0(n1554), .Y(n700) );
  DFFQXL \block_reg[4][108]  ( .D(n700), .CK(clk), .Q(\block[4][108] ) );
  CLKMX2X2 \block_reg[4][107]/U3  ( .A(\block[4][107] ), .B(block_next[107]), 
        .S0(n1554), .Y(n699) );
  DFFQXL \block_reg[4][107]  ( .D(n699), .CK(clk), .Q(\block[4][107] ) );
  CLKMX2X2 \block_reg[4][105]/U3  ( .A(\block[4][105] ), .B(block_next[105]), 
        .S0(n1554), .Y(n698) );
  DFFQXL \block_reg[4][105]  ( .D(n698), .CK(clk), .Q(\block[4][105] ) );
  CLKMX2X2 \block_reg[3][115]/U3  ( .A(\block[3][115] ), .B(block_next[115]), 
        .S0(n1571), .Y(n697) );
  DFFQXL \block_reg[3][115]  ( .D(n697), .CK(clk), .Q(\block[3][115] ) );
  CLKMX2X2 \block_reg[3][114]/U3  ( .A(\block[3][114] ), .B(block_next[114]), 
        .S0(n1571), .Y(n696) );
  DFFQXL \block_reg[3][114]  ( .D(n696), .CK(clk), .Q(\block[3][114] ) );
  CLKMX2X2 \block_reg[3][113]/U3  ( .A(\block[3][113] ), .B(block_next[113]), 
        .S0(n1571), .Y(n695) );
  DFFQXL \block_reg[3][113]  ( .D(n695), .CK(clk), .Q(\block[3][113] ) );
  CLKMX2X2 \block_reg[3][112]/U3  ( .A(\block[3][112] ), .B(block_next[112]), 
        .S0(n1571), .Y(n694) );
  DFFQXL \block_reg[3][112]  ( .D(n694), .CK(clk), .Q(\block[3][112] ) );
  CLKMX2X2 \block_reg[3][111]/U3  ( .A(\block[3][111] ), .B(block_next[111]), 
        .S0(n1571), .Y(n693) );
  DFFQXL \block_reg[3][111]  ( .D(n693), .CK(clk), .Q(\block[3][111] ) );
  CLKMX2X2 \block_reg[3][110]/U3  ( .A(\block[3][110] ), .B(block_next[110]), 
        .S0(n1571), .Y(n692) );
  DFFQXL \block_reg[3][110]  ( .D(n692), .CK(clk), .Q(\block[3][110] ) );
  CLKMX2X2 \block_reg[3][109]/U3  ( .A(\block[3][109] ), .B(block_next[109]), 
        .S0(n1571), .Y(n691) );
  DFFQXL \block_reg[3][109]  ( .D(n691), .CK(clk), .Q(\block[3][109] ) );
  CLKMX2X2 \block_reg[3][108]/U3  ( .A(\block[3][108] ), .B(block_next[108]), 
        .S0(n1571), .Y(n690) );
  DFFQXL \block_reg[3][108]  ( .D(n690), .CK(clk), .Q(\block[3][108] ) );
  CLKMX2X2 \block_reg[3][107]/U3  ( .A(\block[3][107] ), .B(block_next[107]), 
        .S0(n1571), .Y(n689) );
  DFFQXL \block_reg[3][107]  ( .D(n689), .CK(clk), .Q(\block[3][107] ) );
  CLKMX2X2 \block_reg[3][105]/U3  ( .A(\block[3][105] ), .B(block_next[105]), 
        .S0(n1571), .Y(n688) );
  DFFQXL \block_reg[3][105]  ( .D(n688), .CK(clk), .Q(\block[3][105] ) );
  CLKMX2X2 \block_reg[2][115]/U3  ( .A(\block[2][115] ), .B(block_next[115]), 
        .S0(n1584), .Y(n687) );
  DFFQXL \block_reg[2][115]  ( .D(n687), .CK(clk), .Q(\block[2][115] ) );
  CLKMX2X2 \block_reg[2][114]/U3  ( .A(\block[2][114] ), .B(block_next[114]), 
        .S0(n1584), .Y(n686) );
  DFFQXL \block_reg[2][114]  ( .D(n686), .CK(clk), .Q(\block[2][114] ) );
  CLKMX2X2 \block_reg[2][113]/U3  ( .A(\block[2][113] ), .B(block_next[113]), 
        .S0(n1584), .Y(n685) );
  DFFQXL \block_reg[2][113]  ( .D(n685), .CK(clk), .Q(\block[2][113] ) );
  CLKMX2X2 \block_reg[2][112]/U3  ( .A(\block[2][112] ), .B(block_next[112]), 
        .S0(n1584), .Y(n684) );
  DFFQXL \block_reg[2][112]  ( .D(n684), .CK(clk), .Q(\block[2][112] ) );
  CLKMX2X2 \block_reg[2][111]/U3  ( .A(\block[2][111] ), .B(block_next[111]), 
        .S0(n1584), .Y(n683) );
  DFFQXL \block_reg[2][111]  ( .D(n683), .CK(clk), .Q(\block[2][111] ) );
  CLKMX2X2 \block_reg[2][110]/U3  ( .A(\block[2][110] ), .B(block_next[110]), 
        .S0(n1584), .Y(n682) );
  DFFQXL \block_reg[2][110]  ( .D(n682), .CK(clk), .Q(\block[2][110] ) );
  CLKMX2X2 \block_reg[2][109]/U3  ( .A(\block[2][109] ), .B(block_next[109]), 
        .S0(n1584), .Y(n681) );
  DFFQXL \block_reg[2][109]  ( .D(n681), .CK(clk), .Q(\block[2][109] ) );
  CLKMX2X2 \block_reg[2][108]/U3  ( .A(\block[2][108] ), .B(block_next[108]), 
        .S0(n1584), .Y(n680) );
  DFFQXL \block_reg[2][108]  ( .D(n680), .CK(clk), .Q(\block[2][108] ) );
  CLKMX2X2 \block_reg[2][107]/U3  ( .A(\block[2][107] ), .B(block_next[107]), 
        .S0(n1584), .Y(n679) );
  DFFQXL \block_reg[2][107]  ( .D(n679), .CK(clk), .Q(\block[2][107] ) );
  CLKMX2X2 \block_reg[2][105]/U3  ( .A(\block[2][105] ), .B(block_next[105]), 
        .S0(n1584), .Y(n678) );
  DFFQXL \block_reg[2][105]  ( .D(n678), .CK(clk), .Q(\block[2][105] ) );
  CLKMX2X2 \block_reg[1][115]/U3  ( .A(\block[1][115] ), .B(block_next[115]), 
        .S0(n1598), .Y(n677) );
  DFFQXL \block_reg[1][115]  ( .D(n677), .CK(clk), .Q(\block[1][115] ) );
  CLKMX2X2 \block_reg[1][114]/U3  ( .A(\block[1][114] ), .B(block_next[114]), 
        .S0(n1598), .Y(n676) );
  DFFQXL \block_reg[1][114]  ( .D(n676), .CK(clk), .Q(\block[1][114] ) );
  CLKMX2X2 \block_reg[1][113]/U3  ( .A(\block[1][113] ), .B(block_next[113]), 
        .S0(n1598), .Y(n675) );
  DFFQXL \block_reg[1][113]  ( .D(n675), .CK(clk), .Q(\block[1][113] ) );
  CLKMX2X2 \block_reg[1][112]/U3  ( .A(\block[1][112] ), .B(block_next[112]), 
        .S0(n1598), .Y(n674) );
  DFFQXL \block_reg[1][112]  ( .D(n674), .CK(clk), .Q(\block[1][112] ) );
  CLKMX2X2 \block_reg[1][111]/U3  ( .A(\block[1][111] ), .B(block_next[111]), 
        .S0(n1598), .Y(n673) );
  DFFQXL \block_reg[1][111]  ( .D(n673), .CK(clk), .Q(\block[1][111] ) );
  CLKMX2X2 \block_reg[1][110]/U3  ( .A(\block[1][110] ), .B(block_next[110]), 
        .S0(n1598), .Y(n672) );
  DFFQXL \block_reg[1][110]  ( .D(n672), .CK(clk), .Q(\block[1][110] ) );
  CLKMX2X2 \block_reg[1][109]/U3  ( .A(\block[1][109] ), .B(block_next[109]), 
        .S0(n1598), .Y(n671) );
  DFFQXL \block_reg[1][109]  ( .D(n671), .CK(clk), .Q(\block[1][109] ) );
  CLKMX2X2 \block_reg[1][108]/U3  ( .A(\block[1][108] ), .B(block_next[108]), 
        .S0(n1598), .Y(n670) );
  DFFQXL \block_reg[1][108]  ( .D(n670), .CK(clk), .Q(\block[1][108] ) );
  CLKMX2X2 \block_reg[1][107]/U3  ( .A(\block[1][107] ), .B(block_next[107]), 
        .S0(n1598), .Y(n669) );
  DFFQXL \block_reg[1][107]  ( .D(n669), .CK(clk), .Q(\block[1][107] ) );
  CLKMX2X2 \block_reg[1][105]/U3  ( .A(\block[1][105] ), .B(block_next[105]), 
        .S0(n1598), .Y(n668) );
  DFFQXL \block_reg[1][105]  ( .D(n668), .CK(clk), .Q(\block[1][105] ) );
  DFFQXL \block_reg[0][118]  ( .D(n667), .CK(clk), .Q(\block[0][118] ) );
  DFFQXL \block_reg[0][117]  ( .D(n666), .CK(clk), .Q(\block[0][117] ) );
  DFFQXL \block_reg[0][116]  ( .D(n665), .CK(clk), .Q(\block[0][116] ) );
  CLKMX2X2 \block_reg[0][115]/U3  ( .A(\block[0][115] ), .B(block_next[115]), 
        .S0(n1613), .Y(n664) );
  DFFQXL \block_reg[0][115]  ( .D(n664), .CK(clk), .Q(\block[0][115] ) );
  CLKMX2X2 \block_reg[0][114]/U3  ( .A(\block[0][114] ), .B(block_next[114]), 
        .S0(n1613), .Y(n663) );
  DFFQXL \block_reg[0][114]  ( .D(n663), .CK(clk), .Q(\block[0][114] ) );
  CLKMX2X2 \block_reg[0][113]/U3  ( .A(\block[0][113] ), .B(block_next[113]), 
        .S0(n1613), .Y(n662) );
  DFFQXL \block_reg[0][113]  ( .D(n662), .CK(clk), .Q(\block[0][113] ) );
  CLKMX2X2 \block_reg[0][112]/U3  ( .A(\block[0][112] ), .B(block_next[112]), 
        .S0(n1613), .Y(n661) );
  DFFQXL \block_reg[0][112]  ( .D(n661), .CK(clk), .Q(\block[0][112] ) );
  CLKMX2X2 \block_reg[0][111]/U3  ( .A(\block[0][111] ), .B(block_next[111]), 
        .S0(n1613), .Y(n660) );
  DFFQXL \block_reg[0][111]  ( .D(n660), .CK(clk), .Q(\block[0][111] ) );
  CLKMX2X2 \block_reg[0][110]/U3  ( .A(\block[0][110] ), .B(block_next[110]), 
        .S0(n1613), .Y(n659) );
  DFFQXL \block_reg[0][110]  ( .D(n659), .CK(clk), .Q(\block[0][110] ) );
  CLKMX2X2 \block_reg[0][109]/U3  ( .A(\block[0][109] ), .B(block_next[109]), 
        .S0(n1613), .Y(n658) );
  DFFQXL \block_reg[0][109]  ( .D(n658), .CK(clk), .Q(\block[0][109] ) );
  CLKMX2X2 \block_reg[0][108]/U3  ( .A(\block[0][108] ), .B(block_next[108]), 
        .S0(n1613), .Y(n657) );
  DFFQXL \block_reg[0][108]  ( .D(n657), .CK(clk), .Q(\block[0][108] ) );
  CLKMX2X2 \block_reg[0][107]/U3  ( .A(\block[0][107] ), .B(block_next[107]), 
        .S0(n1613), .Y(n656) );
  DFFQXL \block_reg[0][107]  ( .D(n656), .CK(clk), .Q(\block[0][107] ) );
  DFFQXL \block_reg[0][105]  ( .D(n655), .CK(clk), .Q(\block[0][105] ) );
  CLKMX2X2 \block_reg[7][9]/U3  ( .A(\block[7][9] ), .B(block_next[9]), .S0(
        n1498), .Y(n654) );
  DFFQXL \block_reg[7][9]  ( .D(n654), .CK(clk), .Q(\block[7][9] ) );
  CLKMX2X2 \block_reg[7][8]/U3  ( .A(\block[7][8] ), .B(block_next[8]), .S0(
        n1498), .Y(n653) );
  DFFQXL \block_reg[7][8]  ( .D(n653), .CK(clk), .Q(\block[7][8] ) );
  CLKMX2X2 \block_reg[6][9]/U3  ( .A(\block[6][9] ), .B(block_next[9]), .S0(
        n1513), .Y(n652) );
  DFFQXL \block_reg[6][9]  ( .D(n652), .CK(clk), .Q(\block[6][9] ) );
  CLKMX2X2 \block_reg[6][8]/U3  ( .A(\block[6][8] ), .B(block_next[8]), .S0(
        n1513), .Y(n651) );
  DFFQXL \block_reg[6][8]  ( .D(n651), .CK(clk), .Q(\block[6][8] ) );
  CLKMX2X2 \block_reg[5][9]/U3  ( .A(\block[5][9] ), .B(block_next[9]), .S0(
        n1529), .Y(n650) );
  DFFQXL \block_reg[5][9]  ( .D(n650), .CK(clk), .Q(\block[5][9] ) );
  CLKMX2X2 \block_reg[5][8]/U3  ( .A(\block[5][8] ), .B(block_next[8]), .S0(
        n1529), .Y(n649) );
  DFFQXL \block_reg[5][8]  ( .D(n649), .CK(clk), .Q(\block[5][8] ) );
  CLKMX2X2 \block_reg[4][9]/U3  ( .A(\block[4][9] ), .B(block_next[9]), .S0(
        n1546), .Y(n648) );
  DFFQXL \block_reg[4][9]  ( .D(n648), .CK(clk), .Q(\block[4][9] ) );
  CLKMX2X2 \block_reg[4][8]/U3  ( .A(\block[4][8] ), .B(block_next[8]), .S0(
        n1546), .Y(n647) );
  DFFQXL \block_reg[4][8]  ( .D(n647), .CK(clk), .Q(\block[4][8] ) );
  CLKMX2X2 \block_reg[3][9]/U3  ( .A(\block[3][9] ), .B(block_next[9]), .S0(
        n1563), .Y(n646) );
  DFFQXL \block_reg[3][9]  ( .D(n646), .CK(clk), .Q(\block[3][9] ) );
  CLKMX2X2 \block_reg[3][8]/U3  ( .A(\block[3][8] ), .B(block_next[8]), .S0(
        n1563), .Y(n645) );
  DFFQXL \block_reg[3][8]  ( .D(n645), .CK(clk), .Q(\block[3][8] ) );
  CLKMX2X2 \block_reg[2][9]/U3  ( .A(\block[2][9] ), .B(block_next[9]), .S0(
        n1576), .Y(n644) );
  DFFQXL \block_reg[2][9]  ( .D(n644), .CK(clk), .Q(\block[2][9] ) );
  CLKMX2X2 \block_reg[2][8]/U3  ( .A(\block[2][8] ), .B(block_next[8]), .S0(
        n1576), .Y(n643) );
  DFFQXL \block_reg[2][8]  ( .D(n643), .CK(clk), .Q(\block[2][8] ) );
  CLKMX2X2 \block_reg[1][9]/U3  ( .A(\block[1][9] ), .B(block_next[9]), .S0(
        n1590), .Y(n642) );
  DFFQXL \block_reg[1][9]  ( .D(n642), .CK(clk), .Q(\block[1][9] ) );
  CLKMX2X2 \block_reg[1][8]/U3  ( .A(\block[1][8] ), .B(block_next[8]), .S0(
        n1590), .Y(n641) );
  DFFQXL \block_reg[1][8]  ( .D(n641), .CK(clk), .Q(\block[1][8] ) );
  CLKMX2X2 \block_reg[0][9]/U3  ( .A(\block[0][9] ), .B(block_next[9]), .S0(
        n1605), .Y(n640) );
  DFFQXL \block_reg[0][9]  ( .D(n640), .CK(clk), .Q(\block[0][9] ) );
  CLKMX2X2 \block_reg[0][8]/U3  ( .A(\block[0][8] ), .B(block_next[8]), .S0(
        n1605), .Y(n639) );
  DFFQXL \block_reg[0][8]  ( .D(n639), .CK(clk), .Q(\block[0][8] ) );
  CLKMX2X2 \block_reg[7][39]/U3  ( .A(\block[7][39] ), .B(block_next[39]), 
        .S0(n1500), .Y(n638) );
  DFFQXL \block_reg[7][39]  ( .D(n638), .CK(clk), .Q(\block[7][39] ) );
  DFFQXL \block_reg[7][38]  ( .D(n637), .CK(clk), .Q(\block[7][38] ) );
  CLKMX2X2 \block_reg[7][37]/U3  ( .A(\block[7][37] ), .B(block_next[37]), 
        .S0(n1500), .Y(n636) );
  DFFQXL \block_reg[7][37]  ( .D(n636), .CK(clk), .Q(\block[7][37] ) );
  CLKMX2X2 \block_reg[7][36]/U3  ( .A(\block[7][36] ), .B(block_next[36]), 
        .S0(n1500), .Y(n635) );
  DFFQXL \block_reg[7][36]  ( .D(n635), .CK(clk), .Q(\block[7][36] ) );
  CLKMX2X2 \block_reg[7][35]/U3  ( .A(\block[7][35] ), .B(block_next[35]), 
        .S0(n1500), .Y(n634) );
  DFFQXL \block_reg[7][35]  ( .D(n634), .CK(clk), .Q(\block[7][35] ) );
  CLKMX2X2 \block_reg[7][34]/U3  ( .A(\block[7][34] ), .B(block_next[34]), 
        .S0(n1500), .Y(n633) );
  DFFQXL \block_reg[7][34]  ( .D(n633), .CK(clk), .Q(\block[7][34] ) );
  CLKMX2X2 \block_reg[7][33]/U3  ( .A(\block[7][33] ), .B(block_next[33]), 
        .S0(n1500), .Y(n632) );
  DFFQXL \block_reg[7][33]  ( .D(n632), .CK(clk), .Q(\block[7][33] ) );
  CLKMX2X2 \block_reg[7][32]/U3  ( .A(\block[7][32] ), .B(block_next[32]), 
        .S0(n1500), .Y(n631) );
  DFFQXL \block_reg[7][32]  ( .D(n631), .CK(clk), .Q(\block[7][32] ) );
  CLKMX2X2 \block_reg[6][39]/U3  ( .A(\block[6][39] ), .B(block_next[39]), 
        .S0(n1515), .Y(n630) );
  DFFQXL \block_reg[6][39]  ( .D(n630), .CK(clk), .Q(\block[6][39] ) );
  DFFQXL \block_reg[6][38]  ( .D(n629), .CK(clk), .Q(\block[6][38] ) );
  CLKMX2X2 \block_reg[6][37]/U3  ( .A(\block[6][37] ), .B(block_next[37]), 
        .S0(n1515), .Y(n628) );
  DFFQXL \block_reg[6][37]  ( .D(n628), .CK(clk), .Q(\block[6][37] ) );
  CLKMX2X2 \block_reg[6][36]/U3  ( .A(\block[6][36] ), .B(block_next[36]), 
        .S0(n1515), .Y(n627) );
  DFFQXL \block_reg[6][36]  ( .D(n627), .CK(clk), .Q(\block[6][36] ) );
  CLKMX2X2 \block_reg[6][35]/U3  ( .A(\block[6][35] ), .B(block_next[35]), 
        .S0(n1515), .Y(n626) );
  DFFQXL \block_reg[6][35]  ( .D(n626), .CK(clk), .Q(\block[6][35] ) );
  CLKMX2X2 \block_reg[6][34]/U3  ( .A(\block[6][34] ), .B(block_next[34]), 
        .S0(n1515), .Y(n625) );
  DFFQXL \block_reg[6][34]  ( .D(n625), .CK(clk), .Q(\block[6][34] ) );
  CLKMX2X2 \block_reg[6][33]/U3  ( .A(\block[6][33] ), .B(block_next[33]), 
        .S0(n1515), .Y(n624) );
  DFFQXL \block_reg[6][33]  ( .D(n624), .CK(clk), .Q(\block[6][33] ) );
  CLKMX2X2 \block_reg[6][32]/U3  ( .A(\block[6][32] ), .B(block_next[32]), 
        .S0(n1515), .Y(n623) );
  DFFQXL \block_reg[6][32]  ( .D(n623), .CK(clk), .Q(\block[6][32] ) );
  CLKMX2X2 \block_reg[5][39]/U3  ( .A(\block[5][39] ), .B(block_next[39]), 
        .S0(n1531), .Y(n622) );
  DFFQXL \block_reg[5][39]  ( .D(n622), .CK(clk), .Q(\block[5][39] ) );
  DFFQXL \block_reg[5][38]  ( .D(n621), .CK(clk), .Q(\block[5][38] ) );
  CLKMX2X2 \block_reg[5][37]/U3  ( .A(\block[5][37] ), .B(block_next[37]), 
        .S0(n1531), .Y(n620) );
  DFFQXL \block_reg[5][37]  ( .D(n620), .CK(clk), .Q(\block[5][37] ) );
  CLKMX2X2 \block_reg[5][36]/U3  ( .A(\block[5][36] ), .B(block_next[36]), 
        .S0(n1531), .Y(n619) );
  DFFQXL \block_reg[5][36]  ( .D(n619), .CK(clk), .Q(\block[5][36] ) );
  CLKMX2X2 \block_reg[5][35]/U3  ( .A(\block[5][35] ), .B(block_next[35]), 
        .S0(n1531), .Y(n618) );
  DFFQXL \block_reg[5][35]  ( .D(n618), .CK(clk), .Q(\block[5][35] ) );
  CLKMX2X2 \block_reg[5][34]/U3  ( .A(\block[5][34] ), .B(block_next[34]), 
        .S0(n1531), .Y(n617) );
  DFFQXL \block_reg[5][34]  ( .D(n617), .CK(clk), .Q(\block[5][34] ) );
  CLKMX2X2 \block_reg[5][33]/U3  ( .A(\block[5][33] ), .B(block_next[33]), 
        .S0(n1531), .Y(n616) );
  DFFQXL \block_reg[5][33]  ( .D(n616), .CK(clk), .Q(\block[5][33] ) );
  CLKMX2X2 \block_reg[5][32]/U3  ( .A(\block[5][32] ), .B(block_next[32]), 
        .S0(n1531), .Y(n615) );
  DFFQXL \block_reg[5][32]  ( .D(n615), .CK(clk), .Q(\block[5][32] ) );
  CLKMX2X2 \block_reg[4][39]/U3  ( .A(\block[4][39] ), .B(block_next[39]), 
        .S0(n1548), .Y(n614) );
  DFFQXL \block_reg[4][39]  ( .D(n614), .CK(clk), .Q(\block[4][39] ) );
  DFFQXL \block_reg[4][38]  ( .D(n613), .CK(clk), .Q(\block[4][38] ) );
  CLKMX2X2 \block_reg[4][37]/U3  ( .A(\block[4][37] ), .B(block_next[37]), 
        .S0(n1548), .Y(n612) );
  DFFQXL \block_reg[4][37]  ( .D(n612), .CK(clk), .Q(\block[4][37] ) );
  CLKMX2X2 \block_reg[4][36]/U3  ( .A(\block[4][36] ), .B(block_next[36]), 
        .S0(n1548), .Y(n611) );
  DFFQXL \block_reg[4][36]  ( .D(n611), .CK(clk), .Q(\block[4][36] ) );
  CLKMX2X2 \block_reg[4][35]/U3  ( .A(\block[4][35] ), .B(block_next[35]), 
        .S0(n1548), .Y(n610) );
  DFFQXL \block_reg[4][35]  ( .D(n610), .CK(clk), .Q(\block[4][35] ) );
  CLKMX2X2 \block_reg[4][34]/U3  ( .A(\block[4][34] ), .B(block_next[34]), 
        .S0(n1548), .Y(n609) );
  DFFQXL \block_reg[4][34]  ( .D(n609), .CK(clk), .Q(\block[4][34] ) );
  CLKMX2X2 \block_reg[4][33]/U3  ( .A(\block[4][33] ), .B(block_next[33]), 
        .S0(n1548), .Y(n608) );
  DFFQXL \block_reg[4][33]  ( .D(n608), .CK(clk), .Q(\block[4][33] ) );
  CLKMX2X2 \block_reg[4][32]/U3  ( .A(\block[4][32] ), .B(block_next[32]), 
        .S0(n1548), .Y(n607) );
  DFFQXL \block_reg[4][32]  ( .D(n607), .CK(clk), .Q(\block[4][32] ) );
  CLKMX2X2 \block_reg[3][39]/U3  ( .A(\block[3][39] ), .B(block_next[39]), 
        .S0(n1565), .Y(n606) );
  DFFQXL \block_reg[3][39]  ( .D(n606), .CK(clk), .Q(\block[3][39] ) );
  DFFQXL \block_reg[3][38]  ( .D(n605), .CK(clk), .Q(\block[3][38] ) );
  CLKMX2X2 \block_reg[3][37]/U3  ( .A(\block[3][37] ), .B(block_next[37]), 
        .S0(n1565), .Y(n604) );
  DFFQXL \block_reg[3][37]  ( .D(n604), .CK(clk), .Q(\block[3][37] ) );
  CLKMX2X2 \block_reg[3][36]/U3  ( .A(\block[3][36] ), .B(block_next[36]), 
        .S0(n1565), .Y(n603) );
  DFFQXL \block_reg[3][36]  ( .D(n603), .CK(clk), .Q(\block[3][36] ) );
  CLKMX2X2 \block_reg[3][35]/U3  ( .A(\block[3][35] ), .B(block_next[35]), 
        .S0(n1565), .Y(n602) );
  DFFQXL \block_reg[3][35]  ( .D(n602), .CK(clk), .Q(\block[3][35] ) );
  CLKMX2X2 \block_reg[3][34]/U3  ( .A(\block[3][34] ), .B(block_next[34]), 
        .S0(n1565), .Y(n601) );
  DFFQXL \block_reg[3][34]  ( .D(n601), .CK(clk), .Q(\block[3][34] ) );
  CLKMX2X2 \block_reg[3][33]/U3  ( .A(\block[3][33] ), .B(block_next[33]), 
        .S0(n1565), .Y(n600) );
  DFFQXL \block_reg[3][33]  ( .D(n600), .CK(clk), .Q(\block[3][33] ) );
  CLKMX2X2 \block_reg[3][32]/U3  ( .A(\block[3][32] ), .B(block_next[32]), 
        .S0(n1565), .Y(n599) );
  DFFQXL \block_reg[3][32]  ( .D(n599), .CK(clk), .Q(\block[3][32] ) );
  CLKMX2X2 \block_reg[2][39]/U3  ( .A(\block[2][39] ), .B(block_next[39]), 
        .S0(n1578), .Y(n598) );
  DFFQXL \block_reg[2][39]  ( .D(n598), .CK(clk), .Q(\block[2][39] ) );
  DFFQXL \block_reg[2][38]  ( .D(n597), .CK(clk), .Q(\block[2][38] ) );
  CLKMX2X2 \block_reg[2][37]/U3  ( .A(\block[2][37] ), .B(block_next[37]), 
        .S0(n1578), .Y(n596) );
  DFFQXL \block_reg[2][37]  ( .D(n596), .CK(clk), .Q(\block[2][37] ) );
  CLKMX2X2 \block_reg[2][36]/U3  ( .A(\block[2][36] ), .B(block_next[36]), 
        .S0(n1578), .Y(n595) );
  DFFQXL \block_reg[2][36]  ( .D(n595), .CK(clk), .Q(\block[2][36] ) );
  CLKMX2X2 \block_reg[2][35]/U3  ( .A(\block[2][35] ), .B(block_next[35]), 
        .S0(n1578), .Y(n594) );
  DFFQXL \block_reg[2][35]  ( .D(n594), .CK(clk), .Q(\block[2][35] ) );
  CLKMX2X2 \block_reg[2][34]/U3  ( .A(\block[2][34] ), .B(block_next[34]), 
        .S0(n1578), .Y(n593) );
  DFFQXL \block_reg[2][34]  ( .D(n593), .CK(clk), .Q(\block[2][34] ) );
  CLKMX2X2 \block_reg[2][33]/U3  ( .A(\block[2][33] ), .B(block_next[33]), 
        .S0(n1578), .Y(n592) );
  DFFQXL \block_reg[2][33]  ( .D(n592), .CK(clk), .Q(\block[2][33] ) );
  CLKMX2X2 \block_reg[2][32]/U3  ( .A(\block[2][32] ), .B(block_next[32]), 
        .S0(n1578), .Y(n591) );
  DFFQXL \block_reg[2][32]  ( .D(n591), .CK(clk), .Q(\block[2][32] ) );
  CLKMX2X2 \block_reg[1][39]/U3  ( .A(\block[1][39] ), .B(block_next[39]), 
        .S0(n1592), .Y(n590) );
  DFFQXL \block_reg[1][39]  ( .D(n590), .CK(clk), .Q(\block[1][39] ) );
  DFFQXL \block_reg[1][38]  ( .D(n589), .CK(clk), .Q(\block[1][38] ) );
  CLKMX2X2 \block_reg[1][37]/U3  ( .A(\block[1][37] ), .B(block_next[37]), 
        .S0(n1592), .Y(n588) );
  DFFQXL \block_reg[1][37]  ( .D(n588), .CK(clk), .Q(\block[1][37] ) );
  CLKMX2X2 \block_reg[1][36]/U3  ( .A(\block[1][36] ), .B(block_next[36]), 
        .S0(n1592), .Y(n587) );
  DFFQXL \block_reg[1][36]  ( .D(n587), .CK(clk), .Q(\block[1][36] ) );
  CLKMX2X2 \block_reg[1][35]/U3  ( .A(\block[1][35] ), .B(block_next[35]), 
        .S0(n1592), .Y(n586) );
  DFFQXL \block_reg[1][35]  ( .D(n586), .CK(clk), .Q(\block[1][35] ) );
  CLKMX2X2 \block_reg[1][34]/U3  ( .A(\block[1][34] ), .B(block_next[34]), 
        .S0(n1592), .Y(n585) );
  DFFQXL \block_reg[1][34]  ( .D(n585), .CK(clk), .Q(\block[1][34] ) );
  CLKMX2X2 \block_reg[1][33]/U3  ( .A(\block[1][33] ), .B(block_next[33]), 
        .S0(n1592), .Y(n584) );
  DFFQXL \block_reg[1][33]  ( .D(n584), .CK(clk), .Q(\block[1][33] ) );
  CLKMX2X2 \block_reg[1][32]/U3  ( .A(\block[1][32] ), .B(block_next[32]), 
        .S0(n1592), .Y(n583) );
  DFFQXL \block_reg[1][32]  ( .D(n583), .CK(clk), .Q(\block[1][32] ) );
  CLKMX2X2 \block_reg[0][39]/U3  ( .A(\block[0][39] ), .B(block_next[39]), 
        .S0(n1607), .Y(n582) );
  DFFQXL \block_reg[0][39]  ( .D(n582), .CK(clk), .Q(\block[0][39] ) );
  CLKMX2X2 \block_reg[0][37]/U3  ( .A(\block[0][37] ), .B(block_next[37]), 
        .S0(n1607), .Y(n580) );
  DFFQXL \block_reg[0][37]  ( .D(n580), .CK(clk), .Q(\block[0][37] ) );
  CLKMX2X2 \block_reg[0][36]/U3  ( .A(\block[0][36] ), .B(block_next[36]), 
        .S0(n1607), .Y(n579) );
  DFFQXL \block_reg[0][36]  ( .D(n579), .CK(clk), .Q(\block[0][36] ) );
  CLKMX2X2 \block_reg[0][35]/U3  ( .A(\block[0][35] ), .B(block_next[35]), 
        .S0(n1607), .Y(n578) );
  DFFQXL \block_reg[0][35]  ( .D(n578), .CK(clk), .Q(\block[0][35] ) );
  CLKMX2X2 \block_reg[0][34]/U3  ( .A(\block[0][34] ), .B(block_next[34]), 
        .S0(n1607), .Y(n577) );
  DFFQXL \block_reg[0][34]  ( .D(n577), .CK(clk), .Q(\block[0][34] ) );
  CLKMX2X2 \block_reg[0][33]/U3  ( .A(\block[0][33] ), .B(block_next[33]), 
        .S0(n1607), .Y(n576) );
  DFFQXL \block_reg[0][33]  ( .D(n576), .CK(clk), .Q(\block[0][33] ) );
  CLKMX2X2 \block_reg[0][32]/U3  ( .A(\block[0][32] ), .B(block_next[32]), 
        .S0(n1607), .Y(n575) );
  DFFQXL \block_reg[0][32]  ( .D(n575), .CK(clk), .Q(\block[0][32] ) );
  CLKMX2X2 \block_reg[7][7]/U3  ( .A(\block[7][7] ), .B(n38), .S0(n1498), .Y(
        n574) );
  DFFQXL \block_reg[7][7]  ( .D(n574), .CK(clk), .Q(\block[7][7] ) );
  CLKMX2X2 \block_reg[7][6]/U3  ( .A(\block[7][6] ), .B(block_next[6]), .S0(
        n1498), .Y(n573) );
  DFFQXL \block_reg[7][6]  ( .D(n573), .CK(clk), .Q(\block[7][6] ) );
  CLKMX2X2 \block_reg[7][5]/U3  ( .A(\block[7][5] ), .B(block_next[5]), .S0(
        n1498), .Y(n572) );
  DFFQXL \block_reg[7][5]  ( .D(n572), .CK(clk), .Q(\block[7][5] ) );
  CLKMX2X2 \block_reg[7][4]/U3  ( .A(\block[7][4] ), .B(block_next[4]), .S0(
        n1498), .Y(n571) );
  DFFQXL \block_reg[7][4]  ( .D(n571), .CK(clk), .Q(\block[7][4] ) );
  CLKMX2X2 \block_reg[7][3]/U3  ( .A(\block[7][3] ), .B(block_next[3]), .S0(
        n1498), .Y(n570) );
  DFFQXL \block_reg[7][3]  ( .D(n570), .CK(clk), .Q(\block[7][3] ) );
  CLKMX2X2 \block_reg[7][2]/U3  ( .A(\block[7][2] ), .B(block_next[2]), .S0(
        n1498), .Y(n569) );
  DFFQXL \block_reg[7][2]  ( .D(n569), .CK(clk), .Q(\block[7][2] ) );
  CLKMX2X2 \block_reg[7][1]/U3  ( .A(\block[7][1] ), .B(n47), .S0(n1498), .Y(
        n568) );
  DFFQXL \block_reg[7][1]  ( .D(n568), .CK(clk), .Q(\block[7][1] ) );
  CLKMX2X2 \block_reg[7][0]/U3  ( .A(\block[7][0] ), .B(block_next[0]), .S0(
        n1497), .Y(n567) );
  DFFQXL \block_reg[7][0]  ( .D(n567), .CK(clk), .Q(\block[7][0] ) );
  CLKMX2X2 \block_reg[6][7]/U3  ( .A(\block[6][7] ), .B(n38), .S0(n1513), .Y(
        n566) );
  DFFQXL \block_reg[6][7]  ( .D(n566), .CK(clk), .Q(\block[6][7] ) );
  CLKMX2X2 \block_reg[6][6]/U3  ( .A(\block[6][6] ), .B(block_next[6]), .S0(
        n1513), .Y(n565) );
  DFFQXL \block_reg[6][6]  ( .D(n565), .CK(clk), .Q(\block[6][6] ) );
  CLKMX2X2 \block_reg[6][5]/U3  ( .A(\block[6][5] ), .B(block_next[5]), .S0(
        n1513), .Y(n564) );
  DFFQXL \block_reg[6][5]  ( .D(n564), .CK(clk), .Q(\block[6][5] ) );
  CLKMX2X2 \block_reg[6][4]/U3  ( .A(\block[6][4] ), .B(block_next[4]), .S0(
        n1513), .Y(n563) );
  DFFQXL \block_reg[6][4]  ( .D(n563), .CK(clk), .Q(\block[6][4] ) );
  CLKMX2X2 \block_reg[6][3]/U3  ( .A(\block[6][3] ), .B(block_next[3]), .S0(
        n1513), .Y(n562) );
  DFFQXL \block_reg[6][3]  ( .D(n562), .CK(clk), .Q(\block[6][3] ) );
  CLKMX2X2 \block_reg[6][2]/U3  ( .A(\block[6][2] ), .B(block_next[2]), .S0(
        n1513), .Y(n561) );
  DFFQXL \block_reg[6][2]  ( .D(n561), .CK(clk), .Q(\block[6][2] ) );
  CLKMX2X2 \block_reg[6][1]/U3  ( .A(\block[6][1] ), .B(n47), .S0(n1513), .Y(
        n560) );
  DFFQXL \block_reg[6][1]  ( .D(n560), .CK(clk), .Q(\block[6][1] ) );
  CLKMX2X2 \block_reg[6][0]/U3  ( .A(\block[6][0] ), .B(block_next[0]), .S0(
        n1512), .Y(n559) );
  DFFQXL \block_reg[6][0]  ( .D(n559), .CK(clk), .Q(\block[6][0] ) );
  CLKMX2X2 \block_reg[5][7]/U3  ( .A(\block[5][7] ), .B(n38), .S0(n1529), .Y(
        n558) );
  DFFQXL \block_reg[5][7]  ( .D(n558), .CK(clk), .Q(\block[5][7] ) );
  DFFQXL \block_reg[5][6]  ( .D(n557), .CK(clk), .Q(\block[5][6] ) );
  DFFQXL \block_reg[5][5]  ( .D(n556), .CK(clk), .Q(\block[5][5] ) );
  DFFQXL \block_reg[5][4]  ( .D(n555), .CK(clk), .Q(\block[5][4] ) );
  DFFQXL \block_reg[5][3]  ( .D(n554), .CK(clk), .Q(\block[5][3] ) );
  CLKMX2X2 \block_reg[5][2]/U3  ( .A(\block[5][2] ), .B(block_next[2]), .S0(
        n1529), .Y(n553) );
  DFFQXL \block_reg[5][2]  ( .D(n553), .CK(clk), .Q(\block[5][2] ) );
  CLKMX2X2 \block_reg[5][1]/U3  ( .A(\block[5][1] ), .B(n47), .S0(n1529), .Y(
        n552) );
  DFFQXL \block_reg[5][1]  ( .D(n552), .CK(clk), .Q(\block[5][1] ) );
  CLKMX2X2 \block_reg[5][0]/U3  ( .A(\block[5][0] ), .B(block_next[0]), .S0(
        n1528), .Y(n551) );
  DFFQXL \block_reg[5][0]  ( .D(n551), .CK(clk), .Q(\block[5][0] ) );
  CLKMX2X2 \block_reg[4][7]/U3  ( .A(\block[4][7] ), .B(n38), .S0(n1546), .Y(
        n550) );
  DFFQXL \block_reg[4][7]  ( .D(n550), .CK(clk), .Q(\block[4][7] ) );
  DFFQXL \block_reg[4][6]  ( .D(n549), .CK(clk), .Q(\block[4][6] ) );
  DFFQXL \block_reg[4][5]  ( .D(n548), .CK(clk), .Q(\block[4][5] ) );
  DFFQXL \block_reg[4][4]  ( .D(n547), .CK(clk), .Q(\block[4][4] ) );
  DFFQXL \block_reg[4][3]  ( .D(n546), .CK(clk), .Q(\block[4][3] ) );
  CLKMX2X2 \block_reg[4][2]/U3  ( .A(\block[4][2] ), .B(block_next[2]), .S0(
        n1546), .Y(n545) );
  DFFQXL \block_reg[4][2]  ( .D(n545), .CK(clk), .Q(\block[4][2] ) );
  CLKMX2X2 \block_reg[4][1]/U3  ( .A(\block[4][1] ), .B(n47), .S0(n1546), .Y(
        n544) );
  DFFQXL \block_reg[4][1]  ( .D(n544), .CK(clk), .Q(\block[4][1] ) );
  CLKMX2X2 \block_reg[4][0]/U3  ( .A(\block[4][0] ), .B(block_next[0]), .S0(
        n1545), .Y(n543) );
  DFFQXL \block_reg[4][0]  ( .D(n543), .CK(clk), .Q(\block[4][0] ) );
  CLKMX2X2 \block_reg[3][7]/U3  ( .A(\block[3][7] ), .B(n38), .S0(n1563), .Y(
        n542) );
  DFFQXL \block_reg[3][7]  ( .D(n542), .CK(clk), .Q(\block[3][7] ) );
  DFFQXL \block_reg[3][6]  ( .D(n541), .CK(clk), .Q(\block[3][6] ) );
  DFFQXL \block_reg[3][5]  ( .D(n540), .CK(clk), .Q(\block[3][5] ) );
  DFFQXL \block_reg[3][4]  ( .D(n539), .CK(clk), .Q(\block[3][4] ) );
  DFFQXL \block_reg[3][3]  ( .D(n538), .CK(clk), .Q(\block[3][3] ) );
  CLKMX2X2 \block_reg[3][2]/U3  ( .A(\block[3][2] ), .B(block_next[2]), .S0(
        n1563), .Y(n537) );
  DFFQXL \block_reg[3][2]  ( .D(n537), .CK(clk), .Q(\block[3][2] ) );
  CLKMX2X2 \block_reg[3][1]/U3  ( .A(\block[3][1] ), .B(n47), .S0(n1563), .Y(
        n536) );
  DFFQXL \block_reg[3][1]  ( .D(n536), .CK(clk), .Q(\block[3][1] ) );
  CLKMX2X2 \block_reg[3][0]/U3  ( .A(\block[3][0] ), .B(block_next[0]), .S0(
        n1562), .Y(n535) );
  DFFQXL \block_reg[3][0]  ( .D(n535), .CK(clk), .Q(\block[3][0] ) );
  CLKMX2X2 \block_reg[2][7]/U3  ( .A(\block[2][7] ), .B(n38), .S0(n1576), .Y(
        n534) );
  DFFQXL \block_reg[2][7]  ( .D(n534), .CK(clk), .Q(\block[2][7] ) );
  DFFQXL \block_reg[2][6]  ( .D(n533), .CK(clk), .Q(\block[2][6] ) );
  DFFQXL \block_reg[2][5]  ( .D(n532), .CK(clk), .Q(\block[2][5] ) );
  DFFQXL \block_reg[2][4]  ( .D(n531), .CK(clk), .Q(\block[2][4] ) );
  DFFQXL \block_reg[2][3]  ( .D(n530), .CK(clk), .Q(\block[2][3] ) );
  CLKMX2X2 \block_reg[2][2]/U3  ( .A(\block[2][2] ), .B(block_next[2]), .S0(
        n1576), .Y(n529) );
  DFFQXL \block_reg[2][2]  ( .D(n529), .CK(clk), .Q(\block[2][2] ) );
  CLKMX2X2 \block_reg[2][1]/U3  ( .A(\block[2][1] ), .B(n47), .S0(n1576), .Y(
        n528) );
  DFFQXL \block_reg[2][1]  ( .D(n528), .CK(clk), .Q(\block[2][1] ) );
  DFFQXL \block_reg[2][0]  ( .D(n527), .CK(clk), .Q(\block[2][0] ) );
  CLKMX2X2 \block_reg[1][7]/U3  ( .A(\block[1][7] ), .B(n38), .S0(n1590), .Y(
        n526) );
  DFFQXL \block_reg[1][7]  ( .D(n526), .CK(clk), .Q(\block[1][7] ) );
  DFFQXL \block_reg[1][6]  ( .D(n525), .CK(clk), .Q(\block[1][6] ) );
  DFFQXL \block_reg[1][5]  ( .D(n524), .CK(clk), .Q(\block[1][5] ) );
  DFFQXL \block_reg[1][4]  ( .D(n523), .CK(clk), .Q(\block[1][4] ) );
  DFFQXL \block_reg[1][3]  ( .D(n522), .CK(clk), .Q(\block[1][3] ) );
  CLKMX2X2 \block_reg[1][2]/U3  ( .A(\block[1][2] ), .B(block_next[2]), .S0(
        n1590), .Y(n521) );
  DFFQXL \block_reg[1][2]  ( .D(n521), .CK(clk), .Q(\block[1][2] ) );
  CLKMX2X2 \block_reg[1][1]/U3  ( .A(\block[1][1] ), .B(n47), .S0(n1590), .Y(
        n520) );
  DFFQXL \block_reg[1][1]  ( .D(n520), .CK(clk), .Q(\block[1][1] ) );
  DFFQXL \block_reg[1][0]  ( .D(n519), .CK(clk), .Q(\block[1][0] ) );
  CLKMX2X2 \block_reg[0][7]/U3  ( .A(\block[0][7] ), .B(n38), .S0(n1605), .Y(
        n518) );
  DFFQXL \block_reg[0][7]  ( .D(n518), .CK(clk), .Q(\block[0][7] ) );
  DFFQXL \block_reg[0][6]  ( .D(n517), .CK(clk), .Q(\block[0][6] ) );
  DFFQXL \block_reg[0][5]  ( .D(n516), .CK(clk), .Q(\block[0][5] ) );
  DFFQXL \block_reg[0][4]  ( .D(n515), .CK(clk), .Q(\block[0][4] ) );
  DFFQXL \block_reg[0][3]  ( .D(n514), .CK(clk), .Q(\block[0][3] ) );
  CLKMX2X2 \block_reg[0][2]/U3  ( .A(\block[0][2] ), .B(block_next[2]), .S0(
        n1605), .Y(n513) );
  DFFQXL \block_reg[0][2]  ( .D(n513), .CK(clk), .Q(\block[0][2] ) );
  CLKMX2X2 \block_reg[0][1]/U3  ( .A(\block[0][1] ), .B(n47), .S0(n1605), .Y(
        n512) );
  DFFQXL \block_reg[0][1]  ( .D(n512), .CK(clk), .Q(\block[0][1] ) );
  CLKMX2X2 \block_reg[7][19]/U3  ( .A(\block[7][19] ), .B(n49), .S0(n1499), 
        .Y(n510) );
  DFFQXL \block_reg[7][19]  ( .D(n510), .CK(clk), .Q(\block[7][19] ) );
  DFFQXL \block_reg[7][18]  ( .D(n509), .CK(clk), .Q(\block[7][18] ) );
  CLKMX2X2 \block_reg[7][17]/U3  ( .A(\block[7][17] ), .B(block_next[17]), 
        .S0(n1499), .Y(n508) );
  DFFQXL \block_reg[7][17]  ( .D(n508), .CK(clk), .Q(\block[7][17] ) );
  CLKMX2X2 \block_reg[7][16]/U3  ( .A(\block[7][16] ), .B(n42), .S0(n1499), 
        .Y(n507) );
  DFFQXL \block_reg[7][16]  ( .D(n507), .CK(clk), .Q(\block[7][16] ) );
  CLKMX2X2 \block_reg[7][15]/U3  ( .A(\block[7][15] ), .B(block_next[15]), 
        .S0(n1499), .Y(n506) );
  DFFQXL \block_reg[7][15]  ( .D(n506), .CK(clk), .Q(\block[7][15] ) );
  CLKMX2X2 \block_reg[7][14]/U3  ( .A(\block[7][14] ), .B(n44), .S0(n1499), 
        .Y(n505) );
  DFFQXL \block_reg[7][14]  ( .D(n505), .CK(clk), .Q(\block[7][14] ) );
  CLKMX2X2 \block_reg[7][13]/U3  ( .A(\block[7][13] ), .B(block_next[13]), 
        .S0(n1498), .Y(n504) );
  DFFQXL \block_reg[7][13]  ( .D(n504), .CK(clk), .Q(\block[7][13] ) );
  CLKMX2X2 \block_reg[7][12]/U3  ( .A(\block[7][12] ), .B(n46), .S0(n1498), 
        .Y(n502) );
  DFFQXL \block_reg[7][12]  ( .D(n502), .CK(clk), .Q(\block[7][12] ) );
  CLKMX2X2 \block_reg[7][11]/U3  ( .A(\block[7][11] ), .B(block_next[11]), 
        .S0(n1498), .Y(n470) );
  DFFQXL \block_reg[7][11]  ( .D(n470), .CK(clk), .Q(\block[7][11] ) );
  CLKMX2X2 \block_reg[7][10]/U3  ( .A(\block[7][10] ), .B(n48), .S0(n1498), 
        .Y(n469) );
  DFFQXL \block_reg[7][10]  ( .D(n469), .CK(clk), .Q(\block[7][10] ) );
  CLKMX2X2 \block_reg[6][19]/U3  ( .A(\block[6][19] ), .B(n49), .S0(n1514), 
        .Y(n468) );
  DFFQXL \block_reg[6][19]  ( .D(n468), .CK(clk), .Q(\block[6][19] ) );
  CLKMX2X2 \block_reg[6][18]/U3  ( .A(\block[6][18] ), .B(n35), .S0(n1514), 
        .Y(n467) );
  DFFQXL \block_reg[6][18]  ( .D(n467), .CK(clk), .Q(\block[6][18] ) );
  CLKMX2X2 \block_reg[6][17]/U3  ( .A(\block[6][17] ), .B(block_next[17]), 
        .S0(n1514), .Y(n466) );
  DFFQXL \block_reg[6][17]  ( .D(n466), .CK(clk), .Q(\block[6][17] ) );
  CLKMX2X2 \block_reg[6][16]/U3  ( .A(\block[6][16] ), .B(n42), .S0(n1514), 
        .Y(n465) );
  DFFQXL \block_reg[6][16]  ( .D(n465), .CK(clk), .Q(\block[6][16] ) );
  CLKMX2X2 \block_reg[6][15]/U3  ( .A(\block[6][15] ), .B(block_next[15]), 
        .S0(n1514), .Y(n464) );
  DFFQXL \block_reg[6][15]  ( .D(n464), .CK(clk), .Q(\block[6][15] ) );
  CLKMX2X2 \block_reg[6][14]/U3  ( .A(\block[6][14] ), .B(n44), .S0(n1514), 
        .Y(n463) );
  DFFQXL \block_reg[6][14]  ( .D(n463), .CK(clk), .Q(\block[6][14] ) );
  CLKMX2X2 \block_reg[6][13]/U3  ( .A(\block[6][13] ), .B(block_next[13]), 
        .S0(n1513), .Y(n462) );
  DFFQXL \block_reg[6][13]  ( .D(n462), .CK(clk), .Q(\block[6][13] ) );
  CLKMX2X2 \block_reg[6][12]/U3  ( .A(\block[6][12] ), .B(n46), .S0(n1513), 
        .Y(n461) );
  DFFQXL \block_reg[6][12]  ( .D(n461), .CK(clk), .Q(\block[6][12] ) );
  CLKMX2X2 \block_reg[6][11]/U3  ( .A(\block[6][11] ), .B(block_next[11]), 
        .S0(n1513), .Y(n460) );
  DFFQXL \block_reg[6][11]  ( .D(n460), .CK(clk), .Q(\block[6][11] ) );
  CLKMX2X2 \block_reg[6][10]/U3  ( .A(\block[6][10] ), .B(n48), .S0(n1513), 
        .Y(n459) );
  DFFQXL \block_reg[6][10]  ( .D(n459), .CK(clk), .Q(\block[6][10] ) );
  CLKMX2X2 \block_reg[5][19]/U3  ( .A(\block[5][19] ), .B(n49), .S0(n1530), 
        .Y(n458) );
  DFFQXL \block_reg[5][19]  ( .D(n458), .CK(clk), .Q(\block[5][19] ) );
  CLKMX2X2 \block_reg[5][18]/U3  ( .A(\block[5][18] ), .B(n35), .S0(n1530), 
        .Y(n457) );
  DFFQXL \block_reg[5][18]  ( .D(n457), .CK(clk), .Q(\block[5][18] ) );
  CLKMX2X2 \block_reg[5][17]/U3  ( .A(\block[5][17] ), .B(block_next[17]), 
        .S0(n1530), .Y(n456) );
  DFFQXL \block_reg[5][17]  ( .D(n456), .CK(clk), .Q(\block[5][17] ) );
  CLKMX2X2 \block_reg[5][16]/U3  ( .A(\block[5][16] ), .B(n42), .S0(n1530), 
        .Y(n455) );
  DFFQXL \block_reg[5][16]  ( .D(n455), .CK(clk), .Q(\block[5][16] ) );
  CLKMX2X2 \block_reg[5][15]/U3  ( .A(\block[5][15] ), .B(block_next[15]), 
        .S0(n1530), .Y(n454) );
  DFFQXL \block_reg[5][15]  ( .D(n454), .CK(clk), .Q(\block[5][15] ) );
  CLKMX2X2 \block_reg[5][14]/U3  ( .A(\block[5][14] ), .B(n44), .S0(n1530), 
        .Y(n453) );
  DFFQXL \block_reg[5][14]  ( .D(n453), .CK(clk), .Q(\block[5][14] ) );
  DFFQXL \block_reg[5][13]  ( .D(n452), .CK(clk), .Q(\block[5][13] ) );
  CLKMX2X2 \block_reg[5][12]/U3  ( .A(\block[5][12] ), .B(n46), .S0(n1529), 
        .Y(n451) );
  DFFQXL \block_reg[5][12]  ( .D(n451), .CK(clk), .Q(\block[5][12] ) );
  DFFQXL \block_reg[5][11]  ( .D(n450), .CK(clk), .Q(\block[5][11] ) );
  CLKMX2X2 \block_reg[5][10]/U3  ( .A(\block[5][10] ), .B(n48), .S0(n1529), 
        .Y(n449) );
  DFFQXL \block_reg[5][10]  ( .D(n449), .CK(clk), .Q(\block[5][10] ) );
  CLKMX2X2 \block_reg[4][19]/U3  ( .A(\block[4][19] ), .B(n49), .S0(n1547), 
        .Y(n448) );
  DFFQXL \block_reg[4][19]  ( .D(n448), .CK(clk), .Q(\block[4][19] ) );
  CLKMX2X2 \block_reg[4][18]/U3  ( .A(\block[4][18] ), .B(n35), .S0(n1547), 
        .Y(n447) );
  DFFQXL \block_reg[4][18]  ( .D(n447), .CK(clk), .Q(\block[4][18] ) );
  CLKMX2X2 \block_reg[4][17]/U3  ( .A(\block[4][17] ), .B(block_next[17]), 
        .S0(n1547), .Y(n446) );
  DFFQXL \block_reg[4][17]  ( .D(n446), .CK(clk), .Q(\block[4][17] ) );
  CLKMX2X2 \block_reg[4][16]/U3  ( .A(\block[4][16] ), .B(n42), .S0(n1547), 
        .Y(n445) );
  DFFQXL \block_reg[4][16]  ( .D(n445), .CK(clk), .Q(\block[4][16] ) );
  CLKMX2X2 \block_reg[4][15]/U3  ( .A(\block[4][15] ), .B(block_next[15]), 
        .S0(n1547), .Y(n444) );
  DFFQXL \block_reg[4][15]  ( .D(n444), .CK(clk), .Q(\block[4][15] ) );
  CLKMX2X2 \block_reg[4][14]/U3  ( .A(\block[4][14] ), .B(n44), .S0(n1547), 
        .Y(n443) );
  DFFQXL \block_reg[4][14]  ( .D(n443), .CK(clk), .Q(\block[4][14] ) );
  DFFQXL \block_reg[4][13]  ( .D(n442), .CK(clk), .Q(\block[4][13] ) );
  CLKMX2X2 \block_reg[4][12]/U3  ( .A(\block[4][12] ), .B(n46), .S0(n1546), 
        .Y(n441) );
  DFFQXL \block_reg[4][12]  ( .D(n441), .CK(clk), .Q(\block[4][12] ) );
  DFFQXL \block_reg[4][11]  ( .D(n440), .CK(clk), .Q(\block[4][11] ) );
  CLKMX2X2 \block_reg[4][10]/U3  ( .A(\block[4][10] ), .B(n48), .S0(n1546), 
        .Y(n439) );
  DFFQXL \block_reg[4][10]  ( .D(n439), .CK(clk), .Q(\block[4][10] ) );
  CLKMX2X2 \block_reg[3][19]/U3  ( .A(\block[3][19] ), .B(n49), .S0(n1564), 
        .Y(n438) );
  DFFQXL \block_reg[3][19]  ( .D(n438), .CK(clk), .Q(\block[3][19] ) );
  CLKMX2X2 \block_reg[3][18]/U3  ( .A(\block[3][18] ), .B(n35), .S0(n1564), 
        .Y(n437) );
  DFFQXL \block_reg[3][18]  ( .D(n437), .CK(clk), .Q(\block[3][18] ) );
  CLKMX2X2 \block_reg[3][17]/U3  ( .A(\block[3][17] ), .B(block_next[17]), 
        .S0(n1564), .Y(n436) );
  DFFQXL \block_reg[3][17]  ( .D(n436), .CK(clk), .Q(\block[3][17] ) );
  CLKMX2X2 \block_reg[3][16]/U3  ( .A(\block[3][16] ), .B(n42), .S0(n1564), 
        .Y(n435) );
  DFFQXL \block_reg[3][16]  ( .D(n435), .CK(clk), .Q(\block[3][16] ) );
  CLKMX2X2 \block_reg[3][15]/U3  ( .A(\block[3][15] ), .B(block_next[15]), 
        .S0(n1564), .Y(n434) );
  DFFQXL \block_reg[3][15]  ( .D(n434), .CK(clk), .Q(\block[3][15] ) );
  CLKMX2X2 \block_reg[3][14]/U3  ( .A(\block[3][14] ), .B(n44), .S0(n1564), 
        .Y(n433) );
  DFFQXL \block_reg[3][14]  ( .D(n433), .CK(clk), .Q(\block[3][14] ) );
  DFFQXL \block_reg[3][13]  ( .D(n432), .CK(clk), .Q(\block[3][13] ) );
  CLKMX2X2 \block_reg[3][12]/U3  ( .A(\block[3][12] ), .B(n46), .S0(n1563), 
        .Y(n431) );
  DFFQXL \block_reg[3][12]  ( .D(n431), .CK(clk), .Q(\block[3][12] ) );
  DFFQXL \block_reg[3][11]  ( .D(n430), .CK(clk), .Q(\block[3][11] ) );
  CLKMX2X2 \block_reg[3][10]/U3  ( .A(\block[3][10] ), .B(n48), .S0(n1563), 
        .Y(n429) );
  DFFQXL \block_reg[3][10]  ( .D(n429), .CK(clk), .Q(\block[3][10] ) );
  CLKMX2X2 \block_reg[2][19]/U3  ( .A(\block[2][19] ), .B(n49), .S0(n1577), 
        .Y(n428) );
  DFFQXL \block_reg[2][19]  ( .D(n428), .CK(clk), .Q(\block[2][19] ) );
  CLKMX2X2 \block_reg[2][18]/U3  ( .A(\block[2][18] ), .B(n35), .S0(n1577), 
        .Y(n427) );
  DFFQXL \block_reg[2][18]  ( .D(n427), .CK(clk), .Q(\block[2][18] ) );
  CLKMX2X2 \block_reg[2][17]/U3  ( .A(\block[2][17] ), .B(block_next[17]), 
        .S0(n1577), .Y(n426) );
  DFFQXL \block_reg[2][17]  ( .D(n426), .CK(clk), .Q(\block[2][17] ) );
  CLKMX2X2 \block_reg[2][16]/U3  ( .A(\block[2][16] ), .B(n42), .S0(n1577), 
        .Y(n425) );
  DFFQXL \block_reg[2][16]  ( .D(n425), .CK(clk), .Q(\block[2][16] ) );
  CLKMX2X2 \block_reg[2][15]/U3  ( .A(\block[2][15] ), .B(block_next[15]), 
        .S0(n1577), .Y(n424) );
  DFFQXL \block_reg[2][15]  ( .D(n424), .CK(clk), .Q(\block[2][15] ) );
  CLKMX2X2 \block_reg[2][14]/U3  ( .A(\block[2][14] ), .B(n44), .S0(n1577), 
        .Y(n423) );
  DFFQXL \block_reg[2][14]  ( .D(n423), .CK(clk), .Q(\block[2][14] ) );
  DFFQXL \block_reg[2][13]  ( .D(n422), .CK(clk), .Q(\block[2][13] ) );
  CLKMX2X2 \block_reg[2][12]/U3  ( .A(\block[2][12] ), .B(n46), .S0(n1576), 
        .Y(n421) );
  DFFQXL \block_reg[2][12]  ( .D(n421), .CK(clk), .Q(\block[2][12] ) );
  DFFQXL \block_reg[2][11]  ( .D(n420), .CK(clk), .Q(\block[2][11] ) );
  CLKMX2X2 \block_reg[2][10]/U3  ( .A(\block[2][10] ), .B(n48), .S0(n1576), 
        .Y(n419) );
  DFFQXL \block_reg[2][10]  ( .D(n419), .CK(clk), .Q(\block[2][10] ) );
  CLKMX2X2 \block_reg[1][19]/U3  ( .A(\block[1][19] ), .B(n49), .S0(n1591), 
        .Y(n418) );
  DFFQXL \block_reg[1][19]  ( .D(n418), .CK(clk), .Q(\block[1][19] ) );
  CLKMX2X2 \block_reg[1][17]/U3  ( .A(\block[1][17] ), .B(block_next[17]), 
        .S0(n1591), .Y(n417) );
  DFFQXL \block_reg[1][17]  ( .D(n417), .CK(clk), .Q(\block[1][17] ) );
  CLKMX2X2 \block_reg[1][16]/U3  ( .A(\block[1][16] ), .B(n42), .S0(n1591), 
        .Y(n416) );
  DFFQXL \block_reg[1][16]  ( .D(n416), .CK(clk), .Q(\block[1][16] ) );
  CLKMX2X2 \block_reg[1][15]/U3  ( .A(\block[1][15] ), .B(block_next[15]), 
        .S0(n1591), .Y(n415) );
  DFFQXL \block_reg[1][15]  ( .D(n415), .CK(clk), .Q(\block[1][15] ) );
  CLKMX2X2 \block_reg[1][14]/U3  ( .A(\block[1][14] ), .B(n44), .S0(n1591), 
        .Y(n414) );
  DFFQXL \block_reg[1][14]  ( .D(n414), .CK(clk), .Q(\block[1][14] ) );
  DFFQXL \block_reg[1][13]  ( .D(n413), .CK(clk), .Q(\block[1][13] ) );
  CLKMX2X2 \block_reg[1][12]/U3  ( .A(\block[1][12] ), .B(n46), .S0(n1590), 
        .Y(n412) );
  DFFQXL \block_reg[1][12]  ( .D(n412), .CK(clk), .Q(\block[1][12] ) );
  DFFQXL \block_reg[1][11]  ( .D(n411), .CK(clk), .Q(\block[1][11] ) );
  CLKMX2X2 \block_reg[1][10]/U3  ( .A(\block[1][10] ), .B(n48), .S0(n1590), 
        .Y(n410) );
  DFFQXL \block_reg[1][10]  ( .D(n410), .CK(clk), .Q(\block[1][10] ) );
  CLKMX2X2 \block_reg[0][19]/U3  ( .A(\block[0][19] ), .B(n49), .S0(n1606), 
        .Y(n409) );
  DFFQXL \block_reg[0][19]  ( .D(n409), .CK(clk), .Q(\block[0][19] ) );
  CLKMX2X2 \block_reg[0][17]/U3  ( .A(\block[0][17] ), .B(block_next[17]), 
        .S0(n1606), .Y(n408) );
  DFFQXL \block_reg[0][17]  ( .D(n408), .CK(clk), .Q(\block[0][17] ) );
  CLKMX2X2 \block_reg[0][16]/U3  ( .A(\block[0][16] ), .B(n42), .S0(n1606), 
        .Y(n407) );
  DFFQXL \block_reg[0][16]  ( .D(n407), .CK(clk), .Q(\block[0][16] ) );
  CLKMX2X2 \block_reg[0][15]/U3  ( .A(\block[0][15] ), .B(block_next[15]), 
        .S0(n1606), .Y(n406) );
  DFFQXL \block_reg[0][15]  ( .D(n406), .CK(clk), .Q(\block[0][15] ) );
  CLKMX2X2 \block_reg[0][14]/U3  ( .A(\block[0][14] ), .B(n44), .S0(n1606), 
        .Y(n405) );
  DFFQXL \block_reg[0][14]  ( .D(n405), .CK(clk), .Q(\block[0][14] ) );
  DFFQXL \block_reg[0][13]  ( .D(n404), .CK(clk), .Q(\block[0][13] ) );
  CLKMX2X2 \block_reg[0][12]/U3  ( .A(\block[0][12] ), .B(n46), .S0(n1605), 
        .Y(n403) );
  DFFQXL \block_reg[0][12]  ( .D(n403), .CK(clk), .Q(\block[0][12] ) );
  DFFQXL \block_reg[0][11]  ( .D(n402), .CK(clk), .Q(\block[0][11] ) );
  CLKMX2X2 \block_reg[0][10]/U3  ( .A(\block[0][10] ), .B(n48), .S0(n1605), 
        .Y(n401) );
  DFFQXL \block_reg[0][10]  ( .D(n401), .CK(clk), .Q(\block[0][10] ) );
  CLKMX2X2 \block_reg[7][63]/U3  ( .A(\block[7][63] ), .B(block_next[63]), 
        .S0(n1502), .Y(n400) );
  DFFQXL \block_reg[7][63]  ( .D(n400), .CK(clk), .Q(\block[7][63] ) );
  CLKMX2X2 \block_reg[7][62]/U3  ( .A(\block[7][62] ), .B(block_next[62]), 
        .S0(n1502), .Y(n399) );
  DFFQXL \block_reg[7][62]  ( .D(n399), .CK(clk), .Q(\block[7][62] ) );
  CLKMX2X2 \block_reg[7][61]/U3  ( .A(\block[7][61] ), .B(block_next[61]), 
        .S0(n1502), .Y(n398) );
  DFFQXL \block_reg[7][61]  ( .D(n398), .CK(clk), .Q(\block[7][61] ) );
  CLKMX2X2 \block_reg[7][60]/U3  ( .A(\block[7][60] ), .B(block_next[60]), 
        .S0(n1502), .Y(n397) );
  DFFQXL \block_reg[7][60]  ( .D(n397), .CK(clk), .Q(\block[7][60] ) );
  CLKMX2X2 \block_reg[7][59]/U3  ( .A(\block[7][59] ), .B(block_next[59]), 
        .S0(n1502), .Y(n396) );
  DFFQXL \block_reg[7][59]  ( .D(n396), .CK(clk), .Q(\block[7][59] ) );
  CLKMX2X2 \block_reg[7][58]/U3  ( .A(\block[7][58] ), .B(block_next[58]), 
        .S0(n1502), .Y(n395) );
  DFFQXL \block_reg[7][58]  ( .D(n395), .CK(clk), .Q(\block[7][58] ) );
  CLKMX2X2 \block_reg[7][57]/U3  ( .A(\block[7][57] ), .B(block_next[57]), 
        .S0(n1502), .Y(n394) );
  DFFQXL \block_reg[7][57]  ( .D(n394), .CK(clk), .Q(\block[7][57] ) );
  CLKMX2X2 \block_reg[7][56]/U3  ( .A(\block[7][56] ), .B(block_next[56]), 
        .S0(n1502), .Y(n393) );
  DFFQXL \block_reg[7][56]  ( .D(n393), .CK(clk), .Q(\block[7][56] ) );
  CLKMX2X2 \block_reg[7][54]/U3  ( .A(\block[7][54] ), .B(block_next[54]), 
        .S0(n1502), .Y(n392) );
  DFFQXL \block_reg[7][54]  ( .D(n392), .CK(clk), .Q(\block[7][54] ) );
  CLKMX2X2 \block_reg[7][53]/U3  ( .A(\block[7][53] ), .B(block_next[53]), 
        .S0(n1502), .Y(n391) );
  DFFQXL \block_reg[7][53]  ( .D(n391), .CK(clk), .Q(\block[7][53] ) );
  CLKMX2X2 \block_reg[7][52]/U3  ( .A(\block[7][52] ), .B(block_next[52]), 
        .S0(n1501), .Y(n390) );
  DFFQXL \block_reg[7][52]  ( .D(n390), .CK(clk), .Q(\block[7][52] ) );
  DFFQXL \block_reg[7][51]  ( .D(n389), .CK(clk), .Q(\block[7][51] ) );
  CLKMX2X2 \block_reg[7][50]/U3  ( .A(\block[7][50] ), .B(block_next[50]), 
        .S0(n1501), .Y(n388) );
  DFFQXL \block_reg[7][50]  ( .D(n388), .CK(clk), .Q(\block[7][50] ) );
  CLKMX2X2 \block_reg[7][49]/U3  ( .A(\block[7][49] ), .B(block_next[49]), 
        .S0(n1501), .Y(n387) );
  DFFQXL \block_reg[7][49]  ( .D(n387), .CK(clk), .Q(\block[7][49] ) );
  CLKMX2X2 \block_reg[7][48]/U3  ( .A(\block[7][48] ), .B(block_next[48]), 
        .S0(n1501), .Y(n386) );
  DFFQXL \block_reg[7][48]  ( .D(n386), .CK(clk), .Q(\block[7][48] ) );
  CLKMX2X2 \block_reg[7][47]/U3  ( .A(\block[7][47] ), .B(block_next[47]), 
        .S0(n1501), .Y(n385) );
  DFFQXL \block_reg[7][47]  ( .D(n385), .CK(clk), .Q(\block[7][47] ) );
  CLKMX2X2 \block_reg[7][46]/U3  ( .A(\block[7][46] ), .B(block_next[46]), 
        .S0(n1501), .Y(n384) );
  DFFQXL \block_reg[7][46]  ( .D(n384), .CK(clk), .Q(\block[7][46] ) );
  CLKMX2X2 \block_reg[7][45]/U3  ( .A(\block[7][45] ), .B(block_next[45]), 
        .S0(n1501), .Y(n383) );
  DFFQXL \block_reg[7][45]  ( .D(n383), .CK(clk), .Q(\block[7][45] ) );
  CLKMX2X2 \block_reg[7][44]/U3  ( .A(\block[7][44] ), .B(block_next[44]), 
        .S0(n1501), .Y(n382) );
  DFFQXL \block_reg[7][44]  ( .D(n382), .CK(clk), .Q(\block[7][44] ) );
  CLKMX2X2 \block_reg[7][43]/U3  ( .A(\block[7][43] ), .B(block_next[43]), 
        .S0(n1501), .Y(n381) );
  DFFQXL \block_reg[7][43]  ( .D(n381), .CK(clk), .Q(\block[7][43] ) );
  CLKMX2X2 \block_reg[7][42]/U3  ( .A(\block[7][42] ), .B(block_next[42]), 
        .S0(n1501), .Y(n380) );
  DFFQXL \block_reg[7][42]  ( .D(n380), .CK(clk), .Q(\block[7][42] ) );
  CLKMX2X2 \block_reg[7][41]/U3  ( .A(\block[7][41] ), .B(block_next[41]), 
        .S0(n1501), .Y(n379) );
  DFFQXL \block_reg[7][41]  ( .D(n379), .CK(clk), .Q(\block[7][41] ) );
  CLKMX2X2 \block_reg[7][40]/U3  ( .A(\block[7][40] ), .B(n39), .S0(n1501), 
        .Y(n378) );
  DFFQXL \block_reg[7][40]  ( .D(n378), .CK(clk), .Q(\block[7][40] ) );
  CLKMX2X2 \block_reg[6][63]/U3  ( .A(\block[6][63] ), .B(block_next[63]), 
        .S0(n1517), .Y(n377) );
  DFFQXL \block_reg[6][63]  ( .D(n377), .CK(clk), .Q(\block[6][63] ) );
  CLKMX2X2 \block_reg[6][62]/U3  ( .A(\block[6][62] ), .B(block_next[62]), 
        .S0(n1517), .Y(n376) );
  DFFQXL \block_reg[6][62]  ( .D(n376), .CK(clk), .Q(\block[6][62] ) );
  CLKMX2X2 \block_reg[6][61]/U3  ( .A(\block[6][61] ), .B(block_next[61]), 
        .S0(n1517), .Y(n375) );
  DFFQXL \block_reg[6][61]  ( .D(n375), .CK(clk), .Q(\block[6][61] ) );
  CLKMX2X2 \block_reg[6][60]/U3  ( .A(\block[6][60] ), .B(block_next[60]), 
        .S0(n1517), .Y(n374) );
  DFFQXL \block_reg[6][60]  ( .D(n374), .CK(clk), .Q(\block[6][60] ) );
  CLKMX2X2 \block_reg[6][59]/U3  ( .A(\block[6][59] ), .B(block_next[59]), 
        .S0(n1517), .Y(n373) );
  DFFQXL \block_reg[6][59]  ( .D(n373), .CK(clk), .Q(\block[6][59] ) );
  CLKMX2X2 \block_reg[6][58]/U3  ( .A(\block[6][58] ), .B(block_next[58]), 
        .S0(n1517), .Y(n372) );
  DFFQXL \block_reg[6][58]  ( .D(n372), .CK(clk), .Q(\block[6][58] ) );
  CLKMX2X2 \block_reg[6][57]/U3  ( .A(\block[6][57] ), .B(block_next[57]), 
        .S0(n1517), .Y(n371) );
  DFFQXL \block_reg[6][57]  ( .D(n371), .CK(clk), .Q(\block[6][57] ) );
  CLKMX2X2 \block_reg[6][56]/U3  ( .A(\block[6][56] ), .B(block_next[56]), 
        .S0(n1517), .Y(n370) );
  DFFQXL \block_reg[6][56]  ( .D(n370), .CK(clk), .Q(\block[6][56] ) );
  CLKMX2X2 \block_reg[6][54]/U3  ( .A(\block[6][54] ), .B(block_next[54]), 
        .S0(n1517), .Y(n369) );
  DFFQXL \block_reg[6][54]  ( .D(n369), .CK(clk), .Q(\block[6][54] ) );
  CLKMX2X2 \block_reg[6][53]/U3  ( .A(\block[6][53] ), .B(block_next[53]), 
        .S0(n1517), .Y(n368) );
  DFFQXL \block_reg[6][53]  ( .D(n368), .CK(clk), .Q(\block[6][53] ) );
  CLKMX2X2 \block_reg[6][52]/U3  ( .A(\block[6][52] ), .B(block_next[52]), 
        .S0(n1516), .Y(n367) );
  DFFQXL \block_reg[6][52]  ( .D(n367), .CK(clk), .Q(\block[6][52] ) );
  DFFQXL \block_reg[6][51]  ( .D(n366), .CK(clk), .Q(\block[6][51] ) );
  CLKMX2X2 \block_reg[6][50]/U3  ( .A(\block[6][50] ), .B(block_next[50]), 
        .S0(n1516), .Y(n365) );
  DFFQXL \block_reg[6][50]  ( .D(n365), .CK(clk), .Q(\block[6][50] ) );
  CLKMX2X2 \block_reg[6][49]/U3  ( .A(\block[6][49] ), .B(block_next[49]), 
        .S0(n1516), .Y(n364) );
  DFFQXL \block_reg[6][49]  ( .D(n364), .CK(clk), .Q(\block[6][49] ) );
  CLKMX2X2 \block_reg[6][48]/U3  ( .A(\block[6][48] ), .B(block_next[48]), 
        .S0(n1516), .Y(n363) );
  DFFQXL \block_reg[6][48]  ( .D(n363), .CK(clk), .Q(\block[6][48] ) );
  CLKMX2X2 \block_reg[6][47]/U3  ( .A(\block[6][47] ), .B(block_next[47]), 
        .S0(n1516), .Y(n362) );
  DFFQXL \block_reg[6][47]  ( .D(n362), .CK(clk), .Q(\block[6][47] ) );
  CLKMX2X2 \block_reg[6][46]/U3  ( .A(\block[6][46] ), .B(block_next[46]), 
        .S0(n1516), .Y(n361) );
  DFFQXL \block_reg[6][46]  ( .D(n361), .CK(clk), .Q(\block[6][46] ) );
  CLKMX2X2 \block_reg[6][45]/U3  ( .A(\block[6][45] ), .B(block_next[45]), 
        .S0(n1516), .Y(n360) );
  DFFQXL \block_reg[6][45]  ( .D(n360), .CK(clk), .Q(\block[6][45] ) );
  CLKMX2X2 \block_reg[6][44]/U3  ( .A(\block[6][44] ), .B(block_next[44]), 
        .S0(n1516), .Y(n359) );
  DFFQXL \block_reg[6][44]  ( .D(n359), .CK(clk), .Q(\block[6][44] ) );
  CLKMX2X2 \block_reg[6][43]/U3  ( .A(\block[6][43] ), .B(block_next[43]), 
        .S0(n1516), .Y(n358) );
  DFFQXL \block_reg[6][43]  ( .D(n358), .CK(clk), .Q(\block[6][43] ) );
  CLKMX2X2 \block_reg[6][42]/U3  ( .A(\block[6][42] ), .B(block_next[42]), 
        .S0(n1516), .Y(n357) );
  DFFQXL \block_reg[6][42]  ( .D(n357), .CK(clk), .Q(\block[6][42] ) );
  CLKMX2X2 \block_reg[6][41]/U3  ( .A(\block[6][41] ), .B(block_next[41]), 
        .S0(n1516), .Y(n356) );
  DFFQXL \block_reg[6][41]  ( .D(n356), .CK(clk), .Q(\block[6][41] ) );
  CLKMX2X2 \block_reg[6][40]/U3  ( .A(\block[6][40] ), .B(n39), .S0(n1516), 
        .Y(n355) );
  DFFQXL \block_reg[6][40]  ( .D(n355), .CK(clk), .Q(\block[6][40] ) );
  CLKMX2X2 \block_reg[5][63]/U3  ( .A(\block[5][63] ), .B(block_next[63]), 
        .S0(n1533), .Y(n354) );
  DFFQXL \block_reg[5][63]  ( .D(n354), .CK(clk), .Q(\block[5][63] ) );
  CLKMX2X2 \block_reg[5][62]/U3  ( .A(\block[5][62] ), .B(block_next[62]), 
        .S0(n1533), .Y(n353) );
  DFFQXL \block_reg[5][62]  ( .D(n353), .CK(clk), .Q(\block[5][62] ) );
  CLKMX2X2 \block_reg[5][61]/U3  ( .A(\block[5][61] ), .B(block_next[61]), 
        .S0(n1533), .Y(n352) );
  DFFQXL \block_reg[5][61]  ( .D(n352), .CK(clk), .Q(\block[5][61] ) );
  CLKMX2X2 \block_reg[5][60]/U3  ( .A(\block[5][60] ), .B(block_next[60]), 
        .S0(n1533), .Y(n351) );
  DFFQXL \block_reg[5][60]  ( .D(n351), .CK(clk), .Q(\block[5][60] ) );
  CLKMX2X2 \block_reg[5][59]/U3  ( .A(\block[5][59] ), .B(block_next[59]), 
        .S0(n1533), .Y(n350) );
  DFFQXL \block_reg[5][59]  ( .D(n350), .CK(clk), .Q(\block[5][59] ) );
  CLKMX2X2 \block_reg[5][58]/U3  ( .A(\block[5][58] ), .B(block_next[58]), 
        .S0(n1533), .Y(n349) );
  DFFQXL \block_reg[5][58]  ( .D(n349), .CK(clk), .Q(\block[5][58] ) );
  CLKMX2X2 \block_reg[5][57]/U3  ( .A(\block[5][57] ), .B(block_next[57]), 
        .S0(n1533), .Y(n348) );
  DFFQXL \block_reg[5][57]  ( .D(n348), .CK(clk), .Q(\block[5][57] ) );
  CLKMX2X2 \block_reg[5][56]/U3  ( .A(\block[5][56] ), .B(block_next[56]), 
        .S0(n1533), .Y(n347) );
  DFFQXL \block_reg[5][56]  ( .D(n347), .CK(clk), .Q(\block[5][56] ) );
  CLKMX2X2 \block_reg[5][54]/U3  ( .A(\block[5][54] ), .B(block_next[54]), 
        .S0(n1533), .Y(n346) );
  DFFQXL \block_reg[5][54]  ( .D(n346), .CK(clk), .Q(\block[5][54] ) );
  CLKMX2X2 \block_reg[5][53]/U3  ( .A(\block[5][53] ), .B(block_next[53]), 
        .S0(n1533), .Y(n345) );
  DFFQXL \block_reg[5][53]  ( .D(n345), .CK(clk), .Q(\block[5][53] ) );
  CLKMX2X2 \block_reg[5][52]/U3  ( .A(\block[5][52] ), .B(block_next[52]), 
        .S0(n1532), .Y(n344) );
  DFFQXL \block_reg[5][52]  ( .D(n344), .CK(clk), .Q(\block[5][52] ) );
  DFFQXL \block_reg[5][51]  ( .D(n343), .CK(clk), .Q(\block[5][51] ) );
  CLKMX2X2 \block_reg[5][50]/U3  ( .A(\block[5][50] ), .B(block_next[50]), 
        .S0(n1532), .Y(n342) );
  DFFQXL \block_reg[5][50]  ( .D(n342), .CK(clk), .Q(\block[5][50] ) );
  CLKMX2X2 \block_reg[5][49]/U3  ( .A(\block[5][49] ), .B(block_next[49]), 
        .S0(n1532), .Y(n341) );
  DFFQXL \block_reg[5][49]  ( .D(n341), .CK(clk), .Q(\block[5][49] ) );
  CLKMX2X2 \block_reg[5][48]/U3  ( .A(\block[5][48] ), .B(block_next[48]), 
        .S0(n1532), .Y(n340) );
  DFFQXL \block_reg[5][48]  ( .D(n340), .CK(clk), .Q(\block[5][48] ) );
  CLKMX2X2 \block_reg[5][47]/U3  ( .A(\block[5][47] ), .B(block_next[47]), 
        .S0(n1532), .Y(n339) );
  DFFQXL \block_reg[5][47]  ( .D(n339), .CK(clk), .Q(\block[5][47] ) );
  CLKMX2X2 \block_reg[5][46]/U3  ( .A(\block[5][46] ), .B(block_next[46]), 
        .S0(n1532), .Y(n338) );
  DFFQXL \block_reg[5][46]  ( .D(n338), .CK(clk), .Q(\block[5][46] ) );
  CLKMX2X2 \block_reg[5][45]/U3  ( .A(\block[5][45] ), .B(block_next[45]), 
        .S0(n1532), .Y(n337) );
  DFFQXL \block_reg[5][45]  ( .D(n337), .CK(clk), .Q(\block[5][45] ) );
  CLKMX2X2 \block_reg[5][44]/U3  ( .A(\block[5][44] ), .B(block_next[44]), 
        .S0(n1532), .Y(n336) );
  DFFQXL \block_reg[5][44]  ( .D(n336), .CK(clk), .Q(\block[5][44] ) );
  CLKMX2X2 \block_reg[5][43]/U3  ( .A(\block[5][43] ), .B(block_next[43]), 
        .S0(n1532), .Y(n335) );
  DFFQXL \block_reg[5][43]  ( .D(n335), .CK(clk), .Q(\block[5][43] ) );
  CLKMX2X2 \block_reg[5][42]/U3  ( .A(\block[5][42] ), .B(block_next[42]), 
        .S0(n1532), .Y(n334) );
  DFFQXL \block_reg[5][42]  ( .D(n334), .CK(clk), .Q(\block[5][42] ) );
  CLKMX2X2 \block_reg[5][41]/U3  ( .A(\block[5][41] ), .B(block_next[41]), 
        .S0(n1532), .Y(n333) );
  DFFQXL \block_reg[5][41]  ( .D(n333), .CK(clk), .Q(\block[5][41] ) );
  CLKMX2X2 \block_reg[5][40]/U3  ( .A(\block[5][40] ), .B(n39), .S0(n1532), 
        .Y(n332) );
  DFFQXL \block_reg[5][40]  ( .D(n332), .CK(clk), .Q(\block[5][40] ) );
  CLKMX2X2 \block_reg[4][63]/U3  ( .A(\block[4][63] ), .B(block_next[63]), 
        .S0(n1550), .Y(n331) );
  DFFQXL \block_reg[4][63]  ( .D(n331), .CK(clk), .Q(\block[4][63] ) );
  CLKMX2X2 \block_reg[4][62]/U3  ( .A(\block[4][62] ), .B(block_next[62]), 
        .S0(n1550), .Y(n330) );
  DFFQXL \block_reg[4][62]  ( .D(n330), .CK(clk), .Q(\block[4][62] ) );
  CLKMX2X2 \block_reg[4][61]/U3  ( .A(\block[4][61] ), .B(block_next[61]), 
        .S0(n1550), .Y(n329) );
  DFFQXL \block_reg[4][61]  ( .D(n329), .CK(clk), .Q(\block[4][61] ) );
  CLKMX2X2 \block_reg[4][60]/U3  ( .A(\block[4][60] ), .B(block_next[60]), 
        .S0(n1550), .Y(n328) );
  DFFQXL \block_reg[4][60]  ( .D(n328), .CK(clk), .Q(\block[4][60] ) );
  CLKMX2X2 \block_reg[4][59]/U3  ( .A(\block[4][59] ), .B(block_next[59]), 
        .S0(n1550), .Y(n327) );
  DFFQXL \block_reg[4][59]  ( .D(n327), .CK(clk), .Q(\block[4][59] ) );
  CLKMX2X2 \block_reg[4][58]/U3  ( .A(\block[4][58] ), .B(block_next[58]), 
        .S0(n1550), .Y(n326) );
  DFFQXL \block_reg[4][58]  ( .D(n326), .CK(clk), .Q(\block[4][58] ) );
  CLKMX2X2 \block_reg[4][57]/U3  ( .A(\block[4][57] ), .B(block_next[57]), 
        .S0(n1550), .Y(n325) );
  DFFQXL \block_reg[4][57]  ( .D(n325), .CK(clk), .Q(\block[4][57] ) );
  CLKMX2X2 \block_reg[4][56]/U3  ( .A(\block[4][56] ), .B(block_next[56]), 
        .S0(n1550), .Y(n324) );
  DFFQXL \block_reg[4][56]  ( .D(n324), .CK(clk), .Q(\block[4][56] ) );
  CLKMX2X2 \block_reg[4][54]/U3  ( .A(\block[4][54] ), .B(block_next[54]), 
        .S0(n1550), .Y(n323) );
  DFFQXL \block_reg[4][54]  ( .D(n323), .CK(clk), .Q(\block[4][54] ) );
  CLKMX2X2 \block_reg[4][53]/U3  ( .A(\block[4][53] ), .B(block_next[53]), 
        .S0(n1550), .Y(n322) );
  DFFQXL \block_reg[4][53]  ( .D(n322), .CK(clk), .Q(\block[4][53] ) );
  CLKMX2X2 \block_reg[4][52]/U3  ( .A(\block[4][52] ), .B(block_next[52]), 
        .S0(n1549), .Y(n321) );
  DFFQXL \block_reg[4][52]  ( .D(n321), .CK(clk), .Q(\block[4][52] ) );
  DFFQXL \block_reg[4][51]  ( .D(n320), .CK(clk), .Q(\block[4][51] ) );
  CLKMX2X2 \block_reg[4][50]/U3  ( .A(\block[4][50] ), .B(block_next[50]), 
        .S0(n1549), .Y(n319) );
  DFFQXL \block_reg[4][50]  ( .D(n319), .CK(clk), .Q(\block[4][50] ) );
  CLKMX2X2 \block_reg[4][49]/U3  ( .A(\block[4][49] ), .B(block_next[49]), 
        .S0(n1549), .Y(n318) );
  DFFQXL \block_reg[4][49]  ( .D(n318), .CK(clk), .Q(\block[4][49] ) );
  CLKMX2X2 \block_reg[4][48]/U3  ( .A(\block[4][48] ), .B(block_next[48]), 
        .S0(n1549), .Y(n317) );
  DFFQXL \block_reg[4][48]  ( .D(n317), .CK(clk), .Q(\block[4][48] ) );
  CLKMX2X2 \block_reg[4][47]/U3  ( .A(\block[4][47] ), .B(block_next[47]), 
        .S0(n1549), .Y(n316) );
  DFFQXL \block_reg[4][47]  ( .D(n316), .CK(clk), .Q(\block[4][47] ) );
  CLKMX2X2 \block_reg[4][46]/U3  ( .A(\block[4][46] ), .B(block_next[46]), 
        .S0(n1549), .Y(n315) );
  DFFQXL \block_reg[4][46]  ( .D(n315), .CK(clk), .Q(\block[4][46] ) );
  CLKMX2X2 \block_reg[4][45]/U3  ( .A(\block[4][45] ), .B(block_next[45]), 
        .S0(n1549), .Y(n314) );
  DFFQXL \block_reg[4][45]  ( .D(n314), .CK(clk), .Q(\block[4][45] ) );
  CLKMX2X2 \block_reg[4][44]/U3  ( .A(\block[4][44] ), .B(block_next[44]), 
        .S0(n1549), .Y(n313) );
  DFFQXL \block_reg[4][44]  ( .D(n313), .CK(clk), .Q(\block[4][44] ) );
  CLKMX2X2 \block_reg[4][43]/U3  ( .A(\block[4][43] ), .B(block_next[43]), 
        .S0(n1549), .Y(n312) );
  DFFQXL \block_reg[4][43]  ( .D(n312), .CK(clk), .Q(\block[4][43] ) );
  CLKMX2X2 \block_reg[4][42]/U3  ( .A(\block[4][42] ), .B(block_next[42]), 
        .S0(n1549), .Y(n311) );
  DFFQXL \block_reg[4][42]  ( .D(n311), .CK(clk), .Q(\block[4][42] ) );
  CLKMX2X2 \block_reg[4][41]/U3  ( .A(\block[4][41] ), .B(block_next[41]), 
        .S0(n1549), .Y(n310) );
  DFFQXL \block_reg[4][41]  ( .D(n310), .CK(clk), .Q(\block[4][41] ) );
  CLKMX2X2 \block_reg[4][40]/U3  ( .A(\block[4][40] ), .B(n39), .S0(n1549), 
        .Y(n309) );
  DFFQXL \block_reg[4][40]  ( .D(n309), .CK(clk), .Q(\block[4][40] ) );
  CLKMX2X2 \block_reg[3][63]/U3  ( .A(\block[3][63] ), .B(block_next[63]), 
        .S0(n1567), .Y(n308) );
  DFFQXL \block_reg[3][63]  ( .D(n308), .CK(clk), .Q(\block[3][63] ) );
  CLKMX2X2 \block_reg[3][62]/U3  ( .A(\block[3][62] ), .B(block_next[62]), 
        .S0(n1567), .Y(n307) );
  DFFQXL \block_reg[3][62]  ( .D(n307), .CK(clk), .Q(\block[3][62] ) );
  CLKMX2X2 \block_reg[3][61]/U3  ( .A(\block[3][61] ), .B(block_next[61]), 
        .S0(n1567), .Y(n306) );
  DFFQXL \block_reg[3][61]  ( .D(n306), .CK(clk), .Q(\block[3][61] ) );
  CLKMX2X2 \block_reg[3][60]/U3  ( .A(\block[3][60] ), .B(block_next[60]), 
        .S0(n1567), .Y(n305) );
  DFFQXL \block_reg[3][60]  ( .D(n305), .CK(clk), .Q(\block[3][60] ) );
  CLKMX2X2 \block_reg[3][59]/U3  ( .A(\block[3][59] ), .B(block_next[59]), 
        .S0(n1567), .Y(n304) );
  DFFQXL \block_reg[3][59]  ( .D(n304), .CK(clk), .Q(\block[3][59] ) );
  CLKMX2X2 \block_reg[3][58]/U3  ( .A(\block[3][58] ), .B(block_next[58]), 
        .S0(n1567), .Y(n303) );
  DFFQXL \block_reg[3][58]  ( .D(n303), .CK(clk), .Q(\block[3][58] ) );
  CLKMX2X2 \block_reg[3][57]/U3  ( .A(\block[3][57] ), .B(block_next[57]), 
        .S0(n1567), .Y(n302) );
  DFFQXL \block_reg[3][57]  ( .D(n302), .CK(clk), .Q(\block[3][57] ) );
  CLKMX2X2 \block_reg[3][56]/U3  ( .A(\block[3][56] ), .B(block_next[56]), 
        .S0(n1567), .Y(n301) );
  DFFQXL \block_reg[3][56]  ( .D(n301), .CK(clk), .Q(\block[3][56] ) );
  CLKMX2X2 \block_reg[3][54]/U3  ( .A(\block[3][54] ), .B(block_next[54]), 
        .S0(n1567), .Y(n300) );
  DFFQXL \block_reg[3][54]  ( .D(n300), .CK(clk), .Q(\block[3][54] ) );
  CLKMX2X2 \block_reg[3][53]/U3  ( .A(\block[3][53] ), .B(block_next[53]), 
        .S0(n1567), .Y(n299) );
  DFFQXL \block_reg[3][53]  ( .D(n299), .CK(clk), .Q(\block[3][53] ) );
  CLKMX2X2 \block_reg[3][52]/U3  ( .A(\block[3][52] ), .B(block_next[52]), 
        .S0(n1566), .Y(n298) );
  DFFQXL \block_reg[3][52]  ( .D(n298), .CK(clk), .Q(\block[3][52] ) );
  DFFQXL \block_reg[3][51]  ( .D(n297), .CK(clk), .Q(\block[3][51] ) );
  CLKMX2X2 \block_reg[3][50]/U3  ( .A(\block[3][50] ), .B(block_next[50]), 
        .S0(n1566), .Y(n296) );
  DFFQXL \block_reg[3][50]  ( .D(n296), .CK(clk), .Q(\block[3][50] ) );
  CLKMX2X2 \block_reg[3][49]/U3  ( .A(\block[3][49] ), .B(block_next[49]), 
        .S0(n1566), .Y(n295) );
  DFFQXL \block_reg[3][49]  ( .D(n295), .CK(clk), .Q(\block[3][49] ) );
  CLKMX2X2 \block_reg[3][48]/U3  ( .A(\block[3][48] ), .B(block_next[48]), 
        .S0(n1566), .Y(n294) );
  DFFQXL \block_reg[3][48]  ( .D(n294), .CK(clk), .Q(\block[3][48] ) );
  CLKMX2X2 \block_reg[3][47]/U3  ( .A(\block[3][47] ), .B(block_next[47]), 
        .S0(n1566), .Y(n293) );
  DFFQXL \block_reg[3][47]  ( .D(n293), .CK(clk), .Q(\block[3][47] ) );
  CLKMX2X2 \block_reg[3][46]/U3  ( .A(\block[3][46] ), .B(block_next[46]), 
        .S0(n1566), .Y(n292) );
  DFFQXL \block_reg[3][46]  ( .D(n292), .CK(clk), .Q(\block[3][46] ) );
  CLKMX2X2 \block_reg[3][45]/U3  ( .A(\block[3][45] ), .B(block_next[45]), 
        .S0(n1566), .Y(n291) );
  DFFQXL \block_reg[3][45]  ( .D(n291), .CK(clk), .Q(\block[3][45] ) );
  CLKMX2X2 \block_reg[3][44]/U3  ( .A(\block[3][44] ), .B(block_next[44]), 
        .S0(n1566), .Y(n290) );
  DFFQXL \block_reg[3][44]  ( .D(n290), .CK(clk), .Q(\block[3][44] ) );
  CLKMX2X2 \block_reg[3][43]/U3  ( .A(\block[3][43] ), .B(block_next[43]), 
        .S0(n1566), .Y(n289) );
  DFFQXL \block_reg[3][43]  ( .D(n289), .CK(clk), .Q(\block[3][43] ) );
  CLKMX2X2 \block_reg[3][42]/U3  ( .A(\block[3][42] ), .B(block_next[42]), 
        .S0(n1566), .Y(n288) );
  DFFQXL \block_reg[3][42]  ( .D(n288), .CK(clk), .Q(\block[3][42] ) );
  CLKMX2X2 \block_reg[3][41]/U3  ( .A(\block[3][41] ), .B(block_next[41]), 
        .S0(n1566), .Y(n287) );
  DFFQXL \block_reg[3][41]  ( .D(n287), .CK(clk), .Q(\block[3][41] ) );
  CLKMX2X2 \block_reg[3][40]/U3  ( .A(\block[3][40] ), .B(n39), .S0(n1566), 
        .Y(n286) );
  DFFQXL \block_reg[3][40]  ( .D(n286), .CK(clk), .Q(\block[3][40] ) );
  CLKMX2X2 \block_reg[2][63]/U3  ( .A(\block[2][63] ), .B(block_next[63]), 
        .S0(n1580), .Y(n285) );
  DFFQXL \block_reg[2][63]  ( .D(n285), .CK(clk), .Q(\block[2][63] ) );
  CLKMX2X2 \block_reg[2][62]/U3  ( .A(\block[2][62] ), .B(block_next[62]), 
        .S0(n1580), .Y(n284) );
  DFFQXL \block_reg[2][62]  ( .D(n284), .CK(clk), .Q(\block[2][62] ) );
  CLKMX2X2 \block_reg[2][61]/U3  ( .A(\block[2][61] ), .B(block_next[61]), 
        .S0(n1580), .Y(n283) );
  DFFQXL \block_reg[2][61]  ( .D(n283), .CK(clk), .Q(\block[2][61] ) );
  CLKMX2X2 \block_reg[2][60]/U3  ( .A(\block[2][60] ), .B(block_next[60]), 
        .S0(n1580), .Y(n282) );
  DFFQXL \block_reg[2][60]  ( .D(n282), .CK(clk), .Q(\block[2][60] ) );
  CLKMX2X2 \block_reg[2][59]/U3  ( .A(\block[2][59] ), .B(block_next[59]), 
        .S0(n1580), .Y(n281) );
  DFFQXL \block_reg[2][59]  ( .D(n281), .CK(clk), .Q(\block[2][59] ) );
  CLKMX2X2 \block_reg[2][58]/U3  ( .A(\block[2][58] ), .B(block_next[58]), 
        .S0(n1580), .Y(n280) );
  DFFQXL \block_reg[2][58]  ( .D(n280), .CK(clk), .Q(\block[2][58] ) );
  CLKMX2X2 \block_reg[2][57]/U3  ( .A(\block[2][57] ), .B(block_next[57]), 
        .S0(n1580), .Y(n279) );
  DFFQXL \block_reg[2][57]  ( .D(n279), .CK(clk), .Q(\block[2][57] ) );
  CLKMX2X2 \block_reg[2][56]/U3  ( .A(\block[2][56] ), .B(block_next[56]), 
        .S0(n1580), .Y(n278) );
  DFFQXL \block_reg[2][56]  ( .D(n278), .CK(clk), .Q(\block[2][56] ) );
  CLKMX2X2 \block_reg[2][54]/U3  ( .A(\block[2][54] ), .B(block_next[54]), 
        .S0(n1580), .Y(n277) );
  DFFQXL \block_reg[2][54]  ( .D(n277), .CK(clk), .Q(\block[2][54] ) );
  CLKMX2X2 \block_reg[2][53]/U3  ( .A(\block[2][53] ), .B(block_next[53]), 
        .S0(n1580), .Y(n276) );
  DFFQXL \block_reg[2][53]  ( .D(n276), .CK(clk), .Q(\block[2][53] ) );
  CLKMX2X2 \block_reg[2][52]/U3  ( .A(\block[2][52] ), .B(block_next[52]), 
        .S0(n1579), .Y(n275) );
  DFFQXL \block_reg[2][52]  ( .D(n275), .CK(clk), .Q(\block[2][52] ) );
  DFFQXL \block_reg[2][51]  ( .D(n274), .CK(clk), .Q(\block[2][51] ) );
  CLKMX2X2 \block_reg[2][50]/U3  ( .A(\block[2][50] ), .B(block_next[50]), 
        .S0(n1579), .Y(n273) );
  DFFQXL \block_reg[2][50]  ( .D(n273), .CK(clk), .Q(\block[2][50] ) );
  CLKMX2X2 \block_reg[2][49]/U3  ( .A(\block[2][49] ), .B(block_next[49]), 
        .S0(n1579), .Y(n272) );
  DFFQXL \block_reg[2][49]  ( .D(n272), .CK(clk), .Q(\block[2][49] ) );
  CLKMX2X2 \block_reg[2][48]/U3  ( .A(\block[2][48] ), .B(block_next[48]), 
        .S0(n1579), .Y(n271) );
  DFFQXL \block_reg[2][48]  ( .D(n271), .CK(clk), .Q(\block[2][48] ) );
  CLKMX2X2 \block_reg[2][47]/U3  ( .A(\block[2][47] ), .B(block_next[47]), 
        .S0(n1579), .Y(n270) );
  DFFQXL \block_reg[2][47]  ( .D(n270), .CK(clk), .Q(\block[2][47] ) );
  CLKMX2X2 \block_reg[2][46]/U3  ( .A(\block[2][46] ), .B(block_next[46]), 
        .S0(n1579), .Y(n269) );
  DFFQXL \block_reg[2][46]  ( .D(n269), .CK(clk), .Q(\block[2][46] ) );
  CLKMX2X2 \block_reg[2][45]/U3  ( .A(\block[2][45] ), .B(block_next[45]), 
        .S0(n1579), .Y(n268) );
  DFFQXL \block_reg[2][45]  ( .D(n268), .CK(clk), .Q(\block[2][45] ) );
  CLKMX2X2 \block_reg[2][44]/U3  ( .A(\block[2][44] ), .B(block_next[44]), 
        .S0(n1579), .Y(n267) );
  DFFQXL \block_reg[2][44]  ( .D(n267), .CK(clk), .Q(\block[2][44] ) );
  CLKMX2X2 \block_reg[2][43]/U3  ( .A(\block[2][43] ), .B(block_next[43]), 
        .S0(n1579), .Y(n266) );
  DFFQXL \block_reg[2][43]  ( .D(n266), .CK(clk), .Q(\block[2][43] ) );
  CLKMX2X2 \block_reg[2][42]/U3  ( .A(\block[2][42] ), .B(block_next[42]), 
        .S0(n1579), .Y(n265) );
  DFFQXL \block_reg[2][42]  ( .D(n265), .CK(clk), .Q(\block[2][42] ) );
  CLKMX2X2 \block_reg[2][41]/U3  ( .A(\block[2][41] ), .B(block_next[41]), 
        .S0(n1579), .Y(n264) );
  DFFQXL \block_reg[2][41]  ( .D(n264), .CK(clk), .Q(\block[2][41] ) );
  CLKMX2X2 \block_reg[2][40]/U3  ( .A(\block[2][40] ), .B(n39), .S0(n1579), 
        .Y(n263) );
  DFFQXL \block_reg[2][40]  ( .D(n263), .CK(clk), .Q(\block[2][40] ) );
  CLKMX2X2 \block_reg[1][63]/U3  ( .A(\block[1][63] ), .B(block_next[63]), 
        .S0(n1594), .Y(n262) );
  DFFQXL \block_reg[1][63]  ( .D(n262), .CK(clk), .Q(\block[1][63] ) );
  CLKMX2X2 \block_reg[1][62]/U3  ( .A(\block[1][62] ), .B(block_next[62]), 
        .S0(n1594), .Y(n261) );
  DFFQXL \block_reg[1][62]  ( .D(n261), .CK(clk), .Q(\block[1][62] ) );
  CLKMX2X2 \block_reg[1][61]/U3  ( .A(\block[1][61] ), .B(block_next[61]), 
        .S0(n1594), .Y(n260) );
  DFFQXL \block_reg[1][61]  ( .D(n260), .CK(clk), .Q(\block[1][61] ) );
  CLKMX2X2 \block_reg[1][60]/U3  ( .A(\block[1][60] ), .B(block_next[60]), 
        .S0(n1594), .Y(n259) );
  DFFQXL \block_reg[1][60]  ( .D(n259), .CK(clk), .Q(\block[1][60] ) );
  CLKMX2X2 \block_reg[1][59]/U3  ( .A(\block[1][59] ), .B(block_next[59]), 
        .S0(n1594), .Y(n258) );
  DFFQXL \block_reg[1][59]  ( .D(n258), .CK(clk), .Q(\block[1][59] ) );
  CLKMX2X2 \block_reg[1][58]/U3  ( .A(\block[1][58] ), .B(block_next[58]), 
        .S0(n1594), .Y(n257) );
  DFFQXL \block_reg[1][58]  ( .D(n257), .CK(clk), .Q(\block[1][58] ) );
  CLKMX2X2 \block_reg[1][57]/U3  ( .A(\block[1][57] ), .B(block_next[57]), 
        .S0(n1594), .Y(n256) );
  DFFQXL \block_reg[1][57]  ( .D(n256), .CK(clk), .Q(\block[1][57] ) );
  CLKMX2X2 \block_reg[1][56]/U3  ( .A(\block[1][56] ), .B(block_next[56]), 
        .S0(n1594), .Y(n255) );
  DFFQXL \block_reg[1][56]  ( .D(n255), .CK(clk), .Q(\block[1][56] ) );
  CLKMX2X2 \block_reg[1][54]/U3  ( .A(\block[1][54] ), .B(block_next[54]), 
        .S0(n1594), .Y(n254) );
  DFFQXL \block_reg[1][54]  ( .D(n254), .CK(clk), .Q(\block[1][54] ) );
  CLKMX2X2 \block_reg[1][53]/U3  ( .A(\block[1][53] ), .B(block_next[53]), 
        .S0(n1594), .Y(n253) );
  DFFQXL \block_reg[1][53]  ( .D(n253), .CK(clk), .Q(\block[1][53] ) );
  CLKMX2X2 \block_reg[1][52]/U3  ( .A(\block[1][52] ), .B(block_next[52]), 
        .S0(n1593), .Y(n252) );
  DFFQXL \block_reg[1][52]  ( .D(n252), .CK(clk), .Q(\block[1][52] ) );
  DFFQXL \block_reg[1][51]  ( .D(n251), .CK(clk), .Q(\block[1][51] ) );
  CLKMX2X2 \block_reg[1][50]/U3  ( .A(\block[1][50] ), .B(block_next[50]), 
        .S0(n1593), .Y(n250) );
  DFFQXL \block_reg[1][50]  ( .D(n250), .CK(clk), .Q(\block[1][50] ) );
  CLKMX2X2 \block_reg[1][49]/U3  ( .A(\block[1][49] ), .B(block_next[49]), 
        .S0(n1593), .Y(n249) );
  DFFQXL \block_reg[1][49]  ( .D(n249), .CK(clk), .Q(\block[1][49] ) );
  CLKMX2X2 \block_reg[1][48]/U3  ( .A(\block[1][48] ), .B(block_next[48]), 
        .S0(n1593), .Y(n248) );
  DFFQXL \block_reg[1][48]  ( .D(n248), .CK(clk), .Q(\block[1][48] ) );
  CLKMX2X2 \block_reg[1][47]/U3  ( .A(\block[1][47] ), .B(block_next[47]), 
        .S0(n1593), .Y(n247) );
  DFFQXL \block_reg[1][47]  ( .D(n247), .CK(clk), .Q(\block[1][47] ) );
  CLKMX2X2 \block_reg[1][46]/U3  ( .A(\block[1][46] ), .B(block_next[46]), 
        .S0(n1593), .Y(n246) );
  DFFQXL \block_reg[1][46]  ( .D(n246), .CK(clk), .Q(\block[1][46] ) );
  CLKMX2X2 \block_reg[1][45]/U3  ( .A(\block[1][45] ), .B(block_next[45]), 
        .S0(n1593), .Y(n245) );
  DFFQXL \block_reg[1][45]  ( .D(n245), .CK(clk), .Q(\block[1][45] ) );
  CLKMX2X2 \block_reg[1][44]/U3  ( .A(\block[1][44] ), .B(block_next[44]), 
        .S0(n1593), .Y(n244) );
  DFFQXL \block_reg[1][44]  ( .D(n244), .CK(clk), .Q(\block[1][44] ) );
  CLKMX2X2 \block_reg[1][43]/U3  ( .A(\block[1][43] ), .B(block_next[43]), 
        .S0(n1593), .Y(n243) );
  DFFQXL \block_reg[1][43]  ( .D(n243), .CK(clk), .Q(\block[1][43] ) );
  CLKMX2X2 \block_reg[1][42]/U3  ( .A(\block[1][42] ), .B(block_next[42]), 
        .S0(n1593), .Y(n242) );
  DFFQXL \block_reg[1][42]  ( .D(n242), .CK(clk), .Q(\block[1][42] ) );
  CLKMX2X2 \block_reg[1][41]/U3  ( .A(\block[1][41] ), .B(block_next[41]), 
        .S0(n1593), .Y(n241) );
  DFFQXL \block_reg[1][41]  ( .D(n241), .CK(clk), .Q(\block[1][41] ) );
  CLKMX2X2 \block_reg[1][40]/U3  ( .A(\block[1][40] ), .B(n39), .S0(n1593), 
        .Y(n240) );
  DFFQXL \block_reg[1][40]  ( .D(n240), .CK(clk), .Q(\block[1][40] ) );
  CLKMX2X2 \block_reg[0][63]/U3  ( .A(\block[0][63] ), .B(block_next[63]), 
        .S0(n1609), .Y(n239) );
  DFFQXL \block_reg[0][63]  ( .D(n239), .CK(clk), .Q(\block[0][63] ) );
  CLKMX2X2 \block_reg[0][62]/U3  ( .A(\block[0][62] ), .B(block_next[62]), 
        .S0(n1609), .Y(n238) );
  DFFQXL \block_reg[0][62]  ( .D(n238), .CK(clk), .Q(\block[0][62] ) );
  CLKMX2X2 \block_reg[0][61]/U3  ( .A(\block[0][61] ), .B(block_next[61]), 
        .S0(n1609), .Y(n237) );
  DFFQXL \block_reg[0][61]  ( .D(n237), .CK(clk), .Q(\block[0][61] ) );
  CLKMX2X2 \block_reg[0][60]/U3  ( .A(\block[0][60] ), .B(block_next[60]), 
        .S0(n1609), .Y(n236) );
  DFFQXL \block_reg[0][60]  ( .D(n236), .CK(clk), .Q(\block[0][60] ) );
  CLKMX2X2 \block_reg[0][59]/U3  ( .A(\block[0][59] ), .B(block_next[59]), 
        .S0(n1609), .Y(n235) );
  DFFQXL \block_reg[0][59]  ( .D(n235), .CK(clk), .Q(\block[0][59] ) );
  CLKMX2X2 \block_reg[0][58]/U3  ( .A(\block[0][58] ), .B(block_next[58]), 
        .S0(n1609), .Y(n234) );
  DFFQXL \block_reg[0][58]  ( .D(n234), .CK(clk), .Q(\block[0][58] ) );
  CLKMX2X2 \block_reg[0][57]/U3  ( .A(\block[0][57] ), .B(block_next[57]), 
        .S0(n1609), .Y(n233) );
  DFFQXL \block_reg[0][57]  ( .D(n233), .CK(clk), .Q(\block[0][57] ) );
  CLKMX2X2 \block_reg[0][56]/U3  ( .A(\block[0][56] ), .B(block_next[56]), 
        .S0(n1609), .Y(n232) );
  DFFQXL \block_reg[0][56]  ( .D(n232), .CK(clk), .Q(\block[0][56] ) );
  CLKMX2X2 \block_reg[0][54]/U3  ( .A(\block[0][54] ), .B(block_next[54]), 
        .S0(n1609), .Y(n231) );
  DFFQXL \block_reg[0][54]  ( .D(n231), .CK(clk), .Q(\block[0][54] ) );
  CLKMX2X2 \block_reg[0][53]/U3  ( .A(\block[0][53] ), .B(block_next[53]), 
        .S0(n1609), .Y(n230) );
  DFFQXL \block_reg[0][53]  ( .D(n230), .CK(clk), .Q(\block[0][53] ) );
  CLKMX2X2 \block_reg[0][52]/U3  ( .A(\block[0][52] ), .B(block_next[52]), 
        .S0(n1608), .Y(n229) );
  DFFQXL \block_reg[0][52]  ( .D(n229), .CK(clk), .Q(\block[0][52] ) );
  CLKMX2X2 \block_reg[0][50]/U3  ( .A(\block[0][50] ), .B(block_next[50]), 
        .S0(n1608), .Y(n227) );
  DFFQXL \block_reg[0][50]  ( .D(n227), .CK(clk), .Q(\block[0][50] ) );
  CLKMX2X2 \block_reg[0][49]/U3  ( .A(\block[0][49] ), .B(block_next[49]), 
        .S0(n1608), .Y(n226) );
  DFFQXL \block_reg[0][49]  ( .D(n226), .CK(clk), .Q(\block[0][49] ) );
  CLKMX2X2 \block_reg[0][48]/U3  ( .A(\block[0][48] ), .B(block_next[48]), 
        .S0(n1608), .Y(n225) );
  DFFQXL \block_reg[0][48]  ( .D(n225), .CK(clk), .Q(\block[0][48] ) );
  CLKMX2X2 \block_reg[0][47]/U3  ( .A(\block[0][47] ), .B(block_next[47]), 
        .S0(n1608), .Y(n224) );
  DFFQXL \block_reg[0][47]  ( .D(n224), .CK(clk), .Q(\block[0][47] ) );
  CLKMX2X2 \block_reg[0][46]/U3  ( .A(\block[0][46] ), .B(block_next[46]), 
        .S0(n1608), .Y(n223) );
  DFFQXL \block_reg[0][46]  ( .D(n223), .CK(clk), .Q(\block[0][46] ) );
  CLKMX2X2 \block_reg[0][45]/U3  ( .A(\block[0][45] ), .B(block_next[45]), 
        .S0(n1608), .Y(n222) );
  DFFQXL \block_reg[0][45]  ( .D(n222), .CK(clk), .Q(\block[0][45] ) );
  CLKMX2X2 \block_reg[0][44]/U3  ( .A(\block[0][44] ), .B(block_next[44]), 
        .S0(n1608), .Y(n221) );
  DFFQXL \block_reg[0][44]  ( .D(n221), .CK(clk), .Q(\block[0][44] ) );
  CLKMX2X2 \block_reg[0][43]/U3  ( .A(\block[0][43] ), .B(block_next[43]), 
        .S0(n1608), .Y(n220) );
  DFFQXL \block_reg[0][43]  ( .D(n220), .CK(clk), .Q(\block[0][43] ) );
  CLKMX2X2 \block_reg[0][42]/U3  ( .A(\block[0][42] ), .B(block_next[42]), 
        .S0(n1608), .Y(n219) );
  DFFQXL \block_reg[0][42]  ( .D(n219), .CK(clk), .Q(\block[0][42] ) );
  CLKMX2X2 \block_reg[0][41]/U3  ( .A(\block[0][41] ), .B(block_next[41]), 
        .S0(n1608), .Y(n218) );
  DFFQXL \block_reg[0][41]  ( .D(n218), .CK(clk), .Q(\block[0][41] ) );
  CLKMX2X2 \block_reg[0][40]/U3  ( .A(\block[0][40] ), .B(n39), .S0(n1608), 
        .Y(n217) );
  DFFQXL \block_reg[0][40]  ( .D(n217), .CK(clk), .Q(\block[0][40] ) );
  DFFQXL \block_reg[7][31]  ( .D(n216), .CK(clk), .Q(\block[7][31] ) );
  DFFQXL \block_reg[7][30]  ( .D(n215), .CK(clk), .Q(\block[7][30] ) );
  DFFQXL \block_reg[7][29]  ( .D(n214), .CK(clk), .Q(\block[7][29] ) );
  DFFQXL \block_reg[7][28]  ( .D(n213), .CK(clk), .Q(\block[7][28] ) );
  CLKMX2X2 \block_reg[7][27]/U3  ( .A(\block[7][27] ), .B(block_next[27]), 
        .S0(n1500), .Y(n212) );
  DFFQXL \block_reg[7][27]  ( .D(n212), .CK(clk), .Q(\block[7][27] ) );
  DFFQXL \block_reg[7][26]  ( .D(n211), .CK(clk), .Q(\block[7][26] ) );
  DFFQXL \block_reg[7][25]  ( .D(n210), .CK(clk), .Q(\block[7][25] ) );
  DFFQXL \block_reg[7][24]  ( .D(n209), .CK(clk), .Q(\block[7][24] ) );
  DFFQXL \block_reg[7][23]  ( .D(n208), .CK(clk), .Q(\block[7][23] ) );
  DFFQXL \block_reg[7][22]  ( .D(n207), .CK(clk), .Q(\block[7][22] ) );
  DFFQXL \block_reg[7][21]  ( .D(n206), .CK(clk), .Q(\block[7][21] ) );
  DFFQXL \block_reg[7][20]  ( .D(n205), .CK(clk), .Q(\block[7][20] ) );
  DFFQXL \block_reg[6][31]  ( .D(n204), .CK(clk), .Q(\block[6][31] ) );
  DFFQXL \block_reg[6][30]  ( .D(n203), .CK(clk), .Q(\block[6][30] ) );
  DFFQXL \block_reg[6][29]  ( .D(n202), .CK(clk), .Q(\block[6][29] ) );
  DFFQXL \block_reg[6][28]  ( .D(n201), .CK(clk), .Q(\block[6][28] ) );
  CLKMX2X2 \block_reg[6][27]/U3  ( .A(\block[6][27] ), .B(block_next[27]), 
        .S0(n1515), .Y(n200) );
  DFFQXL \block_reg[6][27]  ( .D(n200), .CK(clk), .Q(\block[6][27] ) );
  DFFQXL \block_reg[6][26]  ( .D(n199), .CK(clk), .Q(\block[6][26] ) );
  DFFQXL \block_reg[6][25]  ( .D(n198), .CK(clk), .Q(\block[6][25] ) );
  DFFQXL \block_reg[6][24]  ( .D(n197), .CK(clk), .Q(\block[6][24] ) );
  DFFQXL \block_reg[6][23]  ( .D(n196), .CK(clk), .Q(\block[6][23] ) );
  DFFQXL \block_reg[6][22]  ( .D(n195), .CK(clk), .Q(\block[6][22] ) );
  DFFQXL \block_reg[6][21]  ( .D(n194), .CK(clk), .Q(\block[6][21] ) );
  DFFQXL \block_reg[6][20]  ( .D(n193), .CK(clk), .Q(\block[6][20] ) );
  DFFQXL \block_reg[5][31]  ( .D(n192), .CK(clk), .Q(\block[5][31] ) );
  DFFQXL \block_reg[5][30]  ( .D(n191), .CK(clk), .Q(\block[5][30] ) );
  DFFQXL \block_reg[5][29]  ( .D(n190), .CK(clk), .Q(\block[5][29] ) );
  DFFQXL \block_reg[5][28]  ( .D(n189), .CK(clk), .Q(\block[5][28] ) );
  CLKMX2X2 \block_reg[5][27]/U3  ( .A(\block[5][27] ), .B(block_next[27]), 
        .S0(n1531), .Y(n188) );
  DFFQXL \block_reg[5][27]  ( .D(n188), .CK(clk), .Q(\block[5][27] ) );
  DFFQXL \block_reg[5][26]  ( .D(n187), .CK(clk), .Q(\block[5][26] ) );
  DFFQXL \block_reg[5][25]  ( .D(n186), .CK(clk), .Q(\block[5][25] ) );
  DFFQXL \block_reg[5][24]  ( .D(n185), .CK(clk), .Q(\block[5][24] ) );
  DFFQXL \block_reg[5][23]  ( .D(n184), .CK(clk), .Q(\block[5][23] ) );
  DFFQXL \block_reg[5][22]  ( .D(n183), .CK(clk), .Q(\block[5][22] ) );
  DFFQXL \block_reg[5][21]  ( .D(n182), .CK(clk), .Q(\block[5][21] ) );
  DFFQXL \block_reg[5][20]  ( .D(n181), .CK(clk), .Q(\block[5][20] ) );
  DFFQXL \block_reg[4][31]  ( .D(n180), .CK(clk), .Q(\block[4][31] ) );
  DFFQXL \block_reg[4][30]  ( .D(n179), .CK(clk), .Q(\block[4][30] ) );
  DFFQXL \block_reg[4][29]  ( .D(n178), .CK(clk), .Q(\block[4][29] ) );
  DFFQXL \block_reg[4][28]  ( .D(n177), .CK(clk), .Q(\block[4][28] ) );
  CLKMX2X2 \block_reg[4][27]/U3  ( .A(\block[4][27] ), .B(block_next[27]), 
        .S0(n1548), .Y(n176) );
  DFFQXL \block_reg[4][27]  ( .D(n176), .CK(clk), .Q(\block[4][27] ) );
  DFFQXL \block_reg[4][26]  ( .D(n175), .CK(clk), .Q(\block[4][26] ) );
  DFFQXL \block_reg[4][25]  ( .D(n174), .CK(clk), .Q(\block[4][25] ) );
  DFFQXL \block_reg[4][24]  ( .D(n173), .CK(clk), .Q(\block[4][24] ) );
  DFFQXL \block_reg[4][23]  ( .D(n172), .CK(clk), .Q(\block[4][23] ) );
  DFFQXL \block_reg[4][22]  ( .D(n171), .CK(clk), .Q(\block[4][22] ) );
  DFFQXL \block_reg[4][21]  ( .D(n170), .CK(clk), .Q(\block[4][21] ) );
  DFFQXL \block_reg[4][20]  ( .D(n169), .CK(clk), .Q(\block[4][20] ) );
  DFFQXL \block_reg[3][31]  ( .D(n168), .CK(clk), .Q(\block[3][31] ) );
  DFFQXL \block_reg[3][30]  ( .D(n167), .CK(clk), .Q(\block[3][30] ) );
  DFFQXL \block_reg[3][29]  ( .D(n166), .CK(clk), .Q(\block[3][29] ) );
  DFFQXL \block_reg[3][28]  ( .D(n165), .CK(clk), .Q(\block[3][28] ) );
  CLKMX2X2 \block_reg[3][27]/U3  ( .A(\block[3][27] ), .B(block_next[27]), 
        .S0(n1565), .Y(n164) );
  DFFQXL \block_reg[3][27]  ( .D(n164), .CK(clk), .Q(\block[3][27] ) );
  DFFQXL \block_reg[3][26]  ( .D(n163), .CK(clk), .Q(\block[3][26] ) );
  DFFQXL \block_reg[3][25]  ( .D(n162), .CK(clk), .Q(\block[3][25] ) );
  DFFQXL \block_reg[3][24]  ( .D(n161), .CK(clk), .Q(\block[3][24] ) );
  DFFQXL \block_reg[3][23]  ( .D(n160), .CK(clk), .Q(\block[3][23] ) );
  DFFQXL \block_reg[3][22]  ( .D(n159), .CK(clk), .Q(\block[3][22] ) );
  DFFQXL \block_reg[3][21]  ( .D(n158), .CK(clk), .Q(\block[3][21] ) );
  DFFQXL \block_reg[3][20]  ( .D(n157), .CK(clk), .Q(\block[3][20] ) );
  DFFQXL \block_reg[2][31]  ( .D(n156), .CK(clk), .Q(\block[2][31] ) );
  DFFQXL \block_reg[2][30]  ( .D(n155), .CK(clk), .Q(\block[2][30] ) );
  DFFQXL \block_reg[2][29]  ( .D(n154), .CK(clk), .Q(\block[2][29] ) );
  DFFQXL \block_reg[2][28]  ( .D(n153), .CK(clk), .Q(\block[2][28] ) );
  CLKMX2X2 \block_reg[2][27]/U3  ( .A(\block[2][27] ), .B(block_next[27]), 
        .S0(n1578), .Y(n152) );
  DFFQXL \block_reg[2][27]  ( .D(n152), .CK(clk), .Q(\block[2][27] ) );
  DFFQXL \block_reg[2][26]  ( .D(n151), .CK(clk), .Q(\block[2][26] ) );
  DFFQXL \block_reg[2][25]  ( .D(n150), .CK(clk), .Q(\block[2][25] ) );
  DFFQXL \block_reg[2][24]  ( .D(n149), .CK(clk), .Q(\block[2][24] ) );
  DFFQXL \block_reg[2][23]  ( .D(n148), .CK(clk), .Q(\block[2][23] ) );
  DFFQXL \block_reg[2][22]  ( .D(n147), .CK(clk), .Q(\block[2][22] ) );
  DFFQXL \block_reg[2][21]  ( .D(n146), .CK(clk), .Q(\block[2][21] ) );
  DFFQXL \block_reg[2][20]  ( .D(n145), .CK(clk), .Q(\block[2][20] ) );
  DFFQXL \block_reg[1][31]  ( .D(n144), .CK(clk), .Q(\block[1][31] ) );
  DFFQXL \block_reg[1][30]  ( .D(n143), .CK(clk), .Q(\block[1][30] ) );
  DFFQXL \block_reg[1][29]  ( .D(n142), .CK(clk), .Q(\block[1][29] ) );
  DFFQXL \block_reg[1][28]  ( .D(n141), .CK(clk), .Q(\block[1][28] ) );
  CLKMX2X2 \block_reg[1][27]/U3  ( .A(\block[1][27] ), .B(block_next[27]), 
        .S0(n1592), .Y(n140) );
  DFFQXL \block_reg[1][27]  ( .D(n140), .CK(clk), .Q(\block[1][27] ) );
  DFFQXL \block_reg[1][26]  ( .D(n139), .CK(clk), .Q(\block[1][26] ) );
  DFFQXL \block_reg[1][25]  ( .D(n138), .CK(clk), .Q(\block[1][25] ) );
  DFFQXL \block_reg[1][24]  ( .D(n137), .CK(clk), .Q(\block[1][24] ) );
  DFFQXL \block_reg[1][23]  ( .D(n136), .CK(clk), .Q(\block[1][23] ) );
  DFFQXL \block_reg[1][22]  ( .D(n135), .CK(clk), .Q(\block[1][22] ) );
  DFFQXL \block_reg[1][21]  ( .D(n134), .CK(clk), .Q(\block[1][21] ) );
  DFFQXL \block_reg[1][20]  ( .D(n133), .CK(clk), .Q(\block[1][20] ) );
  DFFQXL \block_reg[0][28]  ( .D(n129), .CK(clk), .Q(\block[0][28] ) );
  CLKMX2X2 \block_reg[0][27]/U3  ( .A(\block[0][27] ), .B(block_next[27]), 
        .S0(n1607), .Y(n128) );
  DFFQXL \block_reg[0][27]  ( .D(n128), .CK(clk), .Q(\block[0][27] ) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n494), .CK(clk), .RN(n1628), .Q(
        blockdirty[7]), .QN(n478) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n490), .CK(clk), .RN(n1628), .Q(
        blockdirty[3]), .QN(n474) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n493), .CK(clk), .RN(n1628), .Q(
        blockdirty[6]), .QN(n477) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n489), .CK(clk), .RN(n1628), .Q(
        blockdirty[2]), .QN(n473) );
  EDFFXL \blocktag_reg[3][17]  ( .D(blocktag_next[17]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][17] ) );
  EDFFXL \blocktag_reg[7][17]  ( .D(blocktag_next[17]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][17] ) );
  EDFFXL \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][16] ) );
  EDFFXL \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][16] ) );
  EDFFXL \blocktag_reg[3][12]  ( .D(blocktag_next[12]), .E(n1561), .CK(clk), 
        .Q(\blocktag[3][12] ) );
  EDFFXL \blocktag_reg[3][14]  ( .D(blocktag_next[14]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][14] ) );
  EDFFXL \blocktag_reg[7][12]  ( .D(blocktag_next[12]), .E(n1496), .CK(clk), 
        .Q(\blocktag[7][12] ) );
  EDFFXL \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][22] ) );
  EDFFXL \blocktag_reg[7][14]  ( .D(blocktag_next[14]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][14] ) );
  EDFFXL \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][22] ) );
  EDFFXL \blocktag_reg[3][10]  ( .D(blocktag_next[10]), .E(n1561), .CK(clk), 
        .Q(\blocktag[3][10] ) );
  EDFFXL \blocktag_reg[7][10]  ( .D(blocktag_next[10]), .E(n1496), .CK(clk), 
        .Q(\blocktag[7][10] ) );
  EDFFXL \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][18] ) );
  EDFFXL \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][18] ) );
  EDFFXL \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFXL \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFXL \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFXL \blocktag_reg[3][5]  ( .D(blocktag_next[5]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFXL \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][2] ) );
  EDFFXL \blocktag_reg[7][5]  ( .D(blocktag_next[5]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFXL \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][6] ) );
  EDFFXL \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][6] ) );
  EDFFXL \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][9] ) );
  EDFFXL \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFXL \blocktag_reg[3][7]  ( .D(blocktag_next[7]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][7] ) );
  EDFFXL \blocktag_reg[7][7]  ( .D(blocktag_next[7]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][7] ) );
  EDFFXL \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFXL \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][1] ) );
  EDFFXL \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFXL \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][8] ) );
  EDFFXL \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFXL \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFXL \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFXL \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][13] ) );
  EDFFXL \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][4] ) );
  EDFFXL \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][4] ) );
  EDFFXL \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n1561), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFXL \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n1496), .CK(clk), 
        .Q(\blocktag[7][11] ) );
  EDFFXL \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][24] ) );
  EDFFXL \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][24] ) );
  EDFFXL \blocktag_reg[3][23]  ( .D(blocktag_next[23]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][23] ) );
  EDFFXL \blocktag_reg[7][23]  ( .D(blocktag_next[23]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][23] ) );
  EDFFXL \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n1561), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFXL \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n1496), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFXL \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][21] ) );
  EDFFXL \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][21] ) );
  EDFFXL \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][19] ) );
  EDFFXL \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][19] ) );
  EDFFXL \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n1562), .CK(clk), 
        .Q(\blocktag[3][20] ) );
  EDFFXL \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n1497), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFXL \blocktag_reg[1][17]  ( .D(blocktag_next[17]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][17] ) );
  EDFFXL \blocktag_reg[5][17]  ( .D(blocktag_next[17]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][17] ) );
  EDFFXL \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][16] ) );
  EDFFXL \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][16] ) );
  EDFFXL \blocktag_reg[1][12]  ( .D(blocktag_next[12]), .E(n1588), .CK(clk), 
        .Q(\blocktag[1][12] ) );
  EDFFXL \blocktag_reg[1][14]  ( .D(blocktag_next[14]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][14] ) );
  EDFFXL \blocktag_reg[5][12]  ( .D(blocktag_next[12]), .E(n1527), .CK(clk), 
        .Q(\blocktag[5][12] ) );
  EDFFXL \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][22] ) );
  EDFFXL \blocktag_reg[5][14]  ( .D(blocktag_next[14]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][14] ) );
  EDFFXL \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][22] ) );
  EDFFXL \blocktag_reg[1][10]  ( .D(blocktag_next[10]), .E(n1588), .CK(clk), 
        .Q(\blocktag[1][10] ) );
  EDFFXL \blocktag_reg[5][10]  ( .D(blocktag_next[10]), .E(n1527), .CK(clk), 
        .Q(\blocktag[5][10] ) );
  EDFFXL \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][18] ) );
  EDFFXL \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][18] ) );
  EDFFXL \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFXL \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFXL \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFXL \blocktag_reg[1][5]  ( .D(blocktag_next[5]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFXL \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][2] ) );
  EDFFXL \blocktag_reg[5][5]  ( .D(blocktag_next[5]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFXL \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][6] ) );
  EDFFXL \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][6] ) );
  EDFFXL \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFXL \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFXL \blocktag_reg[1][7]  ( .D(blocktag_next[7]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][7] ) );
  EDFFXL \blocktag_reg[5][7]  ( .D(blocktag_next[7]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][7] ) );
  EDFFXL \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFXL \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][1] ) );
  EDFFXL \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFXL \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][8] ) );
  EDFFXL \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFXL \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFXL \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFXL \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][13] ) );
  EDFFXL \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][4] ) );
  EDFFXL \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][4] ) );
  EDFFXL \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n1588), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFXL \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n1527), .CK(clk), 
        .Q(\blocktag[5][11] ) );
  EDFFXL \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][24] ) );
  EDFFXL \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][24] ) );
  EDFFXL \blocktag_reg[1][23]  ( .D(blocktag_next[23]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][23] ) );
  EDFFXL \blocktag_reg[5][23]  ( .D(blocktag_next[23]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][23] ) );
  EDFFXL \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n1588), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFXL \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(n1527), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFXL \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][21] ) );
  EDFFXL \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][21] ) );
  EDFFXL \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][19] ) );
  EDFFXL \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][19] ) );
  EDFFXL \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n1589), .CK(clk), 
        .Q(\blocktag[1][20] ) );
  EDFFXL \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n1528), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFXL \blocktag_reg[0][17]  ( .D(blocktag_next[17]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][17] ) );
  EDFFXL \blocktag_reg[4][17]  ( .D(blocktag_next[17]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][17] ) );
  EDFFXL \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][16] ) );
  EDFFXL \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][16] ) );
  EDFFXL \blocktag_reg[0][12]  ( .D(blocktag_next[12]), .E(n1603), .CK(clk), 
        .Q(\blocktag[0][12] ) );
  EDFFXL \blocktag_reg[0][14]  ( .D(blocktag_next[14]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][14] ) );
  EDFFXL \blocktag_reg[4][12]  ( .D(blocktag_next[12]), .E(n1544), .CK(clk), 
        .Q(\blocktag[4][12] ) );
  EDFFXL \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][22] ) );
  EDFFXL \blocktag_reg[4][14]  ( .D(blocktag_next[14]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][14] ) );
  EDFFXL \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][22] ) );
  EDFFXL \blocktag_reg[0][10]  ( .D(blocktag_next[10]), .E(n1603), .CK(clk), 
        .Q(\blocktag[0][10] ) );
  EDFFXL \blocktag_reg[4][10]  ( .D(blocktag_next[10]), .E(n1544), .CK(clk), 
        .Q(\blocktag[4][10] ) );
  EDFFXL \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][18] ) );
  EDFFXL \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][18] ) );
  EDFFXL \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFXL \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFXL \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFXL \blocktag_reg[0][5]  ( .D(blocktag_next[5]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFXL \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][2] ) );
  EDFFXL \blocktag_reg[4][5]  ( .D(blocktag_next[5]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFXL \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][6] ) );
  EDFFXL \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][6] ) );
  EDFFXL \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFXL \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFXL \blocktag_reg[0][7]  ( .D(blocktag_next[7]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][7] ) );
  EDFFXL \blocktag_reg[4][7]  ( .D(blocktag_next[7]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][7] ) );
  EDFFXL \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFXL \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][1] ) );
  EDFFXL \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFXL \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][8] ) );
  EDFFXL \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFXL \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFXL \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFXL \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][13] ) );
  EDFFXL \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][4] ) );
  EDFFXL \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][4] ) );
  EDFFXL \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n1603), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFXL \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n1544), .CK(clk), 
        .Q(\blocktag[4][11] ) );
  EDFFXL \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][24] ) );
  EDFFXL \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][24] ) );
  EDFFXL \blocktag_reg[0][23]  ( .D(blocktag_next[23]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][23] ) );
  EDFFXL \blocktag_reg[4][23]  ( .D(blocktag_next[23]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][23] ) );
  EDFFXL \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n1603), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFXL \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n1544), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFXL \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][21] ) );
  EDFFXL \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][21] ) );
  EDFFXL \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][19] ) );
  EDFFXL \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][19] ) );
  EDFFXL \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n1604), .CK(clk), 
        .Q(\blocktag[0][20] ) );
  EDFFXL \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n1545), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFXL \blocktag_reg[2][17]  ( .D(blocktag_next[17]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][17] ) );
  EDFFXL \blocktag_reg[6][17]  ( .D(blocktag_next[17]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][17] ) );
  EDFFXL \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][16] ) );
  EDFFXL \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][16] ) );
  EDFFXL \blocktag_reg[2][12]  ( .D(blocktag_next[12]), .E(n1574), .CK(clk), 
        .Q(\blocktag[2][12] ) );
  EDFFXL \blocktag_reg[2][14]  ( .D(blocktag_next[14]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][14] ) );
  EDFFXL \blocktag_reg[6][12]  ( .D(blocktag_next[12]), .E(n1511), .CK(clk), 
        .Q(\blocktag[6][12] ) );
  EDFFXL \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][22] ) );
  EDFFXL \blocktag_reg[6][14]  ( .D(blocktag_next[14]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][14] ) );
  EDFFXL \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][22] ) );
  EDFFXL \blocktag_reg[2][10]  ( .D(blocktag_next[10]), .E(n1574), .CK(clk), 
        .Q(\blocktag[2][10] ) );
  EDFFXL \blocktag_reg[6][10]  ( .D(blocktag_next[10]), .E(n1511), .CK(clk), 
        .Q(\blocktag[6][10] ) );
  EDFFXL \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][18] ) );
  EDFFXL \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][18] ) );
  EDFFXL \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFXL \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFXL \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFXL \blocktag_reg[2][5]  ( .D(blocktag_next[5]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFXL \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][2] ) );
  EDFFXL \blocktag_reg[6][5]  ( .D(blocktag_next[5]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFXL \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][6] ) );
  EDFFXL \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][6] ) );
  EDFFXL \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFXL \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFXL \blocktag_reg[2][7]  ( .D(blocktag_next[7]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][7] ) );
  EDFFXL \blocktag_reg[6][7]  ( .D(blocktag_next[7]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][7] ) );
  EDFFXL \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFXL \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][1] ) );
  EDFFXL \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFXL \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][8] ) );
  EDFFXL \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFXL \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFXL \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFXL \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][13] ) );
  EDFFXL \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][4] ) );
  EDFFXL \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][4] ) );
  EDFFXL \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n1574), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFXL \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n1511), .CK(clk), 
        .Q(\blocktag[6][11] ) );
  EDFFXL \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][24] ) );
  EDFFXL \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][24] ) );
  EDFFXL \blocktag_reg[2][23]  ( .D(blocktag_next[23]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][23] ) );
  EDFFXL \blocktag_reg[6][23]  ( .D(blocktag_next[23]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][23] ) );
  EDFFXL \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n1574), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFXL \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n1511), .CK(clk), .Q(
        \blocktag[6][0] ) );
  EDFFXL \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][21] ) );
  EDFFXL \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][21] ) );
  EDFFXL \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][19] ) );
  EDFFXL \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][19] ) );
  EDFFXL \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n1575), .CK(clk), 
        .Q(\blocktag[2][20] ) );
  EDFFXL \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n1512), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n492), .CK(clk), .RN(n1628), .Q(
        blockdirty[5]), .QN(n476) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n488), .CK(clk), .RN(n1628), .Q(
        blockdirty[1]), .QN(n472) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n491), .CK(clk), .RN(n1628), .Q(
        blockdirty[4]), .QN(n475) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n487), .CK(clk), .RN(n1628), .Q(
        blockdirty[0]), .QN(n471) );
  DFFSRXL \blockvalid_reg[6]  ( .D(n501), .CK(clk), .SN(1'b1), .RN(n1629), .Q(
        blockvalid[6]), .QN(n485) );
  DFFSRXL \blockvalid_reg[2]  ( .D(n497), .CK(clk), .SN(1'b1), .RN(n1629), .Q(
        blockvalid[2]), .QN(n481) );
  DFFSRXL \blockvalid_reg[1]  ( .D(n496), .CK(clk), .SN(1'b1), .RN(n1629), .Q(
        blockvalid[1]), .QN(n480) );
  DFFSRXL \blockvalid_reg[0]  ( .D(n495), .CK(clk), .SN(1'b1), .RN(n1629), .Q(
        blockvalid[0]), .QN(n479) );
  EDFFXL \block_reg[7][55]  ( .D(block_next[55]), .E(n1502), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFXL \block_reg[6][55]  ( .D(block_next[55]), .E(n5), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFXL \block_reg[5][55]  ( .D(block_next[55]), .E(n7), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFXL \block_reg[4][55]  ( .D(block_next[55]), .E(n6), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFXL \block_reg[3][55]  ( .D(block_next[55]), .E(n3), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFXL \block_reg[2][55]  ( .D(block_next[55]), .E(n2), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFXL \block_reg[1][55]  ( .D(block_next[55]), .E(n1), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFXL \block_reg[0][55]  ( .D(block_next[55]), .E(n4), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFXL \block_reg[7][117]  ( .D(block_next[117]), .E(n2124), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFXL \block_reg[7][116]  ( .D(block_next[116]), .E(n2124), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFXL \block_reg[6][117]  ( .D(block_next[117]), .E(n5), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFXL \block_reg[6][116]  ( .D(block_next[116]), .E(n5), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFXL \block_reg[5][117]  ( .D(block_next[117]), .E(n7), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFXL \block_reg[5][116]  ( .D(block_next[116]), .E(n7), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFXL \block_reg[4][117]  ( .D(block_next[117]), .E(n6), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFXL \block_reg[4][116]  ( .D(block_next[116]), .E(n6), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFXL \block_reg[3][117]  ( .D(block_next[117]), .E(n3), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFXL \block_reg[3][116]  ( .D(block_next[116]), .E(n3), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFXL \block_reg[2][117]  ( .D(block_next[117]), .E(n2), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFXL \block_reg[2][116]  ( .D(block_next[116]), .E(n2), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFXL \block_reg[1][117]  ( .D(block_next[117]), .E(n1), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFXL \block_reg[1][116]  ( .D(block_next[116]), .E(n1), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFXL \block_reg[7][118]  ( .D(block_next[118]), .E(n2124), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFXL \block_reg[6][118]  ( .D(block_next[118]), .E(n5), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFXL \block_reg[5][118]  ( .D(block_next[118]), .E(n7), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFXL \block_reg[4][118]  ( .D(block_next[118]), .E(n6), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFXL \block_reg[3][118]  ( .D(block_next[118]), .E(n3), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFXL \block_reg[2][118]  ( .D(block_next[118]), .E(n2), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFXL \block_reg[1][118]  ( .D(block_next[118]), .E(n1), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFXL \block_reg[0][124]  ( .D(block_next[124]), .E(n4), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFXL \block_reg[0][123]  ( .D(block_next[123]), .E(n4), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFXL \block_reg[7][124]  ( .D(block_next[124]), .E(n2124), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFXL \block_reg[7][123]  ( .D(block_next[123]), .E(n2124), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFXL \block_reg[6][124]  ( .D(block_next[124]), .E(n5), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFXL \block_reg[6][123]  ( .D(block_next[123]), .E(n5), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFXL \block_reg[5][124]  ( .D(block_next[124]), .E(n7), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFXL \block_reg[5][123]  ( .D(block_next[123]), .E(n7), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFXL \block_reg[4][124]  ( .D(block_next[124]), .E(n6), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFXL \block_reg[4][123]  ( .D(block_next[123]), .E(n6), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFXL \block_reg[3][124]  ( .D(block_next[124]), .E(n3), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFXL \block_reg[3][123]  ( .D(block_next[123]), .E(n3), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFXL \block_reg[2][124]  ( .D(block_next[124]), .E(n2), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFXL \block_reg[2][123]  ( .D(block_next[123]), .E(n2), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFXL \block_reg[1][124]  ( .D(block_next[124]), .E(n1), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFXL \block_reg[1][123]  ( .D(block_next[123]), .E(n1), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFXL \block_reg[0][127]  ( .D(block_next[127]), .E(n4), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFXL \block_reg[0][126]  ( .D(block_next[126]), .E(n4), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFXL \block_reg[0][125]  ( .D(block_next[125]), .E(n4), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFXL \block_reg[0][122]  ( .D(block_next[122]), .E(n4), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFXL \block_reg[0][121]  ( .D(block_next[121]), .E(n4), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFXL \block_reg[0][120]  ( .D(block_next[120]), .E(n4), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFXL \block_reg[7][127]  ( .D(block_next[127]), .E(n2124), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFXL \block_reg[7][126]  ( .D(block_next[126]), .E(n2124), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFXL \block_reg[7][125]  ( .D(block_next[125]), .E(n2124), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFXL \block_reg[7][122]  ( .D(block_next[122]), .E(n2124), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFXL \block_reg[7][121]  ( .D(block_next[121]), .E(n2124), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFXL \block_reg[7][120]  ( .D(block_next[120]), .E(n2124), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFXL \block_reg[6][127]  ( .D(block_next[127]), .E(n5), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFXL \block_reg[6][126]  ( .D(block_next[126]), .E(n5), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFXL \block_reg[6][125]  ( .D(block_next[125]), .E(n5), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFXL \block_reg[6][122]  ( .D(block_next[122]), .E(n5), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFXL \block_reg[6][121]  ( .D(block_next[121]), .E(n5), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFXL \block_reg[6][120]  ( .D(block_next[120]), .E(n5), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFXL \block_reg[5][127]  ( .D(block_next[127]), .E(n7), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFXL \block_reg[5][126]  ( .D(block_next[126]), .E(n7), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFXL \block_reg[5][125]  ( .D(block_next[125]), .E(n7), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFXL \block_reg[5][122]  ( .D(block_next[122]), .E(n7), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFXL \block_reg[5][121]  ( .D(block_next[121]), .E(n7), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFXL \block_reg[5][120]  ( .D(block_next[120]), .E(n7), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFXL \block_reg[4][127]  ( .D(block_next[127]), .E(n6), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFXL \block_reg[4][126]  ( .D(block_next[126]), .E(n6), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFXL \block_reg[4][125]  ( .D(block_next[125]), .E(n6), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFXL \block_reg[4][122]  ( .D(block_next[122]), .E(n6), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFXL \block_reg[4][121]  ( .D(block_next[121]), .E(n6), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFXL \block_reg[4][120]  ( .D(block_next[120]), .E(n6), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFXL \block_reg[3][127]  ( .D(block_next[127]), .E(n3), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFXL \block_reg[3][126]  ( .D(block_next[126]), .E(n3), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFXL \block_reg[3][125]  ( .D(block_next[125]), .E(n3), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFXL \block_reg[3][122]  ( .D(block_next[122]), .E(n3), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFXL \block_reg[3][121]  ( .D(block_next[121]), .E(n3), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFXL \block_reg[3][120]  ( .D(block_next[120]), .E(n3), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFXL \block_reg[2][127]  ( .D(block_next[127]), .E(n2), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFXL \block_reg[2][126]  ( .D(block_next[126]), .E(n2), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFXL \block_reg[2][125]  ( .D(block_next[125]), .E(n2), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFXL \block_reg[2][122]  ( .D(block_next[122]), .E(n2), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFXL \block_reg[2][121]  ( .D(block_next[121]), .E(n2), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFXL \block_reg[2][120]  ( .D(block_next[120]), .E(n2), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFXL \block_reg[1][127]  ( .D(block_next[127]), .E(n1), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFXL \block_reg[1][126]  ( .D(block_next[126]), .E(n1), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFXL \block_reg[1][125]  ( .D(block_next[125]), .E(n1), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFXL \block_reg[1][122]  ( .D(block_next[122]), .E(n1), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFXL \block_reg[1][121]  ( .D(block_next[121]), .E(n1), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFXL \block_reg[1][120]  ( .D(block_next[120]), .E(n1), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFXL \block_reg[0][119]  ( .D(block_next[119]), .E(n4), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFXL \block_reg[7][119]  ( .D(block_next[119]), .E(n2124), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFXL \block_reg[6][119]  ( .D(block_next[119]), .E(n5), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFXL \block_reg[5][119]  ( .D(block_next[119]), .E(n7), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFXL \block_reg[4][119]  ( .D(block_next[119]), .E(n6), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFXL \block_reg[3][119]  ( .D(block_next[119]), .E(n3), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFXL \block_reg[2][119]  ( .D(block_next[119]), .E(n2), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFXL \block_reg[1][119]  ( .D(block_next[119]), .E(n1), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFXL \block_reg[7][96]  ( .D(block_next[96]), .E(n2124), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFXL \block_reg[6][96]  ( .D(block_next[96]), .E(n5), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFXL \block_reg[0][106]  ( .D(block_next[106]), .E(n4), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFXL \block_reg[7][106]  ( .D(block_next[106]), .E(n2124), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFXL \block_reg[6][106]  ( .D(block_next[106]), .E(n5), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFXL \block_reg[5][106]  ( .D(block_next[106]), .E(n7), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFXL \block_reg[4][106]  ( .D(block_next[106]), .E(n6), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFXL \block_reg[3][106]  ( .D(block_next[106]), .E(n3), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFXL \block_reg[2][106]  ( .D(block_next[106]), .E(n2), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFXL \block_reg[1][106]  ( .D(block_next[106]), .E(n1), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFXL \block_reg[5][104]  ( .D(block_next[104]), .E(n7), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFXL \block_reg[4][104]  ( .D(block_next[104]), .E(n6), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFXL \block_reg[3][104]  ( .D(block_next[104]), .E(n3), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFXL \block_reg[2][104]  ( .D(block_next[104]), .E(n2), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFXL \block_reg[1][104]  ( .D(block_next[104]), .E(n1), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFXL \block_reg[0][104]  ( .D(block_next[104]), .E(n4), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFXL \block_reg[7][104]  ( .D(block_next[104]), .E(n2124), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFXL \block_reg[6][104]  ( .D(block_next[104]), .E(n5), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFXL \block_reg[1][18]  ( .D(block_next[18]), .E(n1), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFXL \block_reg[0][18]  ( .D(block_next[18]), .E(n4), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFXL \block_reg[5][98]  ( .D(block_next[98]), .E(n7), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFXL \block_reg[4][98]  ( .D(block_next[98]), .E(n6), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFXL \block_reg[3][98]  ( .D(block_next[98]), .E(n3), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFXL \block_reg[2][98]  ( .D(block_next[98]), .E(n2), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFXL \block_reg[1][98]  ( .D(block_next[98]), .E(n1), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFXL \block_reg[0][98]  ( .D(block_next[98]), .E(n4), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFXL \block_reg[5][97]  ( .D(block_next[97]), .E(n7), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFXL \block_reg[4][97]  ( .D(block_next[97]), .E(n6), .CK(clk), .Q(
        \block[4][97] ) );
  DFFHQX2 \block_reg[0][51]  ( .D(n228), .CK(clk), .Q(\block[0][51] ) );
  DFFHQX2 \block_reg[0][38]  ( .D(n581), .CK(clk), .Q(\block[0][38] ) );
  DFFHQX2 \block_reg[5][71]  ( .D(n1031), .CK(clk), .Q(\block[5][71] ) );
  DFFQXL \block_reg[0][31]  ( .D(n132), .CK(clk), .Q(\block[0][31] ) );
  DFFQXL \block_reg[0][30]  ( .D(n131), .CK(clk), .Q(\block[0][30] ) );
  DFFQXL \block_reg[0][20]  ( .D(n121), .CK(clk), .Q(\block[0][20] ) );
  DFFQXL \block_reg[0][23]  ( .D(n124), .CK(clk), .Q(\block[0][23] ) );
  DFFQXL \block_reg[0][26]  ( .D(n127), .CK(clk), .Q(\block[0][26] ) );
  DFFQXL \block_reg[0][22]  ( .D(n123), .CK(clk), .Q(\block[0][22] ) );
  DFFQXL \block_reg[0][24]  ( .D(n125), .CK(clk), .Q(\block[0][24] ) );
  DFFQXL \block_reg[0][21]  ( .D(n122), .CK(clk), .Q(\block[0][21] ) );
  DFFQXL \block_reg[0][25]  ( .D(n126), .CK(clk), .Q(\block[0][25] ) );
  DFFHQX2 \block_reg[0][67]  ( .D(n987), .CK(clk), .Q(\block[0][67] ) );
  DFFHQX2 \block_reg[7][80]  ( .D(n914), .CK(clk), .Q(\block[7][80] ) );
  DFFHQX2 \block_reg[7][79]  ( .D(n913), .CK(clk), .Q(\block[7][79] ) );
  DFFHQX2 \block_reg[7][85]  ( .D(n919), .CK(clk), .Q(\block[7][85] ) );
  DFFHQX2 \block_reg[7][82]  ( .D(n916), .CK(clk), .Q(\block[7][82] ) );
  DFFHQX2 \block_reg[7][87]  ( .D(n921), .CK(clk), .Q(\block[7][87] ) );
  DFFHQX2 \block_reg[7][81]  ( .D(n915), .CK(clk), .Q(\block[7][81] ) );
  DFFHQX2 \block_reg[7][84]  ( .D(n918), .CK(clk), .Q(\block[7][84] ) );
  DFFHQX2 \block_reg[7][77]  ( .D(n911), .CK(clk), .Q(\block[7][77] ) );
  DFFHQX2 \block_reg[7][83]  ( .D(n917), .CK(clk), .Q(\block[7][83] ) );
  DFFHQX2 \block_reg[2][72]  ( .D(n786), .CK(clk), .Q(\block[2][72] ) );
  DFFHQX2 \block_reg[2][74]  ( .D(n788), .CK(clk), .Q(\block[2][74] ) );
  DFFHQX2 \block_reg[2][73]  ( .D(n787), .CK(clk), .Q(\block[2][73] ) );
  DFFHQX2 \block_reg[2][76]  ( .D(n790), .CK(clk), .Q(\block[2][76] ) );
  DFFHQX4 \block_reg[2][75]  ( .D(n789), .CK(clk), .Q(\block[2][75] ) );
  DFFQXL \block_reg[0][29]  ( .D(n130), .CK(clk), .Q(\block[0][29] ) );
  DFFQXL \block_reg[0][99]  ( .D(n932), .CK(clk), .Q(\block[0][99] ) );
  DFFQX1 \block_reg[0][0]  ( .D(n511), .CK(clk), .Q(\block[0][0] ) );
  CLKINVX2 U3 ( .A(n1664), .Y(n16) );
  MXI4X1 U4 ( .A(\blocktag[4][8] ), .B(\blocktag[5][8] ), .C(\blocktag[6][8] ), 
        .D(\blocktag[7][8] ), .S0(n1446), .S1(n1412), .Y(n1341) );
  INVX4 U5 ( .A(tag[8]), .Y(n1902) );
  MXI4X1 U6 ( .A(\blocktag[0][8] ), .B(\blocktag[1][8] ), .C(\blocktag[2][8] ), 
        .D(\blocktag[3][8] ), .S0(n1446), .S1(n1412), .Y(n1340) );
  INVX3 U7 ( .A(tag[10]), .Y(n1896) );
  MXI4X2 U8 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n1446), .S1(n1412), .Y(
        n1336) );
  MXI4X2 U9 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n1446), .S1(n1412), .Y(
        n1337) );
  MXI2X4 U10 ( .A(n1340), .B(n1341), .S0(n1375), .Y(tag[8]) );
  INVX8 U11 ( .A(tag[11]), .Y(n1893) );
  MXI2X4 U12 ( .A(n1334), .B(n1335), .S0(n1375), .Y(tag[11]) );
  AO22XL U13 ( .A0(proc_addr[18]), .A1(mem_read), .B0(tag[13]), .B1(mem_write), 
        .Y(mem_addr[16]) );
  INVX8 U14 ( .A(tag[13]), .Y(n1887) );
  MXI2X4 U15 ( .A(n1330), .B(n1331), .S0(n1374), .Y(tag[13]) );
  MXI2X4 U16 ( .A(n1336), .B(n1337), .S0(n1375), .Y(tag[10]) );
  INVX3 U17 ( .A(n1619), .Y(n120) );
  BUFX8 U18 ( .A(n2121), .Y(n1491) );
  INVX1 U19 ( .A(mem_write), .Y(n108) );
  INVX1 U20 ( .A(mem_write), .Y(n100) );
  INVX1 U21 ( .A(mem_write), .Y(n86) );
  INVX1 U22 ( .A(mem_write), .Y(n81) );
  INVX1 U23 ( .A(mem_write), .Y(n76) );
  INVX1 U24 ( .A(mem_write), .Y(n72) );
  INVX3 U25 ( .A(n1953), .Y(n2125) );
  INVX3 U26 ( .A(tag[20]), .Y(n1869) );
  INVX3 U27 ( .A(tag[19]), .Y(n1872) );
  INVX3 U28 ( .A(tag[4]), .Y(n1914) );
  BUFX16 U29 ( .A(N33), .Y(n1376) );
  INVX12 U30 ( .A(N31), .Y(n1619) );
  CLKINVX1 U31 ( .A(mem_ready), .Y(n1947) );
  INVX8 U32 ( .A(n1469), .Y(n1465) );
  BUFX16 U33 ( .A(n1750), .Y(n1457) );
  INVX3 U34 ( .A(blockdata[1]), .Y(n1969) );
  CLKINVX12 U35 ( .A(n14), .Y(n29) );
  INVX3 U36 ( .A(tag[21]), .Y(n1866) );
  INVX3 U37 ( .A(tag[23]), .Y(n1860) );
  INVX6 U38 ( .A(tag[6]), .Y(n1908) );
  INVX3 U39 ( .A(tag[17]), .Y(n1877) );
  INVX8 U40 ( .A(n43), .Y(n44) );
  INVX6 U41 ( .A(block_next[14]), .Y(n43) );
  INVX8 U42 ( .A(n41), .Y(n42) );
  INVX6 U43 ( .A(block_next[16]), .Y(n41) );
  NOR2X4 U44 ( .A(n110), .B(n111), .Y(n107) );
  NOR2X4 U45 ( .A(n103), .B(n104), .Y(n99) );
  NOR2X4 U46 ( .A(n89), .B(n90), .Y(n85) );
  NOR2X4 U47 ( .A(n83), .B(n84), .Y(n80) );
  NOR2X4 U48 ( .A(n78), .B(n79), .Y(n75) );
  NOR2X4 U49 ( .A(n73), .B(n74), .Y(n71) );
  OAI221X1 U50 ( .A0(n31), .A1(n1999), .B0(n1493), .B1(n1998), .C0(n1997), .Y(
        proc_rdata[7]) );
  INVXL U51 ( .A(tag[9]), .Y(n1899) );
  BUFX2 U52 ( .A(n1415), .Y(n1379) );
  BUFX2 U53 ( .A(n1416), .Y(n1378) );
  INVX1 U54 ( .A(N32), .Y(n1620) );
  BUFX2 U55 ( .A(n1448), .Y(n1417) );
  INVX16 U56 ( .A(N33), .Y(n1621) );
  BUFX16 U57 ( .A(N32), .Y(n1414) );
  CLKAND2X12 U58 ( .A(n1929), .B(n1628), .Y(n1) );
  CLKAND2X12 U59 ( .A(n1931), .B(n1628), .Y(n2) );
  AND2X8 U60 ( .A(n1933), .B(n1628), .Y(n3) );
  BUFX16 U61 ( .A(n1449), .Y(n1418) );
  CLKAND2X12 U62 ( .A(n1857), .B(n1628), .Y(n4) );
  AND2X8 U63 ( .A(n1940), .B(n1628), .Y(n5) );
  INVX16 U64 ( .A(n1943), .Y(n2124) );
  BUFX2 U65 ( .A(n2124), .Y(n1507) );
  BUFX4 U66 ( .A(n1359), .Y(n1370) );
  BUFX2 U67 ( .A(n4), .Y(n1615) );
  BUFX4 U68 ( .A(n1448), .Y(n1433) );
  AND2X8 U69 ( .A(n1935), .B(n1628), .Y(n6) );
  BUFX2 U70 ( .A(n1), .Y(n1599) );
  AND2X8 U71 ( .A(n1937), .B(n1628), .Y(n7) );
  AND2X4 U72 ( .A(mem_ready), .B(n1950), .Y(n8) );
  BUFX2 U73 ( .A(n2), .Y(n1586) );
  BUFX2 U74 ( .A(n1510), .Y(n1522) );
  BUFX2 U75 ( .A(n1380), .Y(n1385) );
  INVX1 U76 ( .A(mem_read), .Y(n109) );
  INVX1 U77 ( .A(mem_read), .Y(n82) );
  CLKMX2X4 U78 ( .A(n1326), .B(n1327), .S0(n1374), .Y(n9) );
  BUFX2 U79 ( .A(n1360), .Y(n1363) );
  BUFX2 U80 ( .A(n1415), .Y(n1377) );
  AND3X8 U81 ( .A(n1851), .B(n1752), .C(n1751), .Y(n10) );
  BUFX16 U82 ( .A(n1488), .Y(n1479) );
  AND2X6 U83 ( .A(proc_read), .B(n1665), .Y(n11) );
  CLKAND2X12 U84 ( .A(n1752), .B(n1461), .Y(n12) );
  CLKINVX4 U85 ( .A(n1951), .Y(n2126) );
  CLKINVX12 U86 ( .A(proc_addr[29]), .Y(n40) );
  CLKBUFX2 U87 ( .A(n7), .Y(n1526) );
  INVXL U88 ( .A(proc_addr[19]), .Y(n88) );
  CLKBUFX2 U89 ( .A(n1602), .Y(n1614) );
  BUFX4 U90 ( .A(n1614), .Y(n1613) );
  BUFX12 U91 ( .A(n5), .Y(n1510) );
  INVX1 U92 ( .A(proc_reset), .Y(n1629) );
  BUFX6 U93 ( .A(n1629), .Y(n1628) );
  XOR2X4 U94 ( .A(n1884), .B(proc_addr[19]), .Y(n1641) );
  INVX3 U95 ( .A(tag[14]), .Y(n1884) );
  INVXL U96 ( .A(n1382), .Y(n13) );
  BUFX20 U97 ( .A(n1381), .Y(n1382) );
  NAND2XL U98 ( .A(N32), .B(N33), .Y(n1938) );
  CLKBUFX2 U99 ( .A(n1414), .Y(n1415) );
  NAND2X8 U100 ( .A(n1715), .B(n1456), .Y(n1716) );
  INVX12 U101 ( .A(n1716), .Y(n1752) );
  OAI221X4 U102 ( .A0(n31), .A1(n2084), .B0(n1495), .B1(n2083), .C0(n2082), 
        .Y(proc_rdata[24]) );
  MX2X1 U103 ( .A(\block[2][75] ), .B(block_next[75]), .S0(n1581), .Y(n789) );
  OAI221X4 U104 ( .A0(n1458), .A1(n2016), .B0(n1827), .B1(n1459), .C0(n1738), 
        .Y(block_next[75]) );
  MX2X1 U105 ( .A(\block[2][76] ), .B(block_next[76]), .S0(n1581), .Y(n790) );
  MX2X1 U106 ( .A(\block[7][76] ), .B(block_next[76]), .S0(n1503), .Y(n910) );
  MX2X1 U107 ( .A(\block[6][76] ), .B(block_next[76]), .S0(n1518), .Y(n886) );
  MX2X1 U108 ( .A(\block[5][76] ), .B(block_next[76]), .S0(n1534), .Y(n862) );
  MX2X1 U109 ( .A(\block[4][76] ), .B(block_next[76]), .S0(n1551), .Y(n838) );
  MX2X1 U110 ( .A(\block[3][76] ), .B(block_next[76]), .S0(n1568), .Y(n814) );
  MX2X1 U111 ( .A(\block[1][76] ), .B(block_next[76]), .S0(n1595), .Y(n766) );
  MX2X1 U112 ( .A(\block[0][76] ), .B(block_next[76]), .S0(n1610), .Y(n742) );
  OAI221X4 U113 ( .A0(n1458), .A1(n2021), .B0(n1825), .B1(n1459), .C0(n1737), 
        .Y(block_next[76]) );
  MX2X1 U114 ( .A(\block[2][73] ), .B(block_next[73]), .S0(n1581), .Y(n787) );
  MX2X1 U115 ( .A(\block[7][73] ), .B(block_next[73]), .S0(n1503), .Y(n907) );
  MX2X1 U116 ( .A(\block[6][73] ), .B(block_next[73]), .S0(n1518), .Y(n883) );
  MX2X1 U117 ( .A(\block[5][73] ), .B(block_next[73]), .S0(n1534), .Y(n859) );
  MX2X1 U118 ( .A(\block[4][73] ), .B(block_next[73]), .S0(n1551), .Y(n835) );
  MX2X1 U119 ( .A(\block[3][73] ), .B(block_next[73]), .S0(n1568), .Y(n811) );
  MX2X1 U120 ( .A(\block[1][73] ), .B(block_next[73]), .S0(n1595), .Y(n763) );
  MX2X1 U121 ( .A(\block[0][73] ), .B(block_next[73]), .S0(n1610), .Y(n739) );
  OAI221X4 U122 ( .A0(n1458), .A1(n2006), .B0(n1831), .B1(n1459), .C0(n1740), 
        .Y(block_next[73]) );
  MX2X1 U123 ( .A(\block[2][74] ), .B(block_next[74]), .S0(n1581), .Y(n788) );
  MX2X1 U124 ( .A(\block[7][74] ), .B(block_next[74]), .S0(n1503), .Y(n908) );
  MX2X1 U125 ( .A(\block[6][74] ), .B(block_next[74]), .S0(n1518), .Y(n884) );
  MX2X1 U126 ( .A(\block[5][74] ), .B(block_next[74]), .S0(n1534), .Y(n860) );
  MX2X1 U127 ( .A(\block[4][74] ), .B(block_next[74]), .S0(n1551), .Y(n836) );
  MX2X1 U128 ( .A(\block[3][74] ), .B(block_next[74]), .S0(n1568), .Y(n812) );
  MX2X1 U129 ( .A(\block[1][74] ), .B(block_next[74]), .S0(n1595), .Y(n764) );
  MX2X1 U130 ( .A(\block[0][74] ), .B(block_next[74]), .S0(n1610), .Y(n740) );
  OAI221X4 U131 ( .A0(n1458), .A1(n2011), .B0(n1829), .B1(n1459), .C0(n1739), 
        .Y(block_next[74]) );
  MX2X1 U132 ( .A(\block[2][72] ), .B(block_next[72]), .S0(n1581), .Y(n786) );
  MX2X1 U133 ( .A(\block[7][72] ), .B(block_next[72]), .S0(n1503), .Y(n906) );
  MX2X1 U134 ( .A(\block[6][72] ), .B(block_next[72]), .S0(n1518), .Y(n882) );
  MX2X1 U135 ( .A(\block[5][72] ), .B(block_next[72]), .S0(n1534), .Y(n858) );
  MX2X1 U136 ( .A(\block[4][72] ), .B(block_next[72]), .S0(n1551), .Y(n834) );
  MX2X1 U137 ( .A(\block[3][72] ), .B(block_next[72]), .S0(n1568), .Y(n810) );
  MX2X1 U138 ( .A(\block[1][72] ), .B(block_next[72]), .S0(n1595), .Y(n762) );
  MX2X1 U139 ( .A(\block[0][72] ), .B(block_next[72]), .S0(n1610), .Y(n738) );
  OAI221X4 U140 ( .A0(n1458), .A1(n2001), .B0(n1833), .B1(n1459), .C0(n1741), 
        .Y(block_next[72]) );
  INVX3 U141 ( .A(n2118), .Y(n14) );
  NAND3BX1 U142 ( .AN(n1959), .B(proc_addr[1]), .C(n1957), .Y(n2118) );
  MX2X1 U143 ( .A(\block[7][83] ), .B(block_next[83]), .S0(n1504), .Y(n917) );
  MX2X1 U144 ( .A(\block[6][83] ), .B(block_next[83]), .S0(n1519), .Y(n893) );
  MX2X1 U145 ( .A(\block[5][83] ), .B(block_next[83]), .S0(n1535), .Y(n869) );
  MX2X1 U146 ( .A(\block[4][83] ), .B(block_next[83]), .S0(n1552), .Y(n845) );
  MX2X1 U147 ( .A(\block[3][83] ), .B(block_next[83]), .S0(n1569), .Y(n821) );
  MX2X1 U148 ( .A(\block[2][83] ), .B(block_next[83]), .S0(n1582), .Y(n797) );
  MX2X1 U149 ( .A(\block[1][83] ), .B(block_next[83]), .S0(n1596), .Y(n773) );
  MX2X1 U150 ( .A(\block[0][83] ), .B(block_next[83]), .S0(n1611), .Y(n749) );
  OAI221X4 U151 ( .A0(n1458), .A1(n2056), .B0(n1811), .B1(n1460), .C0(n1730), 
        .Y(block_next[83]) );
  MXI4X4 U152 ( .A(\blocktag[0][19] ), .B(\blocktag[1][19] ), .C(
        \blocktag[2][19] ), .D(\blocktag[3][19] ), .S0(n1445), .S1(n1410), .Y(
        n1318) );
  OAI221X4 U153 ( .A0(n1457), .A1(n1981), .B0(n1841), .B1(n1459), .C0(n1745), 
        .Y(block_next[68]) );
  MX2X1 U154 ( .A(\block[7][77] ), .B(block_next[77]), .S0(n1503), .Y(n911) );
  MX2X1 U155 ( .A(\block[6][77] ), .B(block_next[77]), .S0(n1518), .Y(n887) );
  MX2X1 U156 ( .A(\block[5][77] ), .B(block_next[77]), .S0(n1534), .Y(n863) );
  MX2X1 U157 ( .A(\block[4][77] ), .B(block_next[77]), .S0(n1551), .Y(n839) );
  MX2X1 U158 ( .A(\block[3][77] ), .B(block_next[77]), .S0(n1568), .Y(n815) );
  MX2X1 U159 ( .A(\block[2][77] ), .B(block_next[77]), .S0(n1581), .Y(n791) );
  MX2X1 U160 ( .A(\block[1][77] ), .B(block_next[77]), .S0(n1595), .Y(n767) );
  MX2X1 U161 ( .A(\block[0][77] ), .B(block_next[77]), .S0(n1610), .Y(n743) );
  OAI221X4 U162 ( .A0(n1458), .A1(n2026), .B0(n1823), .B1(n1460), .C0(n1736), 
        .Y(block_next[77]) );
  MX2X1 U163 ( .A(\block[7][84] ), .B(block_next[84]), .S0(n1504), .Y(n918) );
  MX2X1 U164 ( .A(\block[6][84] ), .B(block_next[84]), .S0(n1519), .Y(n894) );
  MX2X1 U165 ( .A(\block[5][84] ), .B(block_next[84]), .S0(n1535), .Y(n870) );
  MX2X1 U166 ( .A(\block[4][84] ), .B(block_next[84]), .S0(n1552), .Y(n846) );
  MX2X1 U167 ( .A(\block[3][84] ), .B(block_next[84]), .S0(n1569), .Y(n822) );
  MX2X1 U168 ( .A(\block[2][84] ), .B(block_next[84]), .S0(n1582), .Y(n798) );
  MX2X1 U169 ( .A(\block[1][84] ), .B(block_next[84]), .S0(n1596), .Y(n774) );
  MX2X1 U170 ( .A(\block[0][84] ), .B(block_next[84]), .S0(n1611), .Y(n750) );
  OAI221X4 U171 ( .A0(n1457), .A1(n2061), .B0(n1809), .B1(n1460), .C0(n1729), 
        .Y(block_next[84]) );
  MX2X1 U172 ( .A(\block[7][81] ), .B(block_next[81]), .S0(n1504), .Y(n915) );
  MX2X1 U173 ( .A(\block[6][81] ), .B(block_next[81]), .S0(n1519), .Y(n891) );
  MX2X1 U174 ( .A(\block[5][81] ), .B(block_next[81]), .S0(n1535), .Y(n867) );
  MX2X1 U175 ( .A(\block[4][81] ), .B(block_next[81]), .S0(n1552), .Y(n843) );
  MX2X1 U176 ( .A(\block[3][81] ), .B(block_next[81]), .S0(n1569), .Y(n819) );
  MX2X1 U177 ( .A(\block[2][81] ), .B(block_next[81]), .S0(n1582), .Y(n795) );
  MX2X1 U178 ( .A(\block[1][81] ), .B(block_next[81]), .S0(n1596), .Y(n771) );
  MX2X1 U179 ( .A(\block[0][81] ), .B(block_next[81]), .S0(n1611), .Y(n747) );
  OAI221X4 U180 ( .A0(n1458), .A1(n2046), .B0(n1815), .B1(n1460), .C0(n1732), 
        .Y(block_next[81]) );
  MX2X1 U181 ( .A(\block[7][87] ), .B(block_next[87]), .S0(n1504), .Y(n921) );
  MX2X1 U182 ( .A(\block[6][87] ), .B(block_next[87]), .S0(n1519), .Y(n897) );
  MX2X1 U183 ( .A(\block[5][87] ), .B(block_next[87]), .S0(n1535), .Y(n873) );
  MX2X1 U184 ( .A(\block[4][87] ), .B(block_next[87]), .S0(n1552), .Y(n849) );
  MX2X1 U185 ( .A(\block[3][87] ), .B(block_next[87]), .S0(n1569), .Y(n825) );
  MX2X1 U186 ( .A(\block[2][87] ), .B(block_next[87]), .S0(n1582), .Y(n801) );
  MX2X1 U187 ( .A(\block[1][87] ), .B(block_next[87]), .S0(n1596), .Y(n777) );
  MX2X1 U188 ( .A(\block[0][87] ), .B(block_next[87]), .S0(n1611), .Y(n753) );
  OAI221X4 U189 ( .A0(n1457), .A1(n2076), .B0(n1803), .B1(n1460), .C0(n1726), 
        .Y(block_next[87]) );
  MX2X1 U190 ( .A(\block[7][82] ), .B(block_next[82]), .S0(n1504), .Y(n916) );
  MX2X1 U191 ( .A(\block[6][82] ), .B(block_next[82]), .S0(n1519), .Y(n892) );
  MX2X1 U192 ( .A(\block[5][82] ), .B(block_next[82]), .S0(n1535), .Y(n868) );
  MX2X1 U193 ( .A(\block[4][82] ), .B(block_next[82]), .S0(n1552), .Y(n844) );
  MX2X1 U194 ( .A(\block[3][82] ), .B(block_next[82]), .S0(n1569), .Y(n820) );
  MX2X1 U195 ( .A(\block[2][82] ), .B(block_next[82]), .S0(n1582), .Y(n796) );
  MX2X1 U196 ( .A(\block[1][82] ), .B(block_next[82]), .S0(n1596), .Y(n772) );
  MX2X1 U197 ( .A(\block[0][82] ), .B(block_next[82]), .S0(n1611), .Y(n748) );
  OAI221X4 U198 ( .A0(n1458), .A1(n2051), .B0(n1813), .B1(n1460), .C0(n1731), 
        .Y(block_next[82]) );
  MX2X1 U199 ( .A(\block[7][85] ), .B(block_next[85]), .S0(n1504), .Y(n919) );
  MX2X1 U200 ( .A(\block[6][85] ), .B(block_next[85]), .S0(n1519), .Y(n895) );
  MX2X1 U201 ( .A(\block[5][85] ), .B(block_next[85]), .S0(n1535), .Y(n871) );
  MX2X1 U202 ( .A(\block[4][85] ), .B(block_next[85]), .S0(n1552), .Y(n847) );
  MX2X1 U203 ( .A(\block[3][85] ), .B(block_next[85]), .S0(n1569), .Y(n823) );
  MX2X1 U204 ( .A(\block[2][85] ), .B(block_next[85]), .S0(n1582), .Y(n799) );
  MX2X1 U205 ( .A(\block[1][85] ), .B(block_next[85]), .S0(n1596), .Y(n775) );
  MX2X1 U206 ( .A(\block[0][85] ), .B(block_next[85]), .S0(n1611), .Y(n751) );
  OAI221X4 U207 ( .A0(n1457), .A1(n2066), .B0(n1807), .B1(n1460), .C0(n1728), 
        .Y(block_next[85]) );
  MX2X1 U208 ( .A(\block[7][79] ), .B(block_next[79]), .S0(n1504), .Y(n913) );
  MX2X1 U209 ( .A(\block[6][79] ), .B(block_next[79]), .S0(n1519), .Y(n889) );
  MX2X1 U210 ( .A(\block[5][79] ), .B(block_next[79]), .S0(n1535), .Y(n865) );
  MX2X1 U211 ( .A(\block[4][79] ), .B(block_next[79]), .S0(n1552), .Y(n841) );
  MX2X1 U212 ( .A(\block[3][79] ), .B(block_next[79]), .S0(n1569), .Y(n817) );
  MX2X1 U213 ( .A(\block[2][79] ), .B(block_next[79]), .S0(n1582), .Y(n793) );
  MX2X1 U214 ( .A(\block[1][79] ), .B(block_next[79]), .S0(n1596), .Y(n769) );
  MX2X1 U215 ( .A(\block[0][79] ), .B(block_next[79]), .S0(n1611), .Y(n745) );
  OAI221X4 U216 ( .A0(n1458), .A1(n2036), .B0(n1819), .B1(n1460), .C0(n1734), 
        .Y(block_next[79]) );
  NAND2X8 U217 ( .A(n12), .B(n1467), .Y(n1785) );
  NAND4X4 U218 ( .A(n1715), .B(n1461), .C(n1467), .D(n1472), .Y(n1671) );
  BUFX20 U219 ( .A(n1713), .Y(n1451) );
  INVX12 U220 ( .A(n1671), .Y(n1713) );
  CLKMX2X2 U221 ( .A(\block[0][105] ), .B(block_next[105]), .S0(n1613), .Y(
        n655) );
  BUFX12 U222 ( .A(n1713), .Y(n1450) );
  CLKMX2X2 U223 ( .A(\block[0][116] ), .B(block_next[116]), .S0(n1613), .Y(
        n665) );
  INVX8 U224 ( .A(tag[0]), .Y(n1926) );
  BUFX20 U225 ( .A(n10), .Y(n1463) );
  BUFX2 U226 ( .A(N32), .Y(n1380) );
  MXI4X2 U227 ( .A(\blocktag[4][16] ), .B(\blocktag[5][16] ), .C(
        \blocktag[6][16] ), .D(\blocktag[7][16] ), .S0(n1445), .S1(n1411), .Y(
        n1325) );
  MXI4X2 U228 ( .A(\blocktag[0][16] ), .B(\blocktag[1][16] ), .C(
        \blocktag[2][16] ), .D(\blocktag[3][16] ), .S0(n1445), .S1(n1411), .Y(
        n1324) );
  XOR2X4 U229 ( .A(n1880), .B(proc_addr[21]), .Y(n1643) );
  INVX8 U230 ( .A(tag[16]), .Y(n1880) );
  MXI4X2 U231 ( .A(\blocktag[4][12] ), .B(\blocktag[5][12] ), .C(
        \blocktag[6][12] ), .D(\blocktag[7][12] ), .S0(n1446), .S1(n1411), .Y(
        n1333) );
  MXI4X2 U232 ( .A(\blocktag[0][12] ), .B(\blocktag[1][12] ), .C(
        \blocktag[2][12] ), .D(\blocktag[3][12] ), .S0(n1446), .S1(n1411), .Y(
        n1332) );
  XOR2X4 U233 ( .A(n1890), .B(proc_addr[17]), .Y(n1642) );
  BUFX6 U234 ( .A(n1679), .Y(n15) );
  INVX8 U235 ( .A(n15), .Y(n1924) );
  INVX12 U236 ( .A(n1678), .Y(n1664) );
  NAND2XL U237 ( .A(mem_rdata[75]), .B(n1487), .Y(n1738) );
  NAND2XL U238 ( .A(mem_rdata[38]), .B(n1487), .Y(n1778) );
  NAND2XL U239 ( .A(mem_rdata[112]), .B(n1487), .Y(n1696) );
  NAND2XL U240 ( .A(mem_rdata[63]), .B(n1487), .Y(n1753) );
  NAND2XL U241 ( .A(mem_rdata[13]), .B(n1487), .Y(n1822) );
  BUFX12 U242 ( .A(n1456), .Y(n1454) );
  AND3X8 U243 ( .A(n1673), .B(proc_addr[0]), .C(n1958), .Y(n1470) );
  NAND2X4 U244 ( .A(n1673), .B(n1956), .Y(n1714) );
  MX2X1 U245 ( .A(\block[7][80] ), .B(block_next[80]), .S0(n1504), .Y(n914) );
  MX2X1 U246 ( .A(\block[6][80] ), .B(block_next[80]), .S0(n1519), .Y(n890) );
  MX2X1 U247 ( .A(\block[5][80] ), .B(block_next[80]), .S0(n1535), .Y(n866) );
  MX2X1 U248 ( .A(\block[4][80] ), .B(block_next[80]), .S0(n1552), .Y(n842) );
  MX2X1 U249 ( .A(\block[3][80] ), .B(block_next[80]), .S0(n1569), .Y(n818) );
  MX2X1 U250 ( .A(\block[2][80] ), .B(block_next[80]), .S0(n1582), .Y(n794) );
  MX2X1 U251 ( .A(\block[1][80] ), .B(block_next[80]), .S0(n1596), .Y(n770) );
  MX2X1 U252 ( .A(\block[0][80] ), .B(block_next[80]), .S0(n1611), .Y(n746) );
  OAI221X4 U253 ( .A0(n1458), .A1(n2041), .B0(n1817), .B1(n1460), .C0(n1733), 
        .Y(block_next[80]) );
  MX2X1 U254 ( .A(\block[0][67] ), .B(block_next[67]), .S0(n1610), .Y(n987) );
  MX2X1 U255 ( .A(\block[7][67] ), .B(block_next[67]), .S0(n1503), .Y(n1043)
         );
  MX2X1 U256 ( .A(\block[6][67] ), .B(block_next[67]), .S0(n1518), .Y(n1035)
         );
  MX2X1 U257 ( .A(\block[5][67] ), .B(block_next[67]), .S0(n1534), .Y(n1027)
         );
  MX2X1 U258 ( .A(\block[4][67] ), .B(block_next[67]), .S0(n1551), .Y(n1019)
         );
  MX2X1 U259 ( .A(\block[3][67] ), .B(block_next[67]), .S0(n1568), .Y(n1011)
         );
  MX2X1 U260 ( .A(\block[2][67] ), .B(block_next[67]), .S0(n1581), .Y(n1003)
         );
  MX2X1 U261 ( .A(\block[1][67] ), .B(block_next[67]), .S0(n1595), .Y(n995) );
  OAI221X4 U262 ( .A0(n1457), .A1(n1976), .B0(n1843), .B1(n1459), .C0(n1746), 
        .Y(block_next[67]) );
  CLKINVX6 U263 ( .A(n1675), .Y(n1662) );
  BUFX20 U264 ( .A(n1461), .Y(n1460) );
  BUFX20 U265 ( .A(n1461), .Y(n1459) );
  MX2X1 U266 ( .A(\block[5][71] ), .B(block_next[71]), .S0(n1534), .Y(n1031)
         );
  MX2X1 U267 ( .A(\block[7][71] ), .B(block_next[71]), .S0(n1503), .Y(n1047)
         );
  MX2X1 U268 ( .A(\block[6][71] ), .B(block_next[71]), .S0(n1518), .Y(n1039)
         );
  MX2X1 U269 ( .A(\block[4][71] ), .B(block_next[71]), .S0(n1551), .Y(n1023)
         );
  MX2X1 U270 ( .A(\block[3][71] ), .B(block_next[71]), .S0(n1568), .Y(n1015)
         );
  MX2X1 U271 ( .A(\block[2][71] ), .B(block_next[71]), .S0(n1581), .Y(n1007)
         );
  MX2X1 U272 ( .A(\block[1][71] ), .B(block_next[71]), .S0(n1595), .Y(n999) );
  MX2X1 U273 ( .A(\block[0][71] ), .B(block_next[71]), .S0(n1610), .Y(n991) );
  OAI221X4 U274 ( .A0(n1457), .A1(n1996), .B0(n1835), .B1(n1460), .C0(n1742), 
        .Y(block_next[71]) );
  BUFX12 U275 ( .A(n1924), .Y(n1473) );
  BUFX12 U276 ( .A(n1924), .Y(n1474) );
  CLKMX2X2 U277 ( .A(n1899), .B(n1898), .S0(n1481), .Y(n1900) );
  CLKMX2X2 U278 ( .A(n1860), .B(n1859), .S0(n1481), .Y(n1861) );
  OAI221X4 U279 ( .A0(n1457), .A1(n2071), .B0(n1805), .B1(n1460), .C0(n1727), 
        .Y(block_next[86]) );
  MX2X1 U280 ( .A(\block[7][86] ), .B(block_next[86]), .S0(n1504), .Y(n920) );
  BUFX16 U281 ( .A(n10), .Y(n1464) );
  BUFX20 U282 ( .A(n1751), .Y(n1461) );
  OAI221X4 U283 ( .A0(n1462), .A1(n2075), .B0(n1803), .B1(n1466), .C0(n1761), 
        .Y(block_next[55]) );
  BUFX20 U284 ( .A(n10), .Y(n1462) );
  INVX6 U285 ( .A(n1853), .Y(proc_stall) );
  BUFX20 U286 ( .A(n2125), .Y(mem_read) );
  CLKINVX8 U287 ( .A(n1668), .Y(n1715) );
  OAI211X4 U288 ( .A0(mem_ready), .A1(valid), .B0(n1667), .C0(n1948), .Y(n1668) );
  MX2X1 U289 ( .A(\block[0][99] ), .B(block_next[99]), .S0(n1612), .Y(n932) );
  MX2X1 U290 ( .A(\block[7][99] ), .B(block_next[99]), .S0(n1505), .Y(n979) );
  MX2X1 U291 ( .A(\block[6][99] ), .B(block_next[99]), .S0(n1520), .Y(n972) );
  MX2X1 U292 ( .A(\block[5][99] ), .B(block_next[99]), .S0(n1536), .Y(n965) );
  MX2X1 U293 ( .A(\block[4][99] ), .B(block_next[99]), .S0(n1553), .Y(n959) );
  MX2X1 U294 ( .A(\block[3][99] ), .B(block_next[99]), .S0(n1570), .Y(n953) );
  MX2X1 U295 ( .A(\block[2][99] ), .B(block_next[99]), .S0(n1583), .Y(n946) );
  MX2X1 U296 ( .A(\block[1][99] ), .B(block_next[99]), .S0(n1597), .Y(n939) );
  OAI221X4 U297 ( .A0(n1452), .A1(n1978), .B0(n1843), .B1(n1456), .C0(n1709), 
        .Y(block_next[99]) );
  CLKBUFX20 U298 ( .A(n36), .Y(n17) );
  BUFX6 U299 ( .A(n2116), .Y(n36) );
  OAI221X4 U300 ( .A0(n1452), .A1(n1983), .B0(n1841), .B1(n1456), .C0(n1708), 
        .Y(block_next[100]) );
  BUFX20 U301 ( .A(n1713), .Y(n1452) );
  MX2X1 U302 ( .A(\block[0][100] ), .B(block_next[100]), .S0(n1612), .Y(n933)
         );
  OAI221X4 U303 ( .A0(n1457), .A1(n2101), .B0(n1793), .B1(n1461), .C0(n1721), 
        .Y(block_next[92]) );
  OAI221X4 U304 ( .A0(n1457), .A1(n2106), .B0(n1791), .B1(n1461), .C0(n1720), 
        .Y(block_next[93]) );
  OAI221X4 U305 ( .A0(n1457), .A1(n2111), .B0(n1789), .B1(n1461), .C0(n1719), 
        .Y(block_next[94]) );
  OAI221X4 U306 ( .A0(n1457), .A1(n2117), .B0(n1787), .B1(n1461), .C0(n1718), 
        .Y(block_next[95]) );
  OAI221X4 U307 ( .A0(n1457), .A1(n2096), .B0(n1795), .B1(n1461), .C0(n1722), 
        .Y(block_next[91]) );
  OAI221X4 U308 ( .A0(n1457), .A1(n2081), .B0(n1801), .B1(n1461), .C0(n1725), 
        .Y(block_next[88]) );
  OAI221X4 U309 ( .A0(n1457), .A1(n2086), .B0(n1799), .B1(n1461), .C0(n1724), 
        .Y(block_next[89]) );
  OAI221X4 U310 ( .A0(n1457), .A1(n2091), .B0(n1797), .B1(n1461), .C0(n1723), 
        .Y(block_next[90]) );
  OAI221X4 U311 ( .A0(n1451), .A1(n2053), .B0(n1813), .B1(n1455), .C0(n1694), 
        .Y(block_next[114]) );
  OAI221X4 U312 ( .A0(n1451), .A1(n2023), .B0(n1825), .B1(n1455), .C0(n1700), 
        .Y(block_next[108]) );
  OAI221X4 U313 ( .A0(n1451), .A1(n2018), .B0(n1827), .B1(n1455), .C0(n1701), 
        .Y(block_next[107]) );
  OAI221X4 U314 ( .A0(n1451), .A1(n2028), .B0(n1823), .B1(n1455), .C0(n1699), 
        .Y(block_next[109]) );
  OAI221X4 U315 ( .A0(n1451), .A1(n2033), .B0(n1821), .B1(n1455), .C0(n1698), 
        .Y(block_next[110]) );
  OAI221X4 U316 ( .A0(n1451), .A1(n2038), .B0(n1819), .B1(n1455), .C0(n1697), 
        .Y(block_next[111]) );
  OAI221X4 U317 ( .A0(n1451), .A1(n2043), .B0(n1817), .B1(n1455), .C0(n1696), 
        .Y(block_next[112]) );
  OAI221X4 U318 ( .A0(n1451), .A1(n2048), .B0(n1815), .B1(n1455), .C0(n1695), 
        .Y(block_next[113]) );
  OAI221X4 U319 ( .A0(n1451), .A1(n2058), .B0(n1811), .B1(n1455), .C0(n1693), 
        .Y(block_next[115]) );
  INVX4 U320 ( .A(n1949), .Y(n1666) );
  INVX20 U321 ( .A(n1785), .Y(n1849) );
  INVX3 U322 ( .A(n33), .Y(n1751) );
  MX2X1 U323 ( .A(\block[1][28] ), .B(block_next[28]), .S0(n1592), .Y(n141) );
  MX2X1 U324 ( .A(\block[2][28] ), .B(block_next[28]), .S0(n1578), .Y(n153) );
  MX2X1 U325 ( .A(\block[3][28] ), .B(block_next[28]), .S0(n1565), .Y(n165) );
  MX2X1 U326 ( .A(\block[4][28] ), .B(block_next[28]), .S0(n1548), .Y(n177) );
  MX2X1 U327 ( .A(\block[5][28] ), .B(block_next[28]), .S0(n1531), .Y(n189) );
  MX2X1 U328 ( .A(\block[6][28] ), .B(block_next[28]), .S0(n1515), .Y(n201) );
  MX2X1 U329 ( .A(\block[7][28] ), .B(block_next[28]), .S0(n1500), .Y(n213) );
  NOR3X1 U330 ( .A(n1958), .B(n1854), .C(proc_addr[0]), .Y(n33) );
  CLKINVX8 U331 ( .A(n1854), .Y(n1673) );
  NAND2BX2 U332 ( .AN(n1855), .B(n1854), .Y(n1856) );
  MX2X1 U333 ( .A(\block[0][38] ), .B(block_next[38]), .S0(n1607), .Y(n581) );
  MX2X1 U334 ( .A(\block[7][38] ), .B(block_next[38]), .S0(n1500), .Y(n637) );
  MX2X1 U335 ( .A(\block[6][38] ), .B(block_next[38]), .S0(n1515), .Y(n629) );
  MX2X1 U336 ( .A(\block[5][38] ), .B(block_next[38]), .S0(n1531), .Y(n621) );
  MX2X1 U337 ( .A(\block[4][38] ), .B(block_next[38]), .S0(n1548), .Y(n613) );
  MX2X1 U338 ( .A(\block[3][38] ), .B(block_next[38]), .S0(n1565), .Y(n605) );
  MX2X1 U339 ( .A(\block[2][38] ), .B(block_next[38]), .S0(n1578), .Y(n597) );
  MX2X1 U340 ( .A(\block[1][38] ), .B(block_next[38]), .S0(n1592), .Y(n589) );
  OAI221X4 U341 ( .A0(n1464), .A1(n1990), .B0(n1837), .B1(n1465), .C0(n1778), 
        .Y(block_next[38]) );
  MX2X1 U342 ( .A(\block[0][51] ), .B(block_next[51]), .S0(n1608), .Y(n228) );
  MX2X1 U343 ( .A(\block[7][51] ), .B(block_next[51]), .S0(n1501), .Y(n389) );
  MX2X1 U344 ( .A(\block[6][51] ), .B(block_next[51]), .S0(n1516), .Y(n366) );
  MX2X1 U345 ( .A(\block[5][51] ), .B(block_next[51]), .S0(n1532), .Y(n343) );
  MX2X1 U346 ( .A(\block[4][51] ), .B(block_next[51]), .S0(n1549), .Y(n320) );
  MX2X1 U347 ( .A(\block[3][51] ), .B(block_next[51]), .S0(n1566), .Y(n297) );
  MX2X1 U348 ( .A(\block[2][51] ), .B(block_next[51]), .S0(n1579), .Y(n274) );
  MX2X1 U349 ( .A(\block[1][51] ), .B(block_next[51]), .S0(n1593), .Y(n251) );
  OAI221X4 U350 ( .A0(n1463), .A1(n2055), .B0(n1811), .B1(n1466), .C0(n1765), 
        .Y(block_next[51]) );
  INVX8 U351 ( .A(n1717), .Y(n1750) );
  NAND3BX4 U352 ( .AN(n1468), .B(n1752), .C(n1471), .Y(n1717) );
  NAND2X2 U353 ( .A(n1666), .B(valid), .Y(n1670) );
  NOR2X8 U354 ( .A(n65), .B(n66), .Y(n61) );
  NOR2X2 U355 ( .A(n64), .B(n1919), .Y(n66) );
  NOR2X8 U356 ( .A(n59), .B(n60), .Y(n55) );
  NOR2X2 U357 ( .A(n58), .B(n1874), .Y(n60) );
  NOR2X8 U358 ( .A(n53), .B(n54), .Y(n50) );
  NOR2X2 U359 ( .A(n52), .B(n1859), .Y(n54) );
  NAND2X4 U360 ( .A(n1956), .B(n1955), .Y(n2121) );
  BUFX3 U361 ( .A(n2121), .Y(n1492) );
  BUFX20 U362 ( .A(n1491), .Y(n1494) );
  MX2X1 U363 ( .A(\block[0][31] ), .B(block_next[31]), .S0(n1607), .Y(n132) );
  MX2X1 U364 ( .A(\block[7][31] ), .B(block_next[31]), .S0(n1500), .Y(n216) );
  MX2X1 U365 ( .A(\block[6][31] ), .B(block_next[31]), .S0(n1515), .Y(n204) );
  MX2X1 U366 ( .A(\block[5][31] ), .B(block_next[31]), .S0(n1531), .Y(n192) );
  MX2X1 U367 ( .A(\block[4][31] ), .B(block_next[31]), .S0(n1548), .Y(n180) );
  MX2X1 U368 ( .A(\block[3][31] ), .B(block_next[31]), .S0(n1565), .Y(n168) );
  MX2X1 U369 ( .A(\block[2][31] ), .B(block_next[31]), .S0(n1578), .Y(n156) );
  MX2X1 U370 ( .A(\block[1][31] ), .B(block_next[31]), .S0(n1592), .Y(n144) );
  OAI221X4 U371 ( .A0(n1471), .A1(n1787), .B0(n1849), .B1(n2122), .C0(n1786), 
        .Y(block_next[31]) );
  MX2X1 U372 ( .A(\block[0][29] ), .B(block_next[29]), .S0(n1607), .Y(n130) );
  MX2X1 U373 ( .A(\block[7][29] ), .B(block_next[29]), .S0(n1500), .Y(n214) );
  MX2X1 U374 ( .A(\block[6][29] ), .B(block_next[29]), .S0(n1515), .Y(n202) );
  MX2X1 U375 ( .A(\block[5][29] ), .B(block_next[29]), .S0(n1531), .Y(n190) );
  MX2X1 U376 ( .A(\block[4][29] ), .B(block_next[29]), .S0(n1548), .Y(n178) );
  MX2X1 U377 ( .A(\block[3][29] ), .B(block_next[29]), .S0(n1565), .Y(n166) );
  MX2X1 U378 ( .A(\block[2][29] ), .B(block_next[29]), .S0(n1578), .Y(n154) );
  MX2X1 U379 ( .A(\block[1][29] ), .B(block_next[29]), .S0(n1592), .Y(n142) );
  OAI221X4 U380 ( .A0(n1471), .A1(n1791), .B0(n1849), .B1(n2109), .C0(n1790), 
        .Y(block_next[29]) );
  MX2X1 U381 ( .A(\block[0][30] ), .B(block_next[30]), .S0(n1607), .Y(n131) );
  MX2X1 U382 ( .A(\block[7][30] ), .B(block_next[30]), .S0(n1500), .Y(n215) );
  MX2X1 U383 ( .A(\block[6][30] ), .B(block_next[30]), .S0(n1515), .Y(n203) );
  MX2X1 U384 ( .A(\block[5][30] ), .B(block_next[30]), .S0(n1531), .Y(n191) );
  MX2X1 U385 ( .A(\block[4][30] ), .B(block_next[30]), .S0(n1548), .Y(n179) );
  MX2X1 U386 ( .A(\block[3][30] ), .B(block_next[30]), .S0(n1565), .Y(n167) );
  MX2X1 U387 ( .A(\block[2][30] ), .B(block_next[30]), .S0(n1578), .Y(n155) );
  MX2X1 U388 ( .A(\block[1][30] ), .B(block_next[30]), .S0(n1592), .Y(n143) );
  OAI221X4 U389 ( .A0(n1471), .A1(n1789), .B0(n1849), .B1(n2114), .C0(n1788), 
        .Y(block_next[30]) );
  MX2X1 U390 ( .A(\block[0][25] ), .B(block_next[25]), .S0(n1606), .Y(n126) );
  MX2X1 U391 ( .A(\block[7][25] ), .B(block_next[25]), .S0(n1499), .Y(n210) );
  MX2X1 U392 ( .A(\block[6][25] ), .B(block_next[25]), .S0(n1514), .Y(n198) );
  MX2X1 U393 ( .A(\block[5][25] ), .B(block_next[25]), .S0(n1530), .Y(n186) );
  MX2X1 U394 ( .A(\block[4][25] ), .B(block_next[25]), .S0(n1547), .Y(n174) );
  MX2X1 U395 ( .A(\block[3][25] ), .B(block_next[25]), .S0(n1564), .Y(n162) );
  MX2X1 U396 ( .A(\block[2][25] ), .B(block_next[25]), .S0(n1577), .Y(n150) );
  MX2X1 U397 ( .A(\block[1][25] ), .B(block_next[25]), .S0(n1591), .Y(n138) );
  OAI221X4 U398 ( .A0(n1471), .A1(n1799), .B0(n1849), .B1(n2089), .C0(n1798), 
        .Y(block_next[25]) );
  OAI221X4 U399 ( .A0(n1451), .A1(n2008), .B0(n1831), .B1(n1455), .C0(n1703), 
        .Y(block_next[105]) );
  BUFX12 U400 ( .A(n1453), .Y(n1455) );
  MX2X1 U401 ( .A(\block[0][26] ), .B(block_next[26]), .S0(n1606), .Y(n127) );
  MX2X1 U402 ( .A(\block[7][26] ), .B(block_next[26]), .S0(n1499), .Y(n211) );
  MX2X1 U403 ( .A(\block[6][26] ), .B(block_next[26]), .S0(n1514), .Y(n199) );
  MX2X1 U404 ( .A(\block[5][26] ), .B(block_next[26]), .S0(n1530), .Y(n187) );
  MX2X1 U405 ( .A(\block[4][26] ), .B(block_next[26]), .S0(n1547), .Y(n175) );
  MX2X1 U406 ( .A(\block[3][26] ), .B(block_next[26]), .S0(n1564), .Y(n163) );
  MX2X1 U407 ( .A(\block[2][26] ), .B(block_next[26]), .S0(n1577), .Y(n151) );
  MX2X1 U408 ( .A(\block[1][26] ), .B(block_next[26]), .S0(n1591), .Y(n139) );
  OAI221X4 U409 ( .A0(n1471), .A1(n1797), .B0(n1849), .B1(n2094), .C0(n1796), 
        .Y(block_next[26]) );
  MX2X1 U410 ( .A(\block[0][23] ), .B(block_next[23]), .S0(n1606), .Y(n124) );
  MX2X1 U411 ( .A(\block[7][23] ), .B(block_next[23]), .S0(n1499), .Y(n208) );
  MX2X1 U412 ( .A(\block[6][23] ), .B(block_next[23]), .S0(n1514), .Y(n196) );
  MX2X1 U413 ( .A(\block[5][23] ), .B(block_next[23]), .S0(n1530), .Y(n184) );
  MX2X1 U414 ( .A(\block[4][23] ), .B(block_next[23]), .S0(n1547), .Y(n172) );
  MX2X1 U415 ( .A(\block[3][23] ), .B(block_next[23]), .S0(n1564), .Y(n160) );
  MX2X1 U416 ( .A(\block[2][23] ), .B(block_next[23]), .S0(n1577), .Y(n148) );
  MX2X1 U417 ( .A(\block[1][23] ), .B(block_next[23]), .S0(n1591), .Y(n136) );
  OAI221X4 U418 ( .A0(n1471), .A1(n1803), .B0(n1849), .B1(n2079), .C0(n1802), 
        .Y(block_next[23]) );
  MX2X1 U419 ( .A(\block[0][24] ), .B(block_next[24]), .S0(n1606), .Y(n125) );
  MX2X1 U420 ( .A(\block[7][24] ), .B(block_next[24]), .S0(n1499), .Y(n209) );
  MX2X1 U421 ( .A(\block[6][24] ), .B(block_next[24]), .S0(n1514), .Y(n197) );
  MX2X1 U422 ( .A(\block[5][24] ), .B(block_next[24]), .S0(n1530), .Y(n185) );
  MX2X1 U423 ( .A(\block[4][24] ), .B(block_next[24]), .S0(n1547), .Y(n173) );
  MX2X1 U424 ( .A(\block[3][24] ), .B(block_next[24]), .S0(n1564), .Y(n161) );
  MX2X1 U425 ( .A(\block[2][24] ), .B(block_next[24]), .S0(n1577), .Y(n149) );
  MX2X1 U426 ( .A(\block[1][24] ), .B(block_next[24]), .S0(n1591), .Y(n137) );
  OAI221X4 U427 ( .A0(n1471), .A1(n1801), .B0(n1849), .B1(n2084), .C0(n1800), 
        .Y(block_next[24]) );
  MX2X1 U428 ( .A(\block[0][21] ), .B(block_next[21]), .S0(n1606), .Y(n122) );
  MX2X1 U429 ( .A(\block[7][21] ), .B(block_next[21]), .S0(n1499), .Y(n206) );
  MX2X1 U430 ( .A(\block[6][21] ), .B(block_next[21]), .S0(n1514), .Y(n194) );
  MX2X1 U431 ( .A(\block[5][21] ), .B(block_next[21]), .S0(n1530), .Y(n182) );
  MX2X1 U432 ( .A(\block[4][21] ), .B(block_next[21]), .S0(n1547), .Y(n170) );
  MX2X1 U433 ( .A(\block[3][21] ), .B(block_next[21]), .S0(n1564), .Y(n158) );
  MX2X1 U434 ( .A(\block[2][21] ), .B(block_next[21]), .S0(n1577), .Y(n146) );
  MX2X1 U435 ( .A(\block[1][21] ), .B(block_next[21]), .S0(n1591), .Y(n134) );
  OAI221X4 U436 ( .A0(n1471), .A1(n1807), .B0(n1849), .B1(n2069), .C0(n1806), 
        .Y(block_next[21]) );
  MX2X1 U437 ( .A(\block[0][22] ), .B(block_next[22]), .S0(n1606), .Y(n123) );
  MX2X1 U438 ( .A(\block[7][22] ), .B(block_next[22]), .S0(n1499), .Y(n207) );
  MX2X1 U439 ( .A(\block[6][22] ), .B(block_next[22]), .S0(n1514), .Y(n195) );
  MX2X1 U440 ( .A(\block[5][22] ), .B(block_next[22]), .S0(n1530), .Y(n183) );
  MX2X1 U441 ( .A(\block[4][22] ), .B(block_next[22]), .S0(n1547), .Y(n171) );
  MX2X1 U442 ( .A(\block[3][22] ), .B(block_next[22]), .S0(n1564), .Y(n159) );
  MX2X1 U443 ( .A(\block[2][22] ), .B(block_next[22]), .S0(n1577), .Y(n147) );
  MX2X1 U444 ( .A(\block[1][22] ), .B(block_next[22]), .S0(n1591), .Y(n135) );
  OAI221X4 U445 ( .A0(n1471), .A1(n1805), .B0(n1849), .B1(n2074), .C0(n1804), 
        .Y(block_next[22]) );
  MX2X1 U446 ( .A(\block[0][20] ), .B(block_next[20]), .S0(n1606), .Y(n121) );
  MX2X1 U447 ( .A(\block[7][20] ), .B(block_next[20]), .S0(n1499), .Y(n205) );
  MX2X1 U448 ( .A(\block[6][20] ), .B(block_next[20]), .S0(n1514), .Y(n193) );
  MX2X1 U449 ( .A(\block[5][20] ), .B(block_next[20]), .S0(n1530), .Y(n181) );
  MX2X1 U450 ( .A(\block[4][20] ), .B(block_next[20]), .S0(n1547), .Y(n169) );
  MX2X1 U451 ( .A(\block[3][20] ), .B(block_next[20]), .S0(n1564), .Y(n157) );
  MX2X1 U452 ( .A(\block[2][20] ), .B(block_next[20]), .S0(n1577), .Y(n145) );
  MX2X1 U453 ( .A(\block[1][20] ), .B(block_next[20]), .S0(n1591), .Y(n133) );
  OAI221X4 U454 ( .A0(n1471), .A1(n1809), .B0(n1849), .B1(n2064), .C0(n1808), 
        .Y(block_next[20]) );
  MXI4X1 U455 ( .A(\blocktag[4][13] ), .B(\blocktag[5][13] ), .C(
        \blocktag[6][13] ), .D(\blocktag[7][13] ), .S0(n1445), .S1(n1411), .Y(
        n1331) );
  MXI4X1 U456 ( .A(\blocktag[0][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[3][13] ), .S0(n1445), .S1(n1411), .Y(
        n1330) );
  XOR2X4 U457 ( .A(n1887), .B(proc_addr[18]), .Y(n1660) );
  CLKINVX4 U458 ( .A(n1676), .Y(n1663) );
  NAND4X8 U459 ( .A(n1654), .B(n1653), .C(n1652), .D(n1651), .Y(n1676) );
  NAND3BXL U460 ( .AN(mem_ready), .B(proc_stall), .C(n1950), .Y(n1953) );
  NAND2X2 U461 ( .A(n1951), .B(n1953), .Y(n1952) );
  XOR2X4 U462 ( .A(tag[9]), .B(n1898), .Y(n1634) );
  CLKINVX1 U463 ( .A(proc_addr[14]), .Y(n1898) );
  INVX4 U464 ( .A(n1670), .Y(n1665) );
  XOR2X4 U465 ( .A(n9), .B(proc_addr[20]), .Y(n1661) );
  MXI4X1 U466 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n1445), .S1(n1411), .Y(
        n1327) );
  MXI4X1 U467 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n1445), .S1(n1411), .Y(
        n1326) );
  BUFX20 U468 ( .A(n1491), .Y(n1493) );
  XOR2X2 U469 ( .A(n1914), .B(proc_addr[9]), .Y(n1637) );
  MXI4X2 U470 ( .A(\blocktag[4][4] ), .B(\blocktag[5][4] ), .C(
        \blocktag[6][4] ), .D(\blocktag[7][4] ), .S0(n1447), .S1(n1413), .Y(
        n1349) );
  MXI4X4 U471 ( .A(\blocktag[0][4] ), .B(\blocktag[1][4] ), .C(
        \blocktag[2][4] ), .D(\blocktag[3][4] ), .S0(n1447), .S1(n1413), .Y(
        n1348) );
  INVX4 U472 ( .A(n2137), .Y(n18) );
  CLKINVX20 U473 ( .A(n18), .Y(mem_addr[1]) );
  AND2XL U474 ( .A(N32), .B(n1952), .Y(n2137) );
  INVX8 U475 ( .A(n2139), .Y(n20) );
  CLKINVX20 U476 ( .A(n20), .Y(mem_wdata[108]) );
  CLKAND2X4 U477 ( .A(n1624), .B(blockdata[108]), .Y(n2139) );
  INVX4 U478 ( .A(n2138), .Y(n22) );
  CLKINVX20 U479 ( .A(n22), .Y(mem_addr[0]) );
  AND2XL U480 ( .A(n1618), .B(n1952), .Y(n2138) );
  NAND2X8 U481 ( .A(n1945), .B(n1628), .Y(n1943) );
  INVX20 U486 ( .A(proc_addr[1]), .Y(n1958) );
  OAI221X4 U487 ( .A0(n1452), .A1(n1973), .B0(n1845), .B1(n1714), .C0(n1710), 
        .Y(block_next[98]) );
  INVX3 U488 ( .A(blockdata[98]), .Y(n1973) );
  MX2X1 U489 ( .A(\block[0][96] ), .B(block_next[96]), .S0(n1612), .Y(n930) );
  MX2X1 U490 ( .A(\block[1][96] ), .B(block_next[96]), .S0(n1597), .Y(n937) );
  MX2X1 U491 ( .A(\block[2][96] ), .B(block_next[96]), .S0(n1583), .Y(n944) );
  MX2X1 U492 ( .A(\block[3][96] ), .B(block_next[96]), .S0(n1570), .Y(n951) );
  MX2X1 U493 ( .A(\block[4][96] ), .B(block_next[96]), .S0(n1553), .Y(n958) );
  MX2X1 U494 ( .A(\block[5][96] ), .B(block_next[96]), .S0(n1536), .Y(n964) );
  OAI221X4 U495 ( .A0(n1452), .A1(n1963), .B0(n1850), .B1(n1456), .C0(n1712), 
        .Y(block_next[96]) );
  INVXL U496 ( .A(n1908), .Y(n28) );
  INVX4 U497 ( .A(n2123), .Y(n30) );
  INVX20 U498 ( .A(n30), .Y(n31) );
  MX2XL U499 ( .A(n1308), .B(n1309), .S0(n1373), .Y(n32) );
  INVX1 U500 ( .A(n32), .Y(n34) );
  MXI4X4 U501 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n1445), .S1(n1411), .Y(
        n1329) );
  MXI4X4 U502 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n1445), .S1(n1411), .Y(
        n1328) );
  OAI221X4 U503 ( .A0(n1471), .A1(n1813), .B0(n1849), .B1(n2054), .C0(n1812), 
        .Y(n35) );
  BUFX16 U504 ( .A(n1473), .Y(n1488) );
  BUFX20 U505 ( .A(n1474), .Y(n1490) );
  BUFX20 U506 ( .A(n1474), .Y(n1489) );
  BUFX16 U507 ( .A(n1924), .Y(n1487) );
  BUFX16 U508 ( .A(n1473), .Y(n1486) );
  BUFX20 U509 ( .A(n1488), .Y(n1480) );
  BUFX20 U510 ( .A(n1489), .Y(n1478) );
  BUFX20 U511 ( .A(n1490), .Y(n1476) );
  BUFX20 U512 ( .A(n1490), .Y(n1475) );
  BUFX20 U513 ( .A(n1489), .Y(n1477) );
  BUFX12 U514 ( .A(n1473), .Y(n1484) );
  BUFX12 U515 ( .A(n1474), .Y(n1483) );
  BUFX20 U516 ( .A(n1487), .Y(n1482) );
  BUFX16 U517 ( .A(n1487), .Y(n1481) );
  BUFX16 U518 ( .A(n1486), .Y(n1485) );
  OAI221X4 U519 ( .A0(n1452), .A1(n1998), .B0(n1835), .B1(n1456), .C0(n1705), 
        .Y(block_next[103]) );
  NAND2XL U520 ( .A(mem_rdata[103]), .B(n1477), .Y(n1705) );
  OAI221X4 U521 ( .A0(n1458), .A1(n1971), .B0(n1845), .B1(n1459), .C0(n1747), 
        .Y(block_next[66]) );
  NAND2XL U522 ( .A(mem_rdata[66]), .B(n1484), .Y(n1747) );
  OAI221X4 U523 ( .A0(n1452), .A1(n1988), .B0(n1839), .B1(n1456), .C0(n1707), 
        .Y(block_next[101]) );
  NAND2XL U524 ( .A(mem_rdata[101]), .B(n1474), .Y(n1707) );
  OAI221X4 U525 ( .A0(n1457), .A1(n1986), .B0(n1839), .B1(n1459), .C0(n1744), 
        .Y(block_next[69]) );
  NAND2XL U526 ( .A(mem_rdata[69]), .B(n1477), .Y(n1744) );
  OAI221X4 U527 ( .A0(n1452), .A1(n1993), .B0(n1837), .B1(n1456), .C0(n1706), 
        .Y(block_next[102]) );
  NAND2XL U528 ( .A(mem_rdata[102]), .B(n1473), .Y(n1706) );
  OAI221X4 U529 ( .A0(n1458), .A1(n1991), .B0(n1837), .B1(n1459), .C0(n1743), 
        .Y(block_next[70]) );
  NAND2XL U530 ( .A(mem_rdata[70]), .B(n1475), .Y(n1743) );
  MXI4XL U531 ( .A(\blocktag[2][21] ), .B(\blocktag[3][21] ), .C(
        \blocktag[0][21] ), .D(\blocktag[1][21] ), .S0(n120), .S1(n1620), .Y(
        n1314) );
  OAI221X4 U532 ( .A0(n1457), .A1(n1966), .B0(n1847), .B1(n1459), .C0(n1748), 
        .Y(block_next[65]) );
  NAND2XL U533 ( .A(mem_rdata[65]), .B(n1487), .Y(n1748) );
  OAI221X4 U534 ( .A0(n1450), .A1(n2098), .B0(n1795), .B1(n1454), .C0(n1685), 
        .Y(block_next[123]) );
  NAND2XL U535 ( .A(mem_rdata[123]), .B(n1485), .Y(n1685) );
  OAI221X4 U536 ( .A0(n1450), .A1(n2120), .B0(n1787), .B1(n1454), .C0(n1680), 
        .Y(block_next[127]) );
  NAND2XL U537 ( .A(mem_rdata[127]), .B(n1477), .Y(n1680) );
  OAI221X4 U538 ( .A0(n1450), .A1(n2108), .B0(n1791), .B1(n1454), .C0(n1683), 
        .Y(block_next[125]) );
  NAND2XL U539 ( .A(mem_rdata[125]), .B(n1484), .Y(n1683) );
  OAI221X4 U540 ( .A0(n1463), .A1(n2045), .B0(n1815), .B1(n1466), .C0(n1767), 
        .Y(block_next[49]) );
  OAI221X4 U541 ( .A0(n1462), .A1(n2065), .B0(n1807), .B1(n1466), .C0(n1763), 
        .Y(block_next[53]) );
  NAND2X2 U542 ( .A(mem_rdata[53]), .B(n1489), .Y(n1763) );
  OAI221X4 U543 ( .A0(n1464), .A1(n1975), .B0(n1843), .B1(n1465), .C0(n1781), 
        .Y(block_next[35]) );
  OAI221X4 U544 ( .A0(n1463), .A1(n2050), .B0(n1813), .B1(n1466), .C0(n1766), 
        .Y(block_next[50]) );
  OAI221X4 U545 ( .A0(n1462), .A1(n2070), .B0(n1805), .B1(n1466), .C0(n1762), 
        .Y(block_next[54]) );
  NAND2X2 U546 ( .A(mem_rdata[54]), .B(n1488), .Y(n1762) );
  OAI221X4 U547 ( .A0(n1464), .A1(n1980), .B0(n1841), .B1(n1465), .C0(n1780), 
        .Y(block_next[36]) );
  OAI221X4 U548 ( .A0(n1463), .A1(n2035), .B0(n1819), .B1(n1466), .C0(n1769), 
        .Y(block_next[47]) );
  OAI221X4 U549 ( .A0(n1462), .A1(n2060), .B0(n1809), .B1(n1466), .C0(n1764), 
        .Y(block_next[52]) );
  OAI221X4 U550 ( .A0(n1450), .A1(n2113), .B0(n1789), .B1(n1454), .C0(n1682), 
        .Y(block_next[126]) );
  NAND2XL U551 ( .A(mem_rdata[126]), .B(n1483), .Y(n1682) );
  OAI221X4 U552 ( .A0(n1463), .A1(n2040), .B0(n1817), .B1(n1466), .C0(n1768), 
        .Y(block_next[48]) );
  OAI221X4 U553 ( .A0(n1464), .A1(n1965), .B0(n1847), .B1(n1465), .C0(n1783), 
        .Y(block_next[33]) );
  OAI221X4 U554 ( .A0(n1463), .A1(n2025), .B0(n1823), .B1(n1466), .C0(n1771), 
        .Y(block_next[45]) );
  OAI221X4 U555 ( .A0(n1464), .A1(n1970), .B0(n1845), .B1(n1465), .C0(n1782), 
        .Y(block_next[34]) );
  OAI221X4 U556 ( .A0(n1450), .A1(n2103), .B0(n1793), .B1(n1454), .C0(n1684), 
        .Y(block_next[124]) );
  NAND2XL U557 ( .A(mem_rdata[124]), .B(n1475), .Y(n1684) );
  OAI221X4 U558 ( .A0(n1463), .A1(n2030), .B0(n1821), .B1(n1466), .C0(n1770), 
        .Y(block_next[46]) );
  CLKINVX8 U559 ( .A(block_next[7]), .Y(n37) );
  INVX16 U560 ( .A(n37), .Y(n38) );
  OAI221X4 U561 ( .A0(n1463), .A1(n2015), .B0(n1827), .B1(n1465), .C0(n1773), 
        .Y(block_next[43]) );
  OAI221X4 U562 ( .A0(n1464), .A1(n1960), .B0(n1850), .B1(n1465), .C0(n1784), 
        .Y(block_next[32]) );
  OAI221X4 U563 ( .A0(n1463), .A1(n2020), .B0(n1825), .B1(n1465), .C0(n1772), 
        .Y(block_next[44]) );
  MX2X1 U564 ( .A(\block[0][5] ), .B(block_next[5]), .S0(n1605), .Y(n516) );
  MX2X1 U565 ( .A(\block[1][5] ), .B(block_next[5]), .S0(n1590), .Y(n524) );
  MX2X1 U566 ( .A(\block[2][5] ), .B(block_next[5]), .S0(n1576), .Y(n532) );
  MX2X1 U567 ( .A(\block[3][5] ), .B(block_next[5]), .S0(n1563), .Y(n540) );
  MX2X1 U568 ( .A(\block[4][5] ), .B(block_next[5]), .S0(n1546), .Y(n548) );
  MX2X1 U569 ( .A(\block[5][5] ), .B(block_next[5]), .S0(n1529), .Y(n556) );
  OAI221X4 U570 ( .A0(n1472), .A1(n1839), .B0(n1849), .B1(n1989), .C0(n1838), 
        .Y(block_next[5]) );
  OAI221X4 U571 ( .A0(n1450), .A1(n2088), .B0(n1799), .B1(n1454), .C0(n1687), 
        .Y(block_next[121]) );
  NAND2XL U572 ( .A(mem_rdata[121]), .B(n1478), .Y(n1687) );
  OAI221X4 U573 ( .A0(n1464), .A1(n1995), .B0(n1835), .B1(n1466), .C0(n1777), 
        .Y(block_next[39]) );
  INVX12 U574 ( .A(n1468), .Y(n1466) );
  OAI221X4 U575 ( .A0(n1463), .A1(n2005), .B0(n1831), .B1(n1465), .C0(n1775), 
        .Y(block_next[41]) );
  OAI221X4 U576 ( .A0(n1458), .A1(n1961), .B0(n1850), .B1(n1459), .C0(n1749), 
        .Y(block_next[64]) );
  NAND2XL U577 ( .A(mem_rdata[64]), .B(n1480), .Y(n1749) );
  OAI221X4 U578 ( .A0(n1463), .A1(n2010), .B0(n1829), .B1(n1465), .C0(n1774), 
        .Y(block_next[42]) );
  BUFX6 U579 ( .A(block_next[40]), .Y(n39) );
  OAI221XL U580 ( .A0(n1463), .A1(n2000), .B0(n1833), .B1(n1465), .C0(n1776), 
        .Y(block_next[40]) );
  OAI221X4 U581 ( .A0(n1450), .A1(n2093), .B0(n1797), .B1(n1454), .C0(n1686), 
        .Y(block_next[122]) );
  NAND2XL U582 ( .A(mem_rdata[122]), .B(n1476), .Y(n1686) );
  XOR2X4 U583 ( .A(tag[24]), .B(n40), .Y(n1650) );
  OAI221X4 U584 ( .A0(n1471), .A1(n1819), .B0(n1849), .B1(n2039), .C0(n1818), 
        .Y(block_next[15]) );
  NAND2XL U585 ( .A(mem_rdata[15]), .B(n1483), .Y(n1818) );
  OAI221X4 U586 ( .A0(n1450), .A1(n2078), .B0(n1803), .B1(n1454), .C0(n1689), 
        .Y(block_next[119]) );
  NAND2XL U587 ( .A(mem_rdata[119]), .B(n1482), .Y(n1689) );
  OAI221X4 U588 ( .A0(n1471), .A1(n1817), .B0(n1849), .B1(n2044), .C0(n1816), 
        .Y(block_next[16]) );
  MX2X1 U589 ( .A(\block[0][6] ), .B(block_next[6]), .S0(n1605), .Y(n517) );
  MX2X1 U590 ( .A(\block[1][6] ), .B(block_next[6]), .S0(n1590), .Y(n525) );
  MX2X1 U591 ( .A(\block[2][6] ), .B(block_next[6]), .S0(n1576), .Y(n533) );
  MX2X1 U592 ( .A(\block[3][6] ), .B(block_next[6]), .S0(n1563), .Y(n541) );
  MX2X1 U593 ( .A(\block[4][6] ), .B(block_next[6]), .S0(n1546), .Y(n549) );
  MX2X1 U594 ( .A(\block[5][6] ), .B(block_next[6]), .S0(n1529), .Y(n557) );
  OAI221X4 U595 ( .A0(n1472), .A1(n1837), .B0(n1849), .B1(n1994), .C0(n1836), 
        .Y(block_next[6]) );
  MX2X1 U596 ( .A(\block[0][13] ), .B(block_next[13]), .S0(n1605), .Y(n404) );
  MX2X1 U597 ( .A(\block[1][13] ), .B(block_next[13]), .S0(n1590), .Y(n413) );
  MX2X1 U598 ( .A(\block[2][13] ), .B(block_next[13]), .S0(n1576), .Y(n422) );
  MX2X1 U599 ( .A(\block[3][13] ), .B(block_next[13]), .S0(n1563), .Y(n432) );
  MX2X1 U600 ( .A(\block[4][13] ), .B(block_next[13]), .S0(n1546), .Y(n442) );
  MX2X1 U601 ( .A(\block[5][13] ), .B(block_next[13]), .S0(n1529), .Y(n452) );
  OAI221X4 U602 ( .A0(n1471), .A1(n1823), .B0(n1849), .B1(n2029), .C0(n1822), 
        .Y(block_next[13]) );
  OAI221X4 U603 ( .A0(n1450), .A1(n2083), .B0(n1801), .B1(n1454), .C0(n1688), 
        .Y(block_next[120]) );
  NAND2XL U604 ( .A(mem_rdata[120]), .B(n1474), .Y(n1688) );
  MX2X1 U605 ( .A(\block[0][3] ), .B(block_next[3]), .S0(n1605), .Y(n514) );
  MX2X1 U606 ( .A(\block[1][3] ), .B(block_next[3]), .S0(n1590), .Y(n522) );
  MX2X1 U607 ( .A(\block[2][3] ), .B(block_next[3]), .S0(n1576), .Y(n530) );
  MX2X1 U608 ( .A(\block[3][3] ), .B(block_next[3]), .S0(n1563), .Y(n538) );
  MX2X1 U609 ( .A(\block[4][3] ), .B(block_next[3]), .S0(n1546), .Y(n546) );
  MX2X1 U610 ( .A(\block[5][3] ), .B(block_next[3]), .S0(n1529), .Y(n554) );
  OAI221X4 U611 ( .A0(n1472), .A1(n1843), .B0(n1849), .B1(n1979), .C0(n1842), 
        .Y(block_next[3]) );
  OAI221X4 U612 ( .A0(n1472), .A1(n1821), .B0(n1849), .B1(n2034), .C0(n1820), 
        .Y(block_next[14]) );
  MX2X1 U613 ( .A(\block[0][11] ), .B(block_next[11]), .S0(n1605), .Y(n402) );
  MX2X1 U614 ( .A(\block[1][11] ), .B(block_next[11]), .S0(n1590), .Y(n411) );
  MX2X1 U615 ( .A(\block[2][11] ), .B(block_next[11]), .S0(n1576), .Y(n420) );
  MX2X1 U616 ( .A(\block[3][11] ), .B(block_next[11]), .S0(n1563), .Y(n430) );
  MX2X1 U617 ( .A(\block[4][11] ), .B(block_next[11]), .S0(n1546), .Y(n440) );
  MX2X1 U618 ( .A(\block[5][11] ), .B(block_next[11]), .S0(n1529), .Y(n450) );
  OAI221X4 U619 ( .A0(n1472), .A1(n1827), .B0(n1849), .B1(n2019), .C0(n1826), 
        .Y(block_next[11]) );
  MX2X1 U620 ( .A(\block[0][4] ), .B(block_next[4]), .S0(n1605), .Y(n515) );
  MX2X1 U621 ( .A(\block[1][4] ), .B(block_next[4]), .S0(n1590), .Y(n523) );
  MX2X1 U622 ( .A(\block[2][4] ), .B(block_next[4]), .S0(n1576), .Y(n531) );
  MX2X1 U623 ( .A(\block[3][4] ), .B(block_next[4]), .S0(n1563), .Y(n539) );
  MX2X1 U624 ( .A(\block[4][4] ), .B(block_next[4]), .S0(n1546), .Y(n547) );
  MX2X1 U625 ( .A(\block[5][4] ), .B(block_next[4]), .S0(n1529), .Y(n555) );
  OAI221X4 U626 ( .A0(n1472), .A1(n1841), .B0(n1849), .B1(n1984), .C0(n1840), 
        .Y(block_next[4]) );
  AO22X1 U627 ( .A0(proc_addr[10]), .A1(mem_read), .B0(tag[5]), .B1(mem_write), 
        .Y(mem_addr[8]) );
  AO22X1 U628 ( .A0(proc_addr[17]), .A1(mem_read), .B0(tag[12]), .B1(mem_write), .Y(mem_addr[15]) );
  INVXL U629 ( .A(proc_stall), .Y(n45) );
  AO22X1 U630 ( .A0(proc_addr[21]), .A1(mem_read), .B0(tag[16]), .B1(mem_write), .Y(mem_addr[19]) );
  BUFX20 U631 ( .A(block_next[12]), .Y(n46) );
  OAI221X4 U632 ( .A0(n1472), .A1(n1825), .B0(n1849), .B1(n2024), .C0(n1824), 
        .Y(block_next[12]) );
  BUFX20 U633 ( .A(block_next[1]), .Y(n47) );
  OAI221X4 U634 ( .A0(n1472), .A1(n1847), .B0(n1849), .B1(n1969), .C0(n1846), 
        .Y(block_next[1]) );
  BUFX20 U635 ( .A(block_next[10]), .Y(n48) );
  OAI221X4 U636 ( .A0(n1472), .A1(n1829), .B0(n1849), .B1(n2014), .C0(n1828), 
        .Y(block_next[10]) );
  OAI221X2 U637 ( .A0(n31), .A1(n2099), .B0(n1495), .B1(n2098), .C0(n2097), 
        .Y(proc_rdata[27]) );
  AND2XL U638 ( .A(n1625), .B(blockdata[37]), .Y(mem_wdata[37]) );
  BUFX20 U639 ( .A(block_next[19]), .Y(n49) );
  OAI221X4 U640 ( .A0(n1471), .A1(n1811), .B0(n1849), .B1(n2059), .C0(n1810), 
        .Y(block_next[19]) );
  AND2XL U641 ( .A(n1625), .B(blockdata[46]), .Y(mem_wdata[46]) );
  AND2XL U642 ( .A(n1625), .B(blockdata[47]), .Y(mem_wdata[47]) );
  AND2XL U643 ( .A(n1625), .B(blockdata[48]), .Y(mem_wdata[48]) );
  AND2XL U644 ( .A(n1625), .B(blockdata[49]), .Y(mem_wdata[49]) );
  AND2XL U645 ( .A(n1626), .B(blockdata[7]), .Y(mem_wdata[7]) );
  AND2XL U646 ( .A(n1625), .B(blockdata[50]), .Y(mem_wdata[50]) );
  AND2XL U647 ( .A(n1626), .B(blockdata[8]), .Y(mem_wdata[8]) );
  AND2XL U648 ( .A(n1625), .B(blockdata[51]), .Y(mem_wdata[51]) );
  AND2XL U649 ( .A(n1626), .B(blockdata[9]), .Y(mem_wdata[9]) );
  AND2XL U650 ( .A(n1625), .B(blockdata[52]), .Y(mem_wdata[52]) );
  AND2XL U651 ( .A(n1624), .B(blockdata[83]), .Y(mem_wdata[83]) );
  AND2XL U652 ( .A(n1626), .B(blockdata[10]), .Y(mem_wdata[10]) );
  AND2XL U653 ( .A(n1625), .B(blockdata[53]), .Y(mem_wdata[53]) );
  AND2XL U654 ( .A(n1624), .B(blockdata[84]), .Y(mem_wdata[84]) );
  AND2XL U655 ( .A(n1626), .B(blockdata[11]), .Y(mem_wdata[11]) );
  AND2XL U656 ( .A(n1625), .B(blockdata[54]), .Y(mem_wdata[54]) );
  AND2XL U657 ( .A(n1624), .B(blockdata[85]), .Y(mem_wdata[85]) );
  AND2XL U658 ( .A(n1626), .B(blockdata[12]), .Y(mem_wdata[12]) );
  AND2XL U659 ( .A(n1625), .B(blockdata[55]), .Y(mem_wdata[55]) );
  AND2XL U660 ( .A(n1624), .B(blockdata[86]), .Y(mem_wdata[86]) );
  AND2XL U661 ( .A(n1626), .B(blockdata[13]), .Y(mem_wdata[13]) );
  AND2XL U662 ( .A(n1625), .B(blockdata[56]), .Y(mem_wdata[56]) );
  AND2XL U663 ( .A(n1624), .B(blockdata[87]), .Y(mem_wdata[87]) );
  AND2XL U664 ( .A(n1626), .B(blockdata[14]), .Y(mem_wdata[14]) );
  AND2XL U665 ( .A(n1625), .B(blockdata[57]), .Y(mem_wdata[57]) );
  AND2XL U666 ( .A(n1624), .B(blockdata[88]), .Y(mem_wdata[88]) );
  AND2XL U667 ( .A(n1626), .B(blockdata[15]), .Y(mem_wdata[15]) );
  AND2XL U668 ( .A(n1625), .B(blockdata[58]), .Y(mem_wdata[58]) );
  AND2XL U669 ( .A(n1624), .B(blockdata[89]), .Y(mem_wdata[89]) );
  AND2XL U670 ( .A(n1626), .B(blockdata[16]), .Y(mem_wdata[16]) );
  AND2XL U671 ( .A(n1625), .B(blockdata[59]), .Y(mem_wdata[59]) );
  AND2XL U672 ( .A(n1624), .B(blockdata[90]), .Y(mem_wdata[90]) );
  AND2XL U673 ( .A(n1626), .B(blockdata[17]), .Y(mem_wdata[17]) );
  AND2XL U674 ( .A(n1625), .B(blockdata[60]), .Y(mem_wdata[60]) );
  AND2XL U675 ( .A(n1624), .B(blockdata[91]), .Y(mem_wdata[91]) );
  AND2XL U676 ( .A(n1626), .B(blockdata[18]), .Y(mem_wdata[18]) );
  AND2XL U677 ( .A(n1625), .B(blockdata[61]), .Y(mem_wdata[61]) );
  OAI221X1 U678 ( .A0(n31), .A1(n1984), .B0(n1493), .B1(n1983), .C0(n1982), 
        .Y(proc_rdata[4]) );
  AND2XL U679 ( .A(n1624), .B(blockdata[92]), .Y(mem_wdata[92]) );
  AND2XL U680 ( .A(n1626), .B(blockdata[19]), .Y(mem_wdata[19]) );
  AND2XL U681 ( .A(n1625), .B(blockdata[62]), .Y(mem_wdata[62]) );
  AND2XL U682 ( .A(n1624), .B(blockdata[93]), .Y(mem_wdata[93]) );
  AND2XL U683 ( .A(n1626), .B(blockdata[20]), .Y(mem_wdata[20]) );
  AND2XL U684 ( .A(n1625), .B(blockdata[63]), .Y(mem_wdata[63]) );
  AND2XL U685 ( .A(n1624), .B(blockdata[94]), .Y(mem_wdata[94]) );
  AND2XL U686 ( .A(n1626), .B(blockdata[21]), .Y(mem_wdata[21]) );
  AND2XL U687 ( .A(n1625), .B(blockdata[64]), .Y(mem_wdata[64]) );
  AND2XL U688 ( .A(n1624), .B(blockdata[95]), .Y(mem_wdata[95]) );
  AND2XL U689 ( .A(n1626), .B(blockdata[22]), .Y(mem_wdata[22]) );
  AND2XL U690 ( .A(n1625), .B(blockdata[65]), .Y(mem_wdata[65]) );
  AND2XL U691 ( .A(n1624), .B(blockdata[96]), .Y(mem_wdata[96]) );
  AND2XL U692 ( .A(n1626), .B(blockdata[23]), .Y(mem_wdata[23]) );
  AND2XL U693 ( .A(n1625), .B(blockdata[66]), .Y(mem_wdata[66]) );
  AND2XL U694 ( .A(n1624), .B(blockdata[97]), .Y(mem_wdata[97]) );
  AND2XL U695 ( .A(n1626), .B(blockdata[24]), .Y(mem_wdata[24]) );
  AND2XL U696 ( .A(n1625), .B(blockdata[67]), .Y(mem_wdata[67]) );
  AND2XL U697 ( .A(n1624), .B(blockdata[98]), .Y(mem_wdata[98]) );
  AND2XL U698 ( .A(n1626), .B(blockdata[25]), .Y(mem_wdata[25]) );
  AND2XL U699 ( .A(n1625), .B(blockdata[68]), .Y(mem_wdata[68]) );
  AND2XL U700 ( .A(n1624), .B(blockdata[99]), .Y(mem_wdata[99]) );
  AND2XL U701 ( .A(n1626), .B(blockdata[26]), .Y(mem_wdata[26]) );
  AND2XL U702 ( .A(n1625), .B(blockdata[69]), .Y(mem_wdata[69]) );
  AND2XL U703 ( .A(n1624), .B(blockdata[100]), .Y(mem_wdata[100]) );
  AND2XL U704 ( .A(n1626), .B(blockdata[27]), .Y(mem_wdata[27]) );
  AND2XL U705 ( .A(n1625), .B(blockdata[70]), .Y(mem_wdata[70]) );
  AND2XL U706 ( .A(n1624), .B(blockdata[101]), .Y(mem_wdata[101]) );
  AND2XL U707 ( .A(n1626), .B(blockdata[28]), .Y(mem_wdata[28]) );
  AND2XL U708 ( .A(n1624), .B(blockdata[102]), .Y(mem_wdata[102]) );
  AND2XL U709 ( .A(n1626), .B(blockdata[29]), .Y(mem_wdata[29]) );
  AND2XL U710 ( .A(n1624), .B(blockdata[103]), .Y(mem_wdata[103]) );
  AND2XL U711 ( .A(n1626), .B(blockdata[30]), .Y(mem_wdata[30]) );
  AND2XL U712 ( .A(n1624), .B(blockdata[104]), .Y(mem_wdata[104]) );
  AND2XL U713 ( .A(n1626), .B(blockdata[31]), .Y(mem_wdata[31]) );
  AND2XL U714 ( .A(n1624), .B(blockdata[105]), .Y(mem_wdata[105]) );
  AND2XL U715 ( .A(n1624), .B(blockdata[106]), .Y(mem_wdata[106]) );
  AND2XL U716 ( .A(n1624), .B(blockdata[107]), .Y(mem_wdata[107]) );
  OAI221X2 U717 ( .A0(n31), .A1(n2049), .B0(n1494), .B1(n2048), .C0(n2047), 
        .Y(proc_rdata[17]) );
  OAI221X1 U718 ( .A0(n31), .A1(n2044), .B0(n1494), .B1(n2043), .C0(n2042), 
        .Y(proc_rdata[16]) );
  OAI221X1 U719 ( .A0(n31), .A1(n2064), .B0(n1494), .B1(n2063), .C0(n2062), 
        .Y(proc_rdata[20]) );
  OAI221X1 U720 ( .A0(n31), .A1(n2029), .B0(n1494), .B1(n2028), .C0(n2027), 
        .Y(proc_rdata[13]) );
  OAI221X1 U721 ( .A0(n31), .A1(n2074), .B0(n1494), .B1(n2073), .C0(n2072), 
        .Y(proc_rdata[22]) );
  OAI221X1 U722 ( .A0(n31), .A1(n2039), .B0(n1494), .B1(n2038), .C0(n2037), 
        .Y(proc_rdata[15]) );
  OAI221X1 U723 ( .A0(n31), .A1(n2034), .B0(n1494), .B1(n2033), .C0(n2032), 
        .Y(proc_rdata[14]) );
  OAI221X1 U724 ( .A0(n31), .A1(n2069), .B0(n1494), .B1(n2068), .C0(n2067), 
        .Y(proc_rdata[21]) );
  OAI221X1 U725 ( .A0(n31), .A1(n2079), .B0(n1494), .B1(n2078), .C0(n2077), 
        .Y(proc_rdata[23]) );
  OAI221X1 U726 ( .A0(n31), .A1(n2054), .B0(n1494), .B1(n2053), .C0(n2052), 
        .Y(proc_rdata[18]) );
  OAI221X2 U727 ( .A0(n31), .A1(n2059), .B0(n1494), .B1(n2058), .C0(n2057), 
        .Y(proc_rdata[19]) );
  OAI221X2 U728 ( .A0(n31), .A1(n2024), .B0(n1494), .B1(n2023), .C0(n2022), 
        .Y(proc_rdata[12]) );
  OAI221X1 U729 ( .A0(n31), .A1(n1979), .B0(n1493), .B1(n1978), .C0(n1977), 
        .Y(proc_rdata[3]) );
  OAI221X1 U730 ( .A0(n31), .A1(n1974), .B0(n1493), .B1(n1973), .C0(n1972), 
        .Y(proc_rdata[2]) );
  OAI221X1 U731 ( .A0(n31), .A1(n2004), .B0(n1493), .B1(n2003), .C0(n2002), 
        .Y(proc_rdata[8]) );
  OAI221X1 U732 ( .A0(n31), .A1(n1964), .B0(n1493), .B1(n1963), .C0(n1962), 
        .Y(proc_rdata[0]) );
  OAI221X1 U733 ( .A0(n31), .A1(n2014), .B0(n1493), .B1(n2013), .C0(n2012), 
        .Y(proc_rdata[10]) );
  OAI221X1 U734 ( .A0(n31), .A1(n2019), .B0(n1493), .B1(n2018), .C0(n2017), 
        .Y(proc_rdata[11]) );
  OAI221X1 U735 ( .A0(n31), .A1(n2009), .B0(n1493), .B1(n2008), .C0(n2007), 
        .Y(proc_rdata[9]) );
  OAI221X2 U736 ( .A0(n31), .A1(n1994), .B0(n1493), .B1(n1993), .C0(n1992), 
        .Y(proc_rdata[6]) );
  OAI221X2 U737 ( .A0(n31), .A1(n1989), .B0(n1493), .B1(n1988), .C0(n1987), 
        .Y(proc_rdata[5]) );
  BUFX20 U738 ( .A(N33), .Y(n1362) );
  NAND4X8 U739 ( .A(n1658), .B(n1660), .C(n1659), .D(n1661), .Y(n1675) );
  OA22XL U740 ( .A0(n29), .A1(n1996), .B0(n17), .B1(n1995), .Y(n1997) );
  NAND4BX2 U741 ( .AN(n1950), .B(n1949), .C(n1948), .D(n1947), .Y(n1951) );
  INVX8 U742 ( .A(tag[12]), .Y(n1890) );
  OA21X4 U743 ( .A0(n45), .A1(n1947), .B0(dirty), .Y(n1855) );
  BUFX16 U744 ( .A(n1714), .Y(n1453) );
  OAI221X4 U745 ( .A0(n1472), .A1(n1845), .B0(n1849), .B1(n1974), .C0(n1844), 
        .Y(block_next[2]) );
  CLKXOR2X2 U746 ( .A(n1908), .B(proc_addr[11]), .Y(n1638) );
  MXI4X2 U747 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(
        \blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n1447), .S1(n1413), .Y(
        n1352) );
  MXI4X2 U748 ( .A(\blocktag[4][2] ), .B(\blocktag[5][2] ), .C(
        \blocktag[6][2] ), .D(\blocktag[7][2] ), .S0(n1447), .S1(n1413), .Y(
        n1353) );
  INVX6 U749 ( .A(tag[22]), .Y(n1863) );
  INVX20 U750 ( .A(n1468), .Y(n1467) );
  BUFX12 U751 ( .A(n1470), .Y(n1468) );
  OAI221X4 U752 ( .A0(n1452), .A1(n1968), .B0(n1847), .B1(n1456), .C0(n1711), 
        .Y(block_next[97]) );
  NAND2X2 U753 ( .A(mem_rdata[97]), .B(n1490), .Y(n1711) );
  MXI4X2 U754 ( .A(\blocktag[0][20] ), .B(\blocktag[1][20] ), .C(
        \blocktag[2][20] ), .D(\blocktag[3][20] ), .S0(n1444), .S1(n1410), .Y(
        n1316) );
  MXI4X2 U755 ( .A(\blocktag[4][23] ), .B(\blocktag[5][23] ), .C(
        \blocktag[6][23] ), .D(\blocktag[7][23] ), .S0(n1444), .S1(n1410), .Y(
        n1311) );
  MXI4X2 U756 ( .A(\blocktag[0][23] ), .B(\blocktag[1][23] ), .C(
        \blocktag[2][23] ), .D(\blocktag[3][23] ), .S0(n1444), .S1(n1410), .Y(
        n1310) );
  MXI4X1 U757 ( .A(\blocktag[4][21] ), .B(\blocktag[5][21] ), .C(
        \blocktag[6][21] ), .D(\blocktag[7][21] ), .S0(n1444), .S1(n1410), .Y(
        n1315) );
  NAND2X4 U758 ( .A(n1638), .B(n1637), .Y(n1639) );
  AND3X8 U759 ( .A(n1650), .B(n1649), .C(n1648), .Y(n1651) );
  MXI4X2 U760 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n1444), .S1(n1410), .Y(
        n1317) );
  INVX1 U761 ( .A(tag[2]), .Y(n63) );
  NAND3X8 U762 ( .A(n1636), .B(n1635), .C(n1634), .Y(n1640) );
  BUFX16 U763 ( .A(n1419), .Y(n1420) );
  MXI4X1 U764 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n1446), .S1(n1412), .Y(
        n1335) );
  MXI4X2 U765 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(
        \blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n1447), .S1(n1413), .Y(
        n1347) );
  MXI4X2 U766 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(
        \blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n1447), .S1(n1413), .Y(
        n1346) );
  CLKXOR2X2 U767 ( .A(n1872), .B(proc_addr[24]), .Y(n1653) );
  AND3X8 U768 ( .A(n1643), .B(n1642), .C(n1641), .Y(n1644) );
  XOR2X4 U769 ( .A(proc_addr[8]), .B(tag[3]), .Y(n1631) );
  MXI4X1 U770 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n1446), .S1(n1412), .Y(
        n1334) );
  MXI4X2 U771 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(
        \blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n1446), .S1(n1412), .Y(
        n1339) );
  OAI221X4 U772 ( .A0(n1462), .A1(n2080), .B0(n1801), .B1(n1467), .C0(n1760), 
        .Y(block_next[56]) );
  OAI221X4 U773 ( .A0(n1462), .A1(n2085), .B0(n1799), .B1(n1467), .C0(n1759), 
        .Y(block_next[57]) );
  OAI221X4 U774 ( .A0(n1462), .A1(n2090), .B0(n1797), .B1(n1467), .C0(n1758), 
        .Y(block_next[58]) );
  OAI221X4 U775 ( .A0(n1462), .A1(n2095), .B0(n1795), .B1(n1467), .C0(n1757), 
        .Y(block_next[59]) );
  OAI221X4 U776 ( .A0(n1462), .A1(n2100), .B0(n1793), .B1(n1467), .C0(n1756), 
        .Y(block_next[60]) );
  OAI221X4 U777 ( .A0(n1462), .A1(n2105), .B0(n1791), .B1(n1467), .C0(n1755), 
        .Y(block_next[61]) );
  OAI221X4 U778 ( .A0(n1462), .A1(n2110), .B0(n1789), .B1(n1467), .C0(n1754), 
        .Y(block_next[62]) );
  OAI221X4 U779 ( .A0(n1462), .A1(n2115), .B0(n1787), .B1(n1467), .C0(n1753), 
        .Y(block_next[63]) );
  CLKBUFX2 U780 ( .A(n1470), .Y(n1469) );
  MX2X1 U781 ( .A(\block[0][0] ), .B(block_next[0]), .S0(n1604), .Y(n511) );
  MX2X1 U782 ( .A(\block[1][0] ), .B(block_next[0]), .S0(n1589), .Y(n519) );
  MX2X1 U783 ( .A(\block[2][0] ), .B(block_next[0]), .S0(n1575), .Y(n527) );
  OAI221X4 U784 ( .A0(n1471), .A1(n1850), .B0(n1849), .B1(n1964), .C0(n1848), 
        .Y(block_next[0]) );
  MX2X1 U785 ( .A(\block[0][117] ), .B(block_next[117]), .S0(n1613), .Y(n666)
         );
  OAI221X4 U786 ( .A0(n1450), .A1(n2068), .B0(n1807), .B1(n1454), .C0(n1691), 
        .Y(block_next[117]) );
  BUFX20 U787 ( .A(n1381), .Y(n1383) );
  BUFX20 U788 ( .A(N32), .Y(n1381) );
  BUFX20 U789 ( .A(n1449), .Y(n1419) );
  BUFX20 U790 ( .A(n1419), .Y(n1421) );
  OAI221X4 U791 ( .A0(n1471), .A1(n1815), .B0(n1849), .B1(n2049), .C0(n1814), 
        .Y(block_next[17]) );
  MX2X1 U792 ( .A(\block[7][18] ), .B(block_next[18]), .S0(n1499), .Y(n509) );
  OAI221X4 U793 ( .A0(n1472), .A1(n1813), .B0(n1849), .B1(n2054), .C0(n1812), 
        .Y(block_next[18]) );
  NOR2X8 U794 ( .A(n1640), .B(n1639), .Y(n1674) );
  MXI4X4 U795 ( .A(\blocktag[0][6] ), .B(\blocktag[1][6] ), .C(
        \blocktag[2][6] ), .D(\blocktag[3][6] ), .S0(n1447), .S1(n1412), .Y(
        n1344) );
  MXI4X2 U796 ( .A(\blocktag[4][17] ), .B(\blocktag[5][17] ), .C(
        \blocktag[6][17] ), .D(\blocktag[7][17] ), .S0(n1445), .S1(n1411), .Y(
        n1323) );
  BUFX20 U797 ( .A(n1622), .Y(n1625) );
  MXI4X4 U798 ( .A(\blocktag[4][6] ), .B(\blocktag[5][6] ), .C(
        \blocktag[6][6] ), .D(\blocktag[7][6] ), .S0(n1446), .S1(n1412), .Y(
        n1345) );
  BUFX20 U799 ( .A(n1420), .Y(n1446) );
  OAI221X4 U800 ( .A0(n1471), .A1(n1795), .B0(n1849), .B1(n2099), .C0(n1794), 
        .Y(block_next[27]) );
  MX2X1 U801 ( .A(\block[0][118] ), .B(block_next[118]), .S0(n1613), .Y(n667)
         );
  OAI221X4 U802 ( .A0(n1450), .A1(n2073), .B0(n1805), .B1(n1454), .C0(n1690), 
        .Y(block_next[118]) );
  MX2X1 U803 ( .A(\block[0][28] ), .B(block_next[28]), .S0(n1607), .Y(n129) );
  OAI221X4 U804 ( .A0(n1471), .A1(n1793), .B0(n1849), .B1(n2104), .C0(n1792), 
        .Y(block_next[28]) );
  MXI4X1 U805 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(
        \blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n1446), .S1(n1412), .Y(
        n1338) );
  INVX1 U806 ( .A(tag[14]), .Y(n87) );
  MXI4X2 U807 ( .A(\blocktag[4][1] ), .B(\blocktag[5][1] ), .C(
        \blocktag[6][1] ), .D(\blocktag[7][1] ), .S0(n1447), .S1(n1413), .Y(
        n1355) );
  XOR2X4 U808 ( .A(n1922), .B(proc_addr[6]), .Y(n1659) );
  INVX6 U809 ( .A(tag[1]), .Y(n1922) );
  MXI4X2 U810 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(
        \blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n1447), .S1(n1413), .Y(
        n1354) );
  AND2XL U811 ( .A(N33), .B(n1952), .Y(mem_addr[2]) );
  NAND4X8 U812 ( .A(n1647), .B(n1646), .C(n1645), .D(n1644), .Y(n1678) );
  NAND4X4 U813 ( .A(n1674), .B(n1664), .C(n1663), .D(n1662), .Y(n1949) );
  BUFX20 U814 ( .A(n1851), .Y(n1471) );
  OAI221X4 U815 ( .A0(n1458), .A1(n2031), .B0(n1821), .B1(n1460), .C0(n1735), 
        .Y(block_next[78]) );
  BUFX20 U816 ( .A(n1750), .Y(n1458) );
  BUFX20 U817 ( .A(n1622), .Y(n1624) );
  OAI221X1 U818 ( .A0(n31), .A1(n1969), .B0(n1493), .B1(n1968), .C0(n1967), 
        .Y(proc_rdata[1]) );
  INVX4 U819 ( .A(tag[7]), .Y(n1905) );
  MXI2X4 U820 ( .A(n1342), .B(n1343), .S0(n1375), .Y(tag[7]) );
  BUFX20 U821 ( .A(n1383), .Y(n1410) );
  BUFX20 U822 ( .A(n1362), .Y(n1374) );
  MXI2X4 U823 ( .A(n1314), .B(n1315), .S0(n1374), .Y(tag[21]) );
  CLKBUFX20 U824 ( .A(n1622), .Y(mem_write) );
  AO22XL U825 ( .A0(proc_addr[22]), .A1(mem_read), .B0(tag[17]), .B1(mem_write), .Y(mem_addr[20]) );
  AO22XL U826 ( .A0(proc_addr[26]), .A1(mem_read), .B0(tag[21]), .B1(mem_write), .Y(mem_addr[24]) );
  MXI4X2 U827 ( .A(\blocktag[4][3] ), .B(\blocktag[5][3] ), .C(
        \blocktag[6][3] ), .D(\blocktag[7][3] ), .S0(n1447), .S1(n1413), .Y(
        n1351) );
  MXI4X2 U828 ( .A(\blocktag[0][3] ), .B(\blocktag[1][3] ), .C(
        \blocktag[2][3] ), .D(\blocktag[3][3] ), .S0(n1447), .S1(n1413), .Y(
        n1350) );
  BUFX20 U829 ( .A(n1382), .Y(n1413) );
  MXI4X4 U830 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n1444), .S1(n1416), .Y(
        n1309) );
  BUFX20 U831 ( .A(n1384), .Y(n1409) );
  BUFX20 U832 ( .A(n1618), .Y(n1449) );
  BUFX20 U833 ( .A(n120), .Y(n1443) );
  NAND2X4 U834 ( .A(dirty), .B(valid), .Y(n1950) );
  BUFX20 U835 ( .A(n1420), .Y(n1447) );
  BUFX20 U836 ( .A(n1382), .Y(n1412) );
  BUFX20 U837 ( .A(n1851), .Y(n1472) );
  OAI221X4 U838 ( .A0(n1451), .A1(n2013), .B0(n1829), .B1(n1455), .C0(n1702), 
        .Y(block_next[106]) );
  MXI4X4 U839 ( .A(\blocktag[0][24] ), .B(\blocktag[1][24] ), .C(
        \blocktag[2][24] ), .D(\blocktag[3][24] ), .S0(n1444), .S1(n1409), .Y(
        n1308) );
  BUFX20 U840 ( .A(n1421), .Y(n1444) );
  OAI221X4 U841 ( .A0(n1450), .A1(n2063), .B0(n1809), .B1(n1454), .C0(n1692), 
        .Y(block_next[116]) );
  MXI2X4 U842 ( .A(n1318), .B(n1319), .S0(n1374), .Y(tag[19]) );
  MXI4X4 U843 ( .A(\blocktag[4][19] ), .B(\blocktag[5][19] ), .C(
        \blocktag[6][19] ), .D(\blocktag[7][19] ), .S0(n1444), .S1(n1410), .Y(
        n1319) );
  NOR2X8 U844 ( .A(n1633), .B(n1632), .Y(n1635) );
  MXI2X4 U845 ( .A(n1352), .B(n1353), .S0(n1375), .Y(tag[2]) );
  MXI2X4 U846 ( .A(n1348), .B(n1349), .S0(n1375), .Y(tag[4]) );
  MXI4X2 U847 ( .A(\blocktag[4][18] ), .B(\blocktag[5][18] ), .C(
        \blocktag[6][18] ), .D(\blocktag[7][18] ), .S0(n1445), .S1(n1410), .Y(
        n1321) );
  BUFX20 U848 ( .A(n1421), .Y(n1445) );
  MXI2X4 U849 ( .A(n1320), .B(n1321), .S0(n1374), .Y(tag[18]) );
  MXI4X2 U850 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n1445), .S1(n1410), .Y(
        n1320) );
  BUFX8 U851 ( .A(N33), .Y(n1361) );
  NAND3BX4 U852 ( .AN(n1670), .B(proc_write), .C(n1669), .Y(n1854) );
  OAI221X4 U853 ( .A0(n1451), .A1(n2003), .B0(n1833), .B1(n1455), .C0(n1704), 
        .Y(block_next[104]) );
  MXI2X4 U854 ( .A(n1310), .B(n1311), .S0(n1374), .Y(tag[23]) );
  BUFX20 U855 ( .A(n1622), .Y(n1626) );
  BUFX12 U856 ( .A(n2126), .Y(n1622) );
  CLKAND2X12 U857 ( .A(n1626), .B(blockdata[32]), .Y(mem_wdata[32]) );
  BUFX20 U858 ( .A(n1362), .Y(n1373) );
  MXI2X2 U859 ( .A(n1306), .B(n1307), .S0(n1373), .Y(dirty) );
  MXI2X4 U860 ( .A(n1328), .B(n1329), .S0(n1374), .Y(tag[14]) );
  BUFX20 U861 ( .A(n1383), .Y(n1411) );
  XOR2X4 U862 ( .A(n1877), .B(proc_addr[22]), .Y(n1656) );
  INVX20 U863 ( .A(n1619), .Y(n1618) );
  MXI2X4 U864 ( .A(n1316), .B(n1317), .S0(n1374), .Y(tag[20]) );
  INVX4 U865 ( .A(blockdata[6]), .Y(n1994) );
  MXI2X1 U866 ( .A(n1290), .B(n1291), .S0(n1373), .Y(blockdata[6]) );
  INVX4 U867 ( .A(blockdata[5]), .Y(n1989) );
  MXI2X1 U868 ( .A(n1292), .B(n1293), .S0(n1373), .Y(blockdata[5]) );
  INVX4 U869 ( .A(blockdata[4]), .Y(n1984) );
  MXI2X1 U870 ( .A(n1294), .B(n1295), .S0(n1373), .Y(blockdata[4]) );
  CLKAND2X12 U871 ( .A(n1624), .B(blockdata[6]), .Y(mem_wdata[6]) );
  INVX4 U872 ( .A(blockdata[3]), .Y(n1979) );
  MXI2X1 U873 ( .A(n1296), .B(n1297), .S0(n1373), .Y(blockdata[3]) );
  CLKAND2X12 U874 ( .A(n1624), .B(blockdata[5]), .Y(mem_wdata[5]) );
  INVX4 U875 ( .A(blockdata[2]), .Y(n1974) );
  MXI2X1 U876 ( .A(n1298), .B(n1299), .S0(n1373), .Y(blockdata[2]) );
  CLKAND2X12 U877 ( .A(n1624), .B(blockdata[4]), .Y(mem_wdata[4]) );
  MXI2X1 U878 ( .A(n1300), .B(n1301), .S0(n1373), .Y(blockdata[1]) );
  INVX20 U879 ( .A(n50), .Y(mem_addr[26]) );
  CLKINVX1 U880 ( .A(mem_write), .Y(n51) );
  INVXL U881 ( .A(mem_read), .Y(n52) );
  NOR2X2 U882 ( .A(n51), .B(n1860), .Y(n53) );
  INVX20 U883 ( .A(n55), .Y(mem_addr[21]) );
  CLKINVX1 U884 ( .A(mem_write), .Y(n56) );
  CLKINVX1 U885 ( .A(tag[18]), .Y(n57) );
  INVXL U886 ( .A(mem_read), .Y(n58) );
  NOR2X2 U887 ( .A(n56), .B(n57), .Y(n59) );
  INVX20 U888 ( .A(n61), .Y(mem_addr[5]) );
  CLKINVX1 U889 ( .A(mem_write), .Y(n62) );
  INVXL U890 ( .A(mem_read), .Y(n64) );
  NOR2X2 U891 ( .A(n62), .B(n63), .Y(n65) );
  CLKAND2X12 U892 ( .A(n1624), .B(blockdata[3]), .Y(mem_wdata[3]) );
  CLKINVX6 U893 ( .A(n2127), .Y(n67) );
  INVX20 U894 ( .A(n67), .Y(mem_addr[27]) );
  AO22X1 U895 ( .A0(proc_addr[29]), .A1(mem_read), .B0(n34), .B1(mem_write), 
        .Y(n2127) );
  CLKINVX6 U896 ( .A(n2128), .Y(n69) );
  INVX20 U897 ( .A(n69), .Y(mem_addr[25]) );
  AO22X1 U898 ( .A0(proc_addr[27]), .A1(mem_read), .B0(tag[22]), .B1(mem_write), .Y(n2128) );
  INVX20 U899 ( .A(n71), .Y(mem_addr[23]) );
  NOR2X2 U900 ( .A(n72), .B(n1869), .Y(n73) );
  NOR2X1 U901 ( .A(n109), .B(n1868), .Y(n74) );
  INVX20 U902 ( .A(n75), .Y(mem_addr[22]) );
  INVXL U903 ( .A(mem_read), .Y(n77) );
  NOR2X2 U904 ( .A(n76), .B(n1872), .Y(n78) );
  NOR2X1 U905 ( .A(n77), .B(n1871), .Y(n79) );
  INVX20 U906 ( .A(n80), .Y(mem_addr[18]) );
  NOR2X2 U907 ( .A(n81), .B(n9), .Y(n83) );
  NOR2X1 U908 ( .A(n82), .B(n1882), .Y(n84) );
  INVX20 U909 ( .A(n85), .Y(mem_addr[17]) );
  NOR2X2 U910 ( .A(n86), .B(n87), .Y(n89) );
  NOR2X1 U911 ( .A(n82), .B(n88), .Y(n90) );
  CLKINVX6 U912 ( .A(n2129), .Y(n91) );
  INVX20 U913 ( .A(n91), .Y(mem_addr[14]) );
  AO22X1 U914 ( .A0(proc_addr[16]), .A1(mem_read), .B0(tag[11]), .B1(mem_write), .Y(n2129) );
  CLKINVX6 U915 ( .A(n2130), .Y(n93) );
  INVX20 U916 ( .A(n93), .Y(mem_addr[13]) );
  AO22X1 U917 ( .A0(proc_addr[15]), .A1(mem_read), .B0(tag[10]), .B1(mem_write), .Y(n2130) );
  CLKINVX6 U918 ( .A(n2131), .Y(n95) );
  INVX20 U919 ( .A(n95), .Y(mem_addr[12]) );
  AO22X1 U920 ( .A0(proc_addr[14]), .A1(mem_read), .B0(tag[9]), .B1(mem_write), 
        .Y(n2131) );
  CLKINVX6 U921 ( .A(n2132), .Y(n97) );
  INVX20 U922 ( .A(n97), .Y(mem_addr[11]) );
  AO22X1 U923 ( .A0(proc_addr[13]), .A1(mem_read), .B0(tag[8]), .B1(mem_write), 
        .Y(n2132) );
  INVX20 U924 ( .A(n99), .Y(mem_addr[10]) );
  INVXL U925 ( .A(tag[7]), .Y(n101) );
  INVXL U926 ( .A(mem_read), .Y(n102) );
  NOR2X2 U927 ( .A(n100), .B(n101), .Y(n103) );
  NOR2X1 U928 ( .A(n102), .B(n1904), .Y(n104) );
  CLKINVX6 U929 ( .A(n2133), .Y(n105) );
  INVX20 U930 ( .A(n105), .Y(mem_addr[9]) );
  AO22X1 U931 ( .A0(proc_addr[11]), .A1(mem_read), .B0(n28), .B1(mem_write), 
        .Y(n2133) );
  INVX20 U932 ( .A(n107), .Y(mem_addr[7]) );
  NOR2X2 U933 ( .A(n108), .B(n1914), .Y(n110) );
  NOR2X1 U934 ( .A(n109), .B(n1913), .Y(n111) );
  CLKINVX6 U935 ( .A(n2134), .Y(n112) );
  INVX20 U936 ( .A(n112), .Y(mem_addr[6]) );
  AO22X1 U937 ( .A0(proc_addr[8]), .A1(mem_read), .B0(tag[3]), .B1(mem_write), 
        .Y(n2134) );
  CLKINVX6 U938 ( .A(n2135), .Y(n114) );
  INVX20 U939 ( .A(n114), .Y(mem_addr[4]) );
  AO22X1 U940 ( .A0(proc_addr[6]), .A1(mem_read), .B0(tag[1]), .B1(mem_write), 
        .Y(n2135) );
  CLKINVX6 U941 ( .A(n2136), .Y(n116) );
  INVX20 U942 ( .A(n116), .Y(mem_addr[3]) );
  AO22X1 U943 ( .A0(proc_addr[5]), .A1(mem_read), .B0(tag[0]), .B1(mem_write), 
        .Y(n2136) );
  CLKAND2X12 U944 ( .A(n1624), .B(blockdata[2]), .Y(mem_wdata[2]) );
  CLKAND2X12 U945 ( .A(n1624), .B(blockdata[1]), .Y(mem_wdata[1]) );
  INVXL U946 ( .A(proc_write), .Y(n1954) );
  CLKBUFX4 U947 ( .A(n1418), .Y(n1430) );
  BUFX4 U948 ( .A(n1510), .Y(n1523) );
  BUFX4 U949 ( .A(n1418), .Y(n1423) );
  BUFX4 U950 ( .A(n1378), .Y(n1387) );
  BUFX2 U951 ( .A(n1379), .Y(n1386) );
  CLKBUFX3 U952 ( .A(n1417), .Y(n1424) );
  BUFX4 U953 ( .A(n1615), .Y(n1616) );
  CLKBUFX2 U954 ( .A(n2), .Y(n1587) );
  CLKBUFX2 U955 ( .A(n4), .Y(n1617) );
  CLKBUFX2 U956 ( .A(n1), .Y(n1601) );
  CLKBUFX4 U957 ( .A(n1377), .Y(n1389) );
  CLKBUFX2 U958 ( .A(n1543), .Y(n1558) );
  INVXL U959 ( .A(n1620), .Y(n118) );
  INVXL U960 ( .A(n1619), .Y(n119) );
  MXI4XL U961 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n1443), .S1(n1409), .Y(n1304) );
  MXI4XL U962 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n1443), .S1(n1409), .Y(n1305) );
  XOR2X4 U963 ( .A(n1860), .B(proc_addr[28]), .Y(n1648) );
  MXI4XL U964 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n1437), .S1(n1402), .Y(n1224) );
  MXI4XL U965 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n1437), .S1(n1402), .Y(n1225) );
  BUFX20 U966 ( .A(n1453), .Y(n1456) );
  NOR2X8 U967 ( .A(n1631), .B(n1630), .Y(n1636) );
  NAND3BX4 U968 ( .AN(proc_addr[0]), .B(n1673), .C(n1958), .Y(n1851) );
  INVX3 U969 ( .A(blockdata[0]), .Y(n1964) );
  INVX3 U970 ( .A(blockdata[38]), .Y(n1990) );
  INVX3 U971 ( .A(blockdata[33]), .Y(n1965) );
  INVX3 U972 ( .A(blockdata[34]), .Y(n1970) );
  INVX3 U973 ( .A(blockdata[35]), .Y(n1975) );
  INVX3 U974 ( .A(blockdata[36]), .Y(n1980) );
  INVX3 U975 ( .A(blockdata[40]), .Y(n2000) );
  INVX3 U976 ( .A(blockdata[41]), .Y(n2005) );
  INVX3 U977 ( .A(blockdata[42]), .Y(n2010) );
  INVX3 U978 ( .A(blockdata[43]), .Y(n2015) );
  INVX3 U979 ( .A(blockdata[45]), .Y(n2025) );
  INVX3 U980 ( .A(n1672), .Y(n1956) );
  INVXL U981 ( .A(proc_addr[26]), .Y(n1865) );
  BUFX8 U982 ( .A(n1380), .Y(n1384) );
  CLKBUFX4 U983 ( .A(n1507), .Y(n1506) );
  CLKBUFX4 U984 ( .A(n1522), .Y(n1521) );
  CLKBUFX4 U985 ( .A(n1555), .Y(n1554) );
  CLKBUFX4 U986 ( .A(n1599), .Y(n1598) );
  CLKBUFX4 U987 ( .A(n1585), .Y(n1584) );
  CLKBUFX4 U988 ( .A(n1538), .Y(n1537) );
  CLKBUFX4 U989 ( .A(n1572), .Y(n1571) );
  BUFX20 U990 ( .A(n1361), .Y(n1375) );
  BUFX8 U991 ( .A(n1364), .Y(n1366) );
  CLKBUFX2 U992 ( .A(n1418), .Y(n1422) );
  CLKBUFX2 U993 ( .A(n1364), .Y(n1365) );
  CLKBUFX2 U994 ( .A(n1414), .Y(n1416) );
  CLKBUFX2 U995 ( .A(n1618), .Y(n1448) );
  INVX3 U996 ( .A(n1942), .Y(n1945) );
  NAND2XL U997 ( .A(n1941), .B(n1618), .Y(n1942) );
  INVX3 U998 ( .A(n1939), .Y(n1940) );
  NAND2XL U999 ( .A(n1941), .B(n1619), .Y(n1939) );
  NAND2X4 U1000 ( .A(n11), .B(n1954), .Y(n1959) );
  INVXL U1001 ( .A(proc_addr[5]), .Y(n1925) );
  MX2XL U1002 ( .A(n1926), .B(n1925), .S0(n1480), .Y(n1927) );
  XOR2X4 U1003 ( .A(n1926), .B(proc_addr[5]), .Y(n1649) );
  XOR2X4 U1004 ( .A(n1893), .B(proc_addr[16]), .Y(n1645) );
  XOR2X4 U1005 ( .A(n1902), .B(proc_addr[13]), .Y(n1646) );
  XOR2X4 U1006 ( .A(proc_addr[23]), .B(tag[18]), .Y(n1630) );
  XOR2X4 U1007 ( .A(tag[2]), .B(proc_addr[7]), .Y(n1633) );
  XOR2X4 U1008 ( .A(tag[5]), .B(proc_addr[10]), .Y(n1632) );
  INVX1 U1009 ( .A(blockdata[81]), .Y(n2046) );
  INVX1 U1010 ( .A(blockdata[82]), .Y(n2051) );
  INVX1 U1011 ( .A(blockdata[72]), .Y(n2001) );
  INVX1 U1012 ( .A(blockdata[73]), .Y(n2006) );
  INVX1 U1013 ( .A(blockdata[74]), .Y(n2011) );
  INVX1 U1014 ( .A(blockdata[75]), .Y(n2016) );
  INVX1 U1015 ( .A(blockdata[76]), .Y(n2021) );
  INVX1 U1016 ( .A(blockdata[78]), .Y(n2031) );
  INVX1 U1017 ( .A(blockdata[79]), .Y(n2036) );
  INVX1 U1018 ( .A(blockdata[80]), .Y(n2041) );
  INVXL U1019 ( .A(blockdata[7]), .Y(n1999) );
  INVX1 U1020 ( .A(blockdata[109]), .Y(n2028) );
  INVX1 U1021 ( .A(blockdata[110]), .Y(n2033) );
  INVX1 U1022 ( .A(blockdata[116]), .Y(n2063) );
  INVX1 U1023 ( .A(blockdata[111]), .Y(n2038) );
  INVX1 U1024 ( .A(blockdata[112]), .Y(n2043) );
  INVX1 U1025 ( .A(blockdata[113]), .Y(n2048) );
  INVX1 U1026 ( .A(blockdata[114]), .Y(n2053) );
  INVX1 U1027 ( .A(blockdata[115]), .Y(n2058) );
  INVX1 U1028 ( .A(blockdata[71]), .Y(n1996) );
  INVX1 U1029 ( .A(blockdata[77]), .Y(n2026) );
  INVX1 U1030 ( .A(blockdata[39]), .Y(n1995) );
  INVXL U1031 ( .A(blockdata[8]), .Y(n2004) );
  INVXL U1032 ( .A(proc_addr[0]), .Y(n1957) );
  INVXL U1033 ( .A(blockdata[20]), .Y(n2064) );
  INVXL U1034 ( .A(blockdata[21]), .Y(n2069) );
  INVXL U1035 ( .A(blockdata[22]), .Y(n2074) );
  INVXL U1036 ( .A(blockdata[23]), .Y(n2079) );
  INVXL U1037 ( .A(blockdata[24]), .Y(n2084) );
  INVXL U1038 ( .A(blockdata[13]), .Y(n2029) );
  INVXL U1039 ( .A(blockdata[14]), .Y(n2034) );
  INVXL U1040 ( .A(blockdata[15]), .Y(n2039) );
  INVXL U1041 ( .A(blockdata[16]), .Y(n2044) );
  INVXL U1042 ( .A(blockdata[17]), .Y(n2049) );
  INVXL U1043 ( .A(blockdata[18]), .Y(n2054) );
  INVXL U1044 ( .A(blockdata[19]), .Y(n2059) );
  INVXL U1045 ( .A(blockdata[25]), .Y(n2089) );
  INVXL U1046 ( .A(blockdata[26]), .Y(n2094) );
  INVXL U1047 ( .A(blockdata[27]), .Y(n2099) );
  INVXL U1048 ( .A(blockdata[28]), .Y(n2104) );
  INVXL U1049 ( .A(blockdata[29]), .Y(n2109) );
  INVXL U1050 ( .A(blockdata[30]), .Y(n2114) );
  INVXL U1051 ( .A(blockdata[10]), .Y(n2014) );
  INVXL U1052 ( .A(blockdata[11]), .Y(n2019) );
  INVXL U1053 ( .A(blockdata[12]), .Y(n2024) );
  INVXL U1054 ( .A(blockdata[31]), .Y(n2122) );
  INVXL U1055 ( .A(blockdata[96]), .Y(n1963) );
  INVXL U1056 ( .A(blockdata[97]), .Y(n1968) );
  INVXL U1057 ( .A(blockdata[99]), .Y(n1978) );
  INVXL U1058 ( .A(blockdata[100]), .Y(n1983) );
  INVXL U1059 ( .A(blockdata[101]), .Y(n1988) );
  INVXL U1060 ( .A(blockdata[102]), .Y(n1993) );
  INVXL U1061 ( .A(blockdata[103]), .Y(n1998) );
  INVXL U1062 ( .A(blockdata[104]), .Y(n2003) );
  INVXL U1063 ( .A(blockdata[105]), .Y(n2008) );
  INVXL U1064 ( .A(blockdata[106]), .Y(n2013) );
  INVXL U1065 ( .A(blockdata[107]), .Y(n2018) );
  INVXL U1066 ( .A(blockdata[108]), .Y(n2023) );
  INVXL U1067 ( .A(blockdata[92]), .Y(n2101) );
  INVXL U1068 ( .A(blockdata[65]), .Y(n1966) );
  INVXL U1069 ( .A(blockdata[66]), .Y(n1971) );
  INVXL U1070 ( .A(blockdata[67]), .Y(n1976) );
  INVXL U1071 ( .A(blockdata[68]), .Y(n1981) );
  INVXL U1072 ( .A(blockdata[93]), .Y(n2106) );
  INVXL U1073 ( .A(blockdata[94]), .Y(n2111) );
  INVXL U1074 ( .A(blockdata[95]), .Y(n2117) );
  INVXL U1075 ( .A(blockdata[60]), .Y(n2100) );
  INVXL U1076 ( .A(blockdata[64]), .Y(n1961) );
  INVXL U1077 ( .A(blockdata[57]), .Y(n2085) );
  INVXL U1078 ( .A(blockdata[58]), .Y(n2090) );
  INVXL U1079 ( .A(blockdata[59]), .Y(n2095) );
  INVXL U1080 ( .A(blockdata[61]), .Y(n2105) );
  INVXL U1081 ( .A(blockdata[62]), .Y(n2110) );
  INVXL U1082 ( .A(blockdata[63]), .Y(n2115) );
  INVXL U1083 ( .A(blockdata[32]), .Y(n1960) );
  INVXL U1084 ( .A(blockdata[87]), .Y(n2076) );
  INVXL U1085 ( .A(blockdata[83]), .Y(n2056) );
  INVXL U1086 ( .A(blockdata[84]), .Y(n2061) );
  INVXL U1087 ( .A(blockdata[85]), .Y(n2066) );
  INVXL U1088 ( .A(blockdata[86]), .Y(n2071) );
  INVXL U1089 ( .A(blockdata[88]), .Y(n2081) );
  INVXL U1090 ( .A(blockdata[89]), .Y(n2086) );
  INVXL U1091 ( .A(blockdata[90]), .Y(n2091) );
  INVXL U1092 ( .A(blockdata[91]), .Y(n2096) );
  INVXL U1093 ( .A(blockdata[51]), .Y(n2055) );
  INVXL U1094 ( .A(blockdata[52]), .Y(n2060) );
  INVXL U1095 ( .A(blockdata[53]), .Y(n2065) );
  INVXL U1096 ( .A(blockdata[54]), .Y(n2070) );
  INVXL U1097 ( .A(blockdata[55]), .Y(n2075) );
  INVXL U1098 ( .A(blockdata[56]), .Y(n2080) );
  INVXL U1099 ( .A(blockdata[46]), .Y(n2030) );
  INVXL U1100 ( .A(blockdata[47]), .Y(n2035) );
  INVXL U1101 ( .A(blockdata[48]), .Y(n2040) );
  INVXL U1102 ( .A(blockdata[49]), .Y(n2045) );
  INVXL U1103 ( .A(blockdata[50]), .Y(n2050) );
  INVXL U1104 ( .A(blockdata[69]), .Y(n1986) );
  INVXL U1105 ( .A(blockdata[70]), .Y(n1991) );
  INVXL U1106 ( .A(blockdata[37]), .Y(n1985) );
  INVX1 U1107 ( .A(blockdata[118]), .Y(n2073) );
  INVX1 U1108 ( .A(blockdata[119]), .Y(n2078) );
  INVX1 U1109 ( .A(blockdata[120]), .Y(n2083) );
  INVX1 U1110 ( .A(blockdata[121]), .Y(n2088) );
  INVX1 U1111 ( .A(blockdata[122]), .Y(n2093) );
  INVX1 U1112 ( .A(blockdata[117]), .Y(n2068) );
  INVX1 U1113 ( .A(blockdata[123]), .Y(n2098) );
  INVX1 U1114 ( .A(blockdata[124]), .Y(n2103) );
  INVX1 U1115 ( .A(blockdata[125]), .Y(n2108) );
  INVX1 U1116 ( .A(blockdata[126]), .Y(n2113) );
  INVX1 U1117 ( .A(blockdata[127]), .Y(n2120) );
  INVXL U1118 ( .A(blockdata[9]), .Y(n2009) );
  XOR2X4 U1119 ( .A(n1866), .B(proc_addr[26]), .Y(n1652) );
  MXI2XL U1120 ( .A(n471), .B(n1946), .S0(n1857), .Y(n487) );
  XOR2X4 U1121 ( .A(n1863), .B(proc_addr[27]), .Y(n1655) );
  XOR2X4 U1122 ( .A(n1896), .B(proc_addr[15]), .Y(n1657) );
  MXI4XL U1123 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n1442), .S1(n1407), .Y(n1283) );
  MXI4XL U1124 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n1442), .S1(n1407), .Y(n1282) );
  MXI4XL U1125 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n1442), .S1(n1407), .Y(n1281) );
  MXI4XL U1126 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n1442), .S1(n1407), .Y(n1280) );
  MXI4XL U1127 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n1442), .S1(n1407), .Y(n1285) );
  MXI4XL U1128 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n1442), .S1(n1407), .Y(n1284) );
  MXI2X1 U1129 ( .A(n1214), .B(n1215), .S0(n1367), .Y(blockdata[44]) );
  MXI4XL U1130 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n1437), .S1(n1402), .Y(n1214) );
  MXI4XL U1131 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n1442), .S1(n1389), .Y(n1058) );
  MXI4XL U1132 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n1430), .S1(n1389), .Y(n1066) );
  MXI4XL U1133 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n1433), .S1(n1389), .Y(n1067) );
  MXI4XL U1134 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n1433), .S1(n1389), .Y(n1064) );
  MXI4XL U1135 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n1433), .S1(n1389), .Y(n1065) );
  MXI4XL U1136 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n1439), .S1(n1389), .Y(n1062) );
  MXI4XL U1137 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n1425), .S1(n1389), .Y(n1063) );
  MXI4XL U1138 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n1425), .S1(n1389), .Y(n1060) );
  MXI4XL U1139 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n1442), .S1(n1389), .Y(n1061) );
  MXI4XL U1140 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n1425), .S1(n1389), .Y(n1068) );
  MXI4XL U1141 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n1433), .S1(n1389), .Y(n1069) );
  CLKBUFX3 U1142 ( .A(n1385), .Y(n1404) );
  CLKBUFX3 U1143 ( .A(n1385), .Y(n1403) );
  CLKBUFX3 U1144 ( .A(n1387), .Y(n1397) );
  CLKBUFX3 U1145 ( .A(n1379), .Y(n1401) );
  CLKBUFX3 U1146 ( .A(n1385), .Y(n1395) );
  CLKBUFX3 U1147 ( .A(n1387), .Y(n1400) );
  CLKBUFX3 U1148 ( .A(n1377), .Y(n1394) );
  CLKBUFX3 U1149 ( .A(n1386), .Y(n1399) );
  CLKBUFX3 U1150 ( .A(n1386), .Y(n1398) );
  CLKBUFX3 U1151 ( .A(n1385), .Y(n1405) );
  CLKBUFX3 U1152 ( .A(n1377), .Y(n1406) );
  CLKBUFX3 U1153 ( .A(n1384), .Y(n1408) );
  CLKBUFX3 U1154 ( .A(n1377), .Y(n1407) );
  CLKBUFX3 U1155 ( .A(n1377), .Y(n1391) );
  CLKBUFX3 U1156 ( .A(n1385), .Y(n1393) );
  CLKBUFX3 U1157 ( .A(n1377), .Y(n1392) );
  CLKBUFX3 U1158 ( .A(n1385), .Y(n1390) );
  CLKBUFX3 U1159 ( .A(n1385), .Y(n1402) );
  CLKBUFX3 U1160 ( .A(n1387), .Y(n1396) );
  CLKBUFX3 U1161 ( .A(n1363), .Y(n1371) );
  CLKBUFX3 U1162 ( .A(n1359), .Y(n1369) );
  CLKBUFX3 U1163 ( .A(n1359), .Y(n1368) );
  CLKBUFX3 U1164 ( .A(n1363), .Y(n1372) );
  CLKBUFX3 U1165 ( .A(n1359), .Y(n1367) );
  CLKBUFX3 U1166 ( .A(n1423), .Y(n1438) );
  CLKBUFX3 U1167 ( .A(n1423), .Y(n1436) );
  CLKBUFX3 U1168 ( .A(n1418), .Y(n1431) );
  CLKBUFX3 U1169 ( .A(n1418), .Y(n1435) );
  CLKBUFX3 U1170 ( .A(n1418), .Y(n1434) );
  CLKBUFX3 U1171 ( .A(n1424), .Y(n1429) );
  CLKBUFX3 U1172 ( .A(n1423), .Y(n1439) );
  CLKBUFX3 U1173 ( .A(n1422), .Y(n1441) );
  CLKBUFX3 U1174 ( .A(n1422), .Y(n1440) );
  CLKBUFX3 U1175 ( .A(n1418), .Y(n1442) );
  CLKBUFX3 U1176 ( .A(n1424), .Y(n1428) );
  CLKBUFX3 U1177 ( .A(n1422), .Y(n1427) );
  CLKBUFX3 U1178 ( .A(n1417), .Y(n1432) );
  CLKBUFX3 U1179 ( .A(n1422), .Y(n1426) );
  CLKBUFX3 U1180 ( .A(n1423), .Y(n1437) );
  CLKBUFX3 U1181 ( .A(n1423), .Y(n1425) );
  CLKBUFX3 U1182 ( .A(n1602), .Y(n1608) );
  CLKBUFX3 U1183 ( .A(n1), .Y(n1593) );
  CLKBUFX3 U1184 ( .A(n1586), .Y(n1579) );
  CLKBUFX3 U1185 ( .A(n1559), .Y(n1566) );
  CLKBUFX3 U1186 ( .A(n1557), .Y(n1549) );
  CLKBUFX3 U1187 ( .A(n1541), .Y(n1532) );
  CLKBUFX3 U1188 ( .A(n1616), .Y(n1606) );
  CLKBUFX3 U1189 ( .A(n1599), .Y(n1591) );
  CLKBUFX3 U1190 ( .A(n1585), .Y(n1577) );
  CLKBUFX3 U1191 ( .A(n1560), .Y(n1564) );
  CLKBUFX3 U1192 ( .A(n1543), .Y(n1547) );
  CLKBUFX3 U1193 ( .A(n1526), .Y(n1530) );
  CLKBUFX3 U1194 ( .A(n1602), .Y(n1607) );
  CLKBUFX3 U1195 ( .A(n1), .Y(n1592) );
  CLKBUFX3 U1196 ( .A(n1586), .Y(n1578) );
  CLKBUFX3 U1197 ( .A(n1559), .Y(n1565) );
  CLKBUFX3 U1198 ( .A(n1557), .Y(n1548) );
  CLKBUFX3 U1199 ( .A(n1541), .Y(n1531) );
  CLKBUFX3 U1200 ( .A(n1616), .Y(n1605) );
  CLKBUFX3 U1201 ( .A(n1), .Y(n1590) );
  CLKBUFX3 U1202 ( .A(n2), .Y(n1576) );
  CLKBUFX3 U1203 ( .A(n1560), .Y(n1563) );
  CLKBUFX3 U1204 ( .A(n1543), .Y(n1546) );
  CLKBUFX3 U1205 ( .A(n1526), .Y(n1529) );
  CLKBUFX3 U1206 ( .A(n1602), .Y(n1611) );
  CLKBUFX3 U1207 ( .A(n1), .Y(n1596) );
  CLKBUFX3 U1208 ( .A(n2), .Y(n1582) );
  CLKBUFX3 U1209 ( .A(n1559), .Y(n1569) );
  CLKBUFX3 U1210 ( .A(n1542), .Y(n1552) );
  CLKBUFX3 U1211 ( .A(n1539), .Y(n1535) );
  CLKBUFX3 U1212 ( .A(n1602), .Y(n1612) );
  CLKBUFX3 U1213 ( .A(n1599), .Y(n1597) );
  CLKBUFX3 U1214 ( .A(n2), .Y(n1583) );
  CLKBUFX3 U1215 ( .A(n1559), .Y(n1570) );
  CLKBUFX3 U1216 ( .A(n1542), .Y(n1553) );
  CLKBUFX3 U1217 ( .A(n1539), .Y(n1536) );
  CLKBUFX3 U1218 ( .A(n1615), .Y(n1609) );
  CLKBUFX3 U1219 ( .A(n1615), .Y(n1610) );
  CLKBUFX3 U1220 ( .A(n1600), .Y(n1594) );
  CLKBUFX3 U1221 ( .A(n1600), .Y(n1595) );
  CLKBUFX3 U1222 ( .A(n2), .Y(n1580) );
  CLKBUFX3 U1223 ( .A(n1586), .Y(n1581) );
  CLKBUFX3 U1224 ( .A(n1573), .Y(n1567) );
  CLKBUFX3 U1225 ( .A(n1573), .Y(n1568) );
  CLKBUFX3 U1226 ( .A(n1556), .Y(n1550) );
  CLKBUFX3 U1227 ( .A(n1556), .Y(n1551) );
  CLKBUFX3 U1228 ( .A(n1540), .Y(n1533) );
  CLKBUFX3 U1229 ( .A(n1540), .Y(n1534) );
  CLKBUFX3 U1230 ( .A(n1523), .Y(n1514) );
  CLKBUFX3 U1231 ( .A(n5), .Y(n1515) );
  CLKBUFX3 U1232 ( .A(n1523), .Y(n1513) );
  CLKBUFX3 U1233 ( .A(n2124), .Y(n1499) );
  CLKBUFX3 U1234 ( .A(n1509), .Y(n1500) );
  CLKBUFX3 U1235 ( .A(n1507), .Y(n1498) );
  CLKBUFX3 U1236 ( .A(n1510), .Y(n1516) );
  CLKBUFX3 U1237 ( .A(n1510), .Y(n1519) );
  CLKBUFX3 U1238 ( .A(n1510), .Y(n1520) );
  CLKBUFX3 U1239 ( .A(n1522), .Y(n1517) );
  CLKBUFX3 U1240 ( .A(n1510), .Y(n1518) );
  CLKBUFX3 U1241 ( .A(n1509), .Y(n1501) );
  CLKBUFX3 U1242 ( .A(n2124), .Y(n1504) );
  CLKBUFX3 U1243 ( .A(n1507), .Y(n1505) );
  CLKBUFX3 U1244 ( .A(n1508), .Y(n1502) );
  CLKBUFX3 U1245 ( .A(n1508), .Y(n1503) );
  CLKBUFX3 U1246 ( .A(n1617), .Y(n1604) );
  CLKBUFX3 U1247 ( .A(n1601), .Y(n1589) );
  CLKBUFX3 U1248 ( .A(n1587), .Y(n1575) );
  CLKBUFX3 U1249 ( .A(n1573), .Y(n1562) );
  CLKBUFX3 U1250 ( .A(n1558), .Y(n1545) );
  CLKBUFX3 U1251 ( .A(n1538), .Y(n1528) );
  CLKBUFX3 U1252 ( .A(n1522), .Y(n1512) );
  CLKBUFX3 U1253 ( .A(n1507), .Y(n1497) );
  CLKBUFX3 U1254 ( .A(n1617), .Y(n1603) );
  CLKBUFX3 U1255 ( .A(n1601), .Y(n1588) );
  CLKBUFX3 U1256 ( .A(n1587), .Y(n1574) );
  CLKBUFX3 U1257 ( .A(n1560), .Y(n1561) );
  CLKBUFX3 U1258 ( .A(n1558), .Y(n1544) );
  CLKBUFX3 U1259 ( .A(n1538), .Y(n1527) );
  CLKBUFX3 U1260 ( .A(n1510), .Y(n1511) );
  CLKBUFX3 U1261 ( .A(n2124), .Y(n1496) );
  CLKBUFX3 U1262 ( .A(n1377), .Y(n1388) );
  CLKBUFX3 U1263 ( .A(n6), .Y(n1557) );
  CLKBUFX3 U1264 ( .A(n1525), .Y(n1541) );
  CLKBUFX3 U1265 ( .A(n1524), .Y(n1539) );
  CLKBUFX3 U1266 ( .A(n1), .Y(n1600) );
  CLKBUFX3 U1267 ( .A(n3), .Y(n1573) );
  CLKBUFX3 U1268 ( .A(n6), .Y(n1556) );
  CLKBUFX3 U1269 ( .A(n1525), .Y(n1540) );
  CLKBUFX3 U1270 ( .A(n2), .Y(n1585) );
  CLKBUFX3 U1271 ( .A(n1559), .Y(n1572) );
  CLKBUFX3 U1272 ( .A(n1542), .Y(n1555) );
  CLKBUFX3 U1273 ( .A(n1524), .Y(n1538) );
  CLKBUFX3 U1274 ( .A(n2124), .Y(n1509) );
  CLKBUFX3 U1275 ( .A(n2124), .Y(n1508) );
  CLKBUFX3 U1276 ( .A(n3), .Y(n1560) );
  CLKBUFX3 U1277 ( .A(n6), .Y(n1543) );
  CLKBUFX3 U1278 ( .A(n7), .Y(n1525) );
  CLKBUFX3 U1279 ( .A(n4), .Y(n1602) );
  CLKBUFX3 U1280 ( .A(n3), .Y(n1559) );
  CLKBUFX3 U1281 ( .A(n6), .Y(n1542) );
  CLKBUFX3 U1282 ( .A(n7), .Y(n1524) );
  CLKBUFX3 U1283 ( .A(n1376), .Y(n1360) );
  CLKBUFX3 U1284 ( .A(n1376), .Y(n1359) );
  CLKBUFX3 U1285 ( .A(n1358), .Y(n1364) );
  CLKBUFX3 U1286 ( .A(n1376), .Y(n1358) );
  CLKINVX1 U1287 ( .A(n1938), .Y(n1941) );
  CLKBUFX3 U1288 ( .A(n1492), .Y(n1495) );
  CLKINVX1 U1289 ( .A(n1681), .Y(n1857) );
  NAND3BXL U1290 ( .AN(N32), .B(n1619), .C(n1621), .Y(n1681) );
  CLKINVX1 U1291 ( .A(n1928), .Y(n1929) );
  NAND3BXL U1292 ( .AN(N32), .B(n1618), .C(n1621), .Y(n1928) );
  CLKINVX1 U1293 ( .A(n1930), .Y(n1931) );
  NAND3BXL U1294 ( .AN(n1618), .B(N32), .C(n1621), .Y(n1930) );
  CLKINVX1 U1295 ( .A(n1932), .Y(n1933) );
  NAND3BXL U1296 ( .AN(n13), .B(n1618), .C(n1621), .Y(n1932) );
  CLKINVX1 U1297 ( .A(n1934), .Y(n1935) );
  NAND3BXL U1298 ( .AN(n1618), .B(N33), .C(n13), .Y(n1934) );
  CLKINVX1 U1299 ( .A(n1936), .Y(n1937) );
  NAND3BXL U1300 ( .AN(n1621), .B(n1618), .C(n13), .Y(n1936) );
  CLKINVX1 U1301 ( .A(n1959), .Y(n1955) );
  MX2XL U1302 ( .A(n1922), .B(n1921), .S0(n1476), .Y(n1923) );
  INVXL U1303 ( .A(proc_addr[6]), .Y(n1921) );
  MX2XL U1304 ( .A(n63), .B(n1919), .S0(n1484), .Y(n1920) );
  INVXL U1305 ( .A(proc_addr[7]), .Y(n1919) );
  MX2XL U1306 ( .A(n1917), .B(n1916), .S0(n1486), .Y(n1918) );
  INVXL U1307 ( .A(proc_addr[8]), .Y(n1916) );
  INVXL U1308 ( .A(tag[3]), .Y(n1917) );
  MX2XL U1309 ( .A(n1914), .B(n1913), .S0(n1483), .Y(n1915) );
  INVXL U1310 ( .A(proc_addr[9]), .Y(n1913) );
  MX2XL U1311 ( .A(n1911), .B(n1910), .S0(n1482), .Y(n1912) );
  INVXL U1312 ( .A(proc_addr[10]), .Y(n1910) );
  INVXL U1313 ( .A(tag[5]), .Y(n1911) );
  MX2XL U1314 ( .A(n1908), .B(n1907), .S0(n1488), .Y(n1909) );
  INVXL U1315 ( .A(proc_addr[11]), .Y(n1907) );
  MX2XL U1316 ( .A(n1905), .B(n1904), .S0(n1483), .Y(n1906) );
  INVXL U1317 ( .A(proc_addr[12]), .Y(n1904) );
  MX2XL U1318 ( .A(n1902), .B(n1901), .S0(n1473), .Y(n1903) );
  INVXL U1319 ( .A(proc_addr[13]), .Y(n1901) );
  MX2XL U1320 ( .A(n1896), .B(n1895), .S0(n1489), .Y(n1897) );
  CLKINVX1 U1321 ( .A(proc_addr[15]), .Y(n1895) );
  MX2XL U1322 ( .A(n1893), .B(n1892), .S0(n1474), .Y(n1894) );
  INVXL U1323 ( .A(proc_addr[16]), .Y(n1892) );
  MX2XL U1324 ( .A(n1890), .B(n1889), .S0(n1485), .Y(n1891) );
  INVXL U1325 ( .A(proc_addr[17]), .Y(n1889) );
  MX2XL U1326 ( .A(n1887), .B(n1886), .S0(n1484), .Y(n1888) );
  INVXL U1327 ( .A(proc_addr[18]), .Y(n1886) );
  MX2XL U1328 ( .A(n1884), .B(n88), .S0(n1489), .Y(n1885) );
  MX2XL U1329 ( .A(n9), .B(n1882), .S0(n1487), .Y(n1883) );
  INVXL U1330 ( .A(proc_addr[20]), .Y(n1882) );
  MX2XL U1331 ( .A(n1880), .B(n1879), .S0(n1487), .Y(n1881) );
  CLKINVX1 U1332 ( .A(proc_addr[21]), .Y(n1879) );
  MX2XL U1333 ( .A(n57), .B(n1874), .S0(n1486), .Y(n1875) );
  INVXL U1334 ( .A(proc_addr[23]), .Y(n1874) );
  MX2XL U1335 ( .A(n1872), .B(n1871), .S0(n1490), .Y(n1873) );
  INVXL U1336 ( .A(proc_addr[24]), .Y(n1871) );
  MX2XL U1337 ( .A(n1869), .B(n1868), .S0(n1483), .Y(n1870) );
  INVXL U1338 ( .A(proc_addr[25]), .Y(n1868) );
  MX2XL U1339 ( .A(n1863), .B(n1862), .S0(n1488), .Y(n1864) );
  INVXL U1340 ( .A(proc_addr[27]), .Y(n1862) );
  INVXL U1341 ( .A(proc_addr[28]), .Y(n1859) );
  MX2XL U1342 ( .A(n32), .B(n40), .S0(n1484), .Y(n1858) );
  NAND2XL U1343 ( .A(n8), .B(proc_stall), .Y(n1679) );
  CLKINVX1 U1344 ( .A(blockdata[44]), .Y(n2020) );
  NAND2X1 U1345 ( .A(mem_rdata[42]), .B(n1483), .Y(n1774) );
  NAND2X1 U1346 ( .A(mem_rdata[43]), .B(n1484), .Y(n1773) );
  NAND2X1 U1347 ( .A(mem_rdata[44]), .B(n1475), .Y(n1772) );
  NAND2X1 U1348 ( .A(mem_rdata[45]), .B(n1489), .Y(n1771) );
  NAND2X1 U1349 ( .A(mem_rdata[46]), .B(n1481), .Y(n1770) );
  NAND2X1 U1350 ( .A(mem_rdata[47]), .B(n1479), .Y(n1769) );
  NAND2X1 U1351 ( .A(mem_rdata[48]), .B(n1479), .Y(n1768) );
  NAND2X1 U1352 ( .A(mem_rdata[49]), .B(n1488), .Y(n1767) );
  NAND2X1 U1353 ( .A(mem_rdata[50]), .B(n1474), .Y(n1766) );
  NAND2X1 U1354 ( .A(mem_rdata[51]), .B(n1487), .Y(n1765) );
  NAND2X1 U1355 ( .A(mem_rdata[52]), .B(n1473), .Y(n1764) );
  NAND2X1 U1356 ( .A(mem_rdata[55]), .B(n1480), .Y(n1761) );
  NAND2X1 U1357 ( .A(mem_rdata[56]), .B(n1481), .Y(n1760) );
  NAND2X1 U1358 ( .A(mem_rdata[57]), .B(n1490), .Y(n1759) );
  NAND2X1 U1359 ( .A(mem_rdata[58]), .B(n1480), .Y(n1758) );
  NAND2X1 U1360 ( .A(mem_rdata[59]), .B(n1484), .Y(n1757) );
  NAND2X1 U1361 ( .A(mem_rdata[60]), .B(n1490), .Y(n1756) );
  NAND2X1 U1362 ( .A(mem_rdata[61]), .B(n1488), .Y(n1755) );
  NAND2X1 U1363 ( .A(mem_rdata[62]), .B(n1473), .Y(n1754) );
  NAND2X1 U1364 ( .A(mem_rdata[32]), .B(n1484), .Y(n1784) );
  NAND2X1 U1365 ( .A(mem_rdata[33]), .B(n1476), .Y(n1783) );
  NAND2X1 U1366 ( .A(mem_rdata[34]), .B(n1483), .Y(n1782) );
  NAND2X1 U1367 ( .A(mem_rdata[35]), .B(n1490), .Y(n1781) );
  NAND2X1 U1368 ( .A(mem_rdata[36]), .B(n1487), .Y(n1780) );
  NAND2X1 U1369 ( .A(mem_rdata[37]), .B(n1477), .Y(n1779) );
  NAND2X1 U1370 ( .A(mem_rdata[39]), .B(n1479), .Y(n1777) );
  NAND2X1 U1371 ( .A(mem_rdata[106]), .B(n1481), .Y(n1702) );
  NAND2X1 U1372 ( .A(mem_rdata[107]), .B(n1482), .Y(n1701) );
  NAND2X1 U1373 ( .A(mem_rdata[108]), .B(n1479), .Y(n1700) );
  NAND2X1 U1374 ( .A(mem_rdata[109]), .B(n1479), .Y(n1699) );
  NAND2X1 U1375 ( .A(mem_rdata[110]), .B(n1486), .Y(n1698) );
  NAND2X1 U1376 ( .A(mem_rdata[111]), .B(n1487), .Y(n1697) );
  NAND2X1 U1377 ( .A(mem_rdata[113]), .B(n1482), .Y(n1695) );
  NAND2X1 U1378 ( .A(mem_rdata[114]), .B(n1476), .Y(n1694) );
  NAND2X1 U1379 ( .A(mem_rdata[115]), .B(n1478), .Y(n1693) );
  NAND2X1 U1380 ( .A(mem_rdata[116]), .B(n1481), .Y(n1692) );
  NAND2X1 U1381 ( .A(mem_rdata[117]), .B(n1481), .Y(n1691) );
  NAND2X1 U1382 ( .A(mem_rdata[118]), .B(n1474), .Y(n1690) );
  NAND2X1 U1383 ( .A(mem_rdata[74]), .B(n1489), .Y(n1739) );
  NAND2X1 U1384 ( .A(mem_rdata[76]), .B(n1485), .Y(n1737) );
  NAND2X1 U1385 ( .A(mem_rdata[77]), .B(n1486), .Y(n1736) );
  NAND2X1 U1386 ( .A(mem_rdata[78]), .B(n1479), .Y(n1735) );
  NAND2X1 U1387 ( .A(mem_rdata[79]), .B(n1489), .Y(n1734) );
  NAND2X1 U1388 ( .A(mem_rdata[80]), .B(n1473), .Y(n1733) );
  NAND2X1 U1389 ( .A(mem_rdata[81]), .B(n1476), .Y(n1732) );
  NAND2X1 U1390 ( .A(mem_rdata[82]), .B(n1483), .Y(n1731) );
  NAND2X1 U1391 ( .A(mem_rdata[83]), .B(n1479), .Y(n1730) );
  NAND2X1 U1392 ( .A(mem_rdata[84]), .B(n1481), .Y(n1729) );
  NAND2X1 U1393 ( .A(mem_rdata[85]), .B(n1474), .Y(n1728) );
  NAND2X1 U1394 ( .A(mem_rdata[86]), .B(n1486), .Y(n1727) );
  NAND2X1 U1395 ( .A(mem_rdata[87]), .B(n1481), .Y(n1726) );
  NAND2X1 U1396 ( .A(mem_rdata[88]), .B(n1474), .Y(n1725) );
  NAND2X1 U1397 ( .A(mem_rdata[89]), .B(n1481), .Y(n1724) );
  NAND2X1 U1398 ( .A(mem_rdata[90]), .B(n1486), .Y(n1723) );
  NAND2X1 U1399 ( .A(mem_rdata[91]), .B(n1479), .Y(n1722) );
  NAND2X1 U1400 ( .A(mem_rdata[92]), .B(n1480), .Y(n1721) );
  NAND2X1 U1401 ( .A(mem_rdata[93]), .B(n1484), .Y(n1720) );
  NAND2X1 U1402 ( .A(mem_rdata[94]), .B(n1479), .Y(n1719) );
  NAND2X1 U1403 ( .A(mem_rdata[95]), .B(n1481), .Y(n1718) );
  NAND2X1 U1404 ( .A(mem_rdata[96]), .B(n1477), .Y(n1712) );
  NAND2X1 U1405 ( .A(mem_rdata[98]), .B(n1481), .Y(n1710) );
  NAND2X1 U1406 ( .A(mem_rdata[99]), .B(n1481), .Y(n1709) );
  NAND2X1 U1407 ( .A(mem_rdata[100]), .B(n1480), .Y(n1708) );
  NAND2X1 U1408 ( .A(mem_rdata[67]), .B(n1482), .Y(n1746) );
  NAND2X1 U1409 ( .A(mem_rdata[68]), .B(n1484), .Y(n1745) );
  NAND2X1 U1410 ( .A(mem_rdata[71]), .B(n1478), .Y(n1742) );
  NAND2X1 U1411 ( .A(mem_rdata[40]), .B(n1473), .Y(n1776) );
  NAND2X1 U1412 ( .A(mem_rdata[41]), .B(n1484), .Y(n1775) );
  NAND2X1 U1413 ( .A(mem_rdata[104]), .B(n1483), .Y(n1704) );
  NAND2X1 U1414 ( .A(mem_rdata[105]), .B(n1479), .Y(n1703) );
  NAND2X1 U1415 ( .A(mem_rdata[72]), .B(n1479), .Y(n1741) );
  NAND2X1 U1416 ( .A(mem_rdata[73]), .B(n1479), .Y(n1740) );
  NAND2X1 U1417 ( .A(mem_rdata[20]), .B(n1477), .Y(n1808) );
  NAND2X1 U1418 ( .A(mem_rdata[21]), .B(n1475), .Y(n1806) );
  NAND2X1 U1419 ( .A(mem_rdata[22]), .B(n1486), .Y(n1804) );
  NAND2X1 U1420 ( .A(mem_rdata[23]), .B(n1484), .Y(n1802) );
  NAND2X1 U1421 ( .A(mem_rdata[24]), .B(n1476), .Y(n1800) );
  NAND2X1 U1422 ( .A(mem_rdata[25]), .B(n1483), .Y(n1798) );
  NAND2X1 U1423 ( .A(mem_rdata[26]), .B(n1483), .Y(n1796) );
  NAND2X1 U1424 ( .A(mem_rdata[27]), .B(n1478), .Y(n1794) );
  NAND2X1 U1425 ( .A(mem_rdata[28]), .B(n1478), .Y(n1792) );
  NAND2X1 U1426 ( .A(mem_rdata[29]), .B(n1485), .Y(n1790) );
  NAND2X1 U1427 ( .A(mem_rdata[30]), .B(n1481), .Y(n1788) );
  NAND2X1 U1428 ( .A(mem_rdata[31]), .B(n1475), .Y(n1786) );
  NAND2X1 U1429 ( .A(mem_rdata[10]), .B(n1482), .Y(n1828) );
  NAND2X1 U1430 ( .A(mem_rdata[11]), .B(n1490), .Y(n1826) );
  NAND2X1 U1431 ( .A(mem_rdata[12]), .B(n1485), .Y(n1824) );
  NAND2X1 U1432 ( .A(mem_rdata[14]), .B(n1476), .Y(n1820) );
  NAND2X1 U1433 ( .A(mem_rdata[16]), .B(n1475), .Y(n1816) );
  NAND2X1 U1434 ( .A(mem_rdata[17]), .B(n1489), .Y(n1814) );
  NAND2X1 U1435 ( .A(mem_rdata[18]), .B(n1480), .Y(n1812) );
  NAND2X1 U1436 ( .A(mem_rdata[19]), .B(n1487), .Y(n1810) );
  NAND2X1 U1437 ( .A(mem_rdata[0]), .B(n1488), .Y(n1848) );
  NAND2X1 U1438 ( .A(mem_rdata[1]), .B(n1482), .Y(n1846) );
  NAND2X1 U1439 ( .A(mem_rdata[2]), .B(n1479), .Y(n1844) );
  NAND2X1 U1440 ( .A(mem_rdata[3]), .B(n1473), .Y(n1842) );
  NAND2X1 U1441 ( .A(mem_rdata[4]), .B(n1477), .Y(n1840) );
  NAND2X1 U1442 ( .A(mem_rdata[5]), .B(n1483), .Y(n1838) );
  NAND2X1 U1443 ( .A(mem_rdata[6]), .B(n1488), .Y(n1836) );
  NAND2X1 U1444 ( .A(mem_rdata[7]), .B(n1478), .Y(n1834) );
  OA22XL U1445 ( .A0(n29), .A1(n1961), .B0(n17), .B1(n1960), .Y(n1962) );
  OA22XL U1446 ( .A0(n29), .A1(n1966), .B0(n17), .B1(n1965), .Y(n1967) );
  OA22XL U1447 ( .A0(n29), .A1(n1971), .B0(n17), .B1(n1970), .Y(n1972) );
  OA22XL U1448 ( .A0(n29), .A1(n1976), .B0(n17), .B1(n1975), .Y(n1977) );
  OA22XL U1449 ( .A0(n29), .A1(n1981), .B0(n17), .B1(n1980), .Y(n1982) );
  OA22XL U1450 ( .A0(n29), .A1(n1986), .B0(n17), .B1(n1985), .Y(n1987) );
  OA22XL U1451 ( .A0(n29), .A1(n1991), .B0(n17), .B1(n1990), .Y(n1992) );
  OA22XL U1452 ( .A0(n29), .A1(n2011), .B0(n17), .B1(n2010), .Y(n2012) );
  OA22XL U1453 ( .A0(n29), .A1(n2016), .B0(n17), .B1(n2015), .Y(n2017) );
  OA22XL U1454 ( .A0(n29), .A1(n2021), .B0(n17), .B1(n2020), .Y(n2022) );
  OA22XL U1455 ( .A0(n29), .A1(n2026), .B0(n17), .B1(n2025), .Y(n2027) );
  OA22XL U1456 ( .A0(n29), .A1(n2031), .B0(n17), .B1(n2030), .Y(n2032) );
  OA22XL U1457 ( .A0(n29), .A1(n2036), .B0(n17), .B1(n2035), .Y(n2037) );
  OA22XL U1458 ( .A0(n29), .A1(n2041), .B0(n17), .B1(n2040), .Y(n2042) );
  OA22XL U1459 ( .A0(n29), .A1(n2046), .B0(n17), .B1(n2045), .Y(n2047) );
  OA22XL U1460 ( .A0(n29), .A1(n2051), .B0(n17), .B1(n2050), .Y(n2052) );
  OA22XL U1461 ( .A0(n29), .A1(n2056), .B0(n17), .B1(n2055), .Y(n2057) );
  OA22XL U1462 ( .A0(n29), .A1(n2061), .B0(n17), .B1(n2060), .Y(n2062) );
  OA22XL U1463 ( .A0(n29), .A1(n2066), .B0(n17), .B1(n2065), .Y(n2067) );
  OA22XL U1464 ( .A0(n29), .A1(n2071), .B0(n17), .B1(n2070), .Y(n2072) );
  OA22XL U1465 ( .A0(n29), .A1(n2076), .B0(n17), .B1(n2075), .Y(n2077) );
  OA22XL U1466 ( .A0(n29), .A1(n2081), .B0(n17), .B1(n2080), .Y(n2082) );
  OAI221XL U1467 ( .A0(n31), .A1(n2089), .B0(n1495), .B1(n2088), .C0(n2087), 
        .Y(proc_rdata[25]) );
  OA22XL U1468 ( .A0(n29), .A1(n2086), .B0(n17), .B1(n2085), .Y(n2087) );
  OAI221XL U1469 ( .A0(n31), .A1(n2094), .B0(n1495), .B1(n2093), .C0(n2092), 
        .Y(proc_rdata[26]) );
  OA22XL U1470 ( .A0(n29), .A1(n2091), .B0(n17), .B1(n2090), .Y(n2092) );
  OA22XL U1471 ( .A0(n29), .A1(n2096), .B0(n17), .B1(n2095), .Y(n2097) );
  OAI221XL U1472 ( .A0(n31), .A1(n2104), .B0(n1495), .B1(n2103), .C0(n2102), 
        .Y(proc_rdata[28]) );
  OA22X1 U1473 ( .A0(n29), .A1(n2101), .B0(n17), .B1(n2100), .Y(n2102) );
  OAI221XL U1474 ( .A0(n31), .A1(n2109), .B0(n1495), .B1(n2108), .C0(n2107), 
        .Y(proc_rdata[29]) );
  OA22XL U1475 ( .A0(n29), .A1(n2106), .B0(n17), .B1(n2105), .Y(n2107) );
  OAI221XL U1476 ( .A0(n31), .A1(n2114), .B0(n1495), .B1(n2113), .C0(n2112), 
        .Y(proc_rdata[30]) );
  OA22XL U1477 ( .A0(n29), .A1(n2111), .B0(n17), .B1(n2110), .Y(n2112) );
  OAI221XL U1478 ( .A0(n31), .A1(n2122), .B0(n1495), .B1(n2120), .C0(n2119), 
        .Y(proc_rdata[31]) );
  OA22XL U1479 ( .A0(n29), .A1(n2117), .B0(n17), .B1(n2115), .Y(n2119) );
  NAND2XL U1480 ( .A(mem_rdata[8]), .B(n1490), .Y(n1832) );
  NAND2XL U1481 ( .A(mem_rdata[9]), .B(n1485), .Y(n1830) );
  OA22XL U1482 ( .A0(n29), .A1(n2001), .B0(n17), .B1(n2000), .Y(n2002) );
  OA22XL U1483 ( .A0(n29), .A1(n2006), .B0(n17), .B1(n2005), .Y(n2007) );
  MX2XL U1484 ( .A(n1866), .B(n1865), .S0(n1475), .Y(n1867) );
  MX2XL U1485 ( .A(n1877), .B(n1876), .S0(n1478), .Y(n1878) );
  INVXL U1486 ( .A(proc_addr[22]), .Y(n1876) );
  MXI2XL U1487 ( .A(n472), .B(n1946), .S0(n1929), .Y(n488) );
  MXI2XL U1488 ( .A(n473), .B(n1946), .S0(n1931), .Y(n489) );
  MXI2XL U1489 ( .A(n474), .B(n1946), .S0(n1933), .Y(n490) );
  MXI2XL U1490 ( .A(n475), .B(n1946), .S0(n1935), .Y(n491) );
  MXI2XL U1491 ( .A(n476), .B(n1946), .S0(n1937), .Y(n492) );
  MXI2XL U1492 ( .A(n477), .B(n1946), .S0(n1940), .Y(n493) );
  MXI2XL U1493 ( .A(n478), .B(n1946), .S0(n1945), .Y(n494) );
  MXI4XL U1494 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n1444), .S1(n1409), .Y(n1307) );
  MXI4XL U1495 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n1444), .S1(n1409), .Y(n1306) );
  INVX1 U1496 ( .A(proc_wdata[22]), .Y(n1805) );
  INVX1 U1497 ( .A(proc_wdata[23]), .Y(n1803) );
  INVX1 U1498 ( .A(proc_wdata[20]), .Y(n1809) );
  INVX1 U1499 ( .A(proc_wdata[21]), .Y(n1807) );
  INVX1 U1500 ( .A(proc_wdata[13]), .Y(n1823) );
  INVX1 U1501 ( .A(proc_wdata[14]), .Y(n1821) );
  INVX1 U1502 ( .A(proc_wdata[15]), .Y(n1819) );
  INVX1 U1503 ( .A(proc_wdata[16]), .Y(n1817) );
  INVX1 U1504 ( .A(proc_wdata[17]), .Y(n1815) );
  INVX1 U1505 ( .A(proc_wdata[18]), .Y(n1813) );
  INVX1 U1506 ( .A(proc_wdata[19]), .Y(n1811) );
  INVX1 U1507 ( .A(proc_wdata[10]), .Y(n1829) );
  INVX1 U1508 ( .A(proc_wdata[11]), .Y(n1827) );
  INVX1 U1509 ( .A(proc_wdata[12]), .Y(n1825) );
  INVX1 U1510 ( .A(proc_wdata[0]), .Y(n1850) );
  INVX1 U1511 ( .A(proc_wdata[24]), .Y(n1801) );
  INVX1 U1512 ( .A(proc_wdata[7]), .Y(n1835) );
  INVX1 U1513 ( .A(proc_wdata[1]), .Y(n1847) );
  INVX1 U1514 ( .A(proc_wdata[2]), .Y(n1845) );
  INVX1 U1515 ( .A(proc_wdata[3]), .Y(n1843) );
  INVX1 U1516 ( .A(proc_wdata[4]), .Y(n1841) );
  INVX1 U1517 ( .A(proc_wdata[6]), .Y(n1837) );
  INVX1 U1518 ( .A(proc_wdata[5]), .Y(n1839) );
  INVX1 U1519 ( .A(proc_wdata[27]), .Y(n1795) );
  INVX1 U1520 ( .A(proc_wdata[28]), .Y(n1793) );
  INVX1 U1521 ( .A(proc_wdata[29]), .Y(n1791) );
  INVX1 U1522 ( .A(proc_wdata[30]), .Y(n1789) );
  INVX1 U1523 ( .A(proc_wdata[31]), .Y(n1787) );
  INVX1 U1524 ( .A(proc_wdata[26]), .Y(n1797) );
  INVX1 U1525 ( .A(proc_wdata[25]), .Y(n1799) );
  INVX1 U1526 ( .A(proc_wdata[8]), .Y(n1833) );
  INVX1 U1527 ( .A(proc_wdata[9]), .Y(n1831) );
  MXI2X1 U1528 ( .A(n479), .B(n1944), .S0(n1857), .Y(n495) );
  MXI2X1 U1529 ( .A(n480), .B(n1944), .S0(n1929), .Y(n496) );
  MXI2X1 U1530 ( .A(n481), .B(n1944), .S0(n1931), .Y(n497) );
  MXI2X1 U1531 ( .A(n482), .B(n1944), .S0(n1933), .Y(n498) );
  MXI2X1 U1532 ( .A(n483), .B(n1944), .S0(n1935), .Y(n499) );
  MXI2X1 U1533 ( .A(n484), .B(n1944), .S0(n1937), .Y(n500) );
  MXI2X1 U1534 ( .A(n485), .B(n1944), .S0(n1940), .Y(n501) );
  MXI2X1 U1535 ( .A(n486), .B(n1944), .S0(n1945), .Y(n503) );
  MXI2X1 U1536 ( .A(n1262), .B(n1263), .S0(n1372), .Y(blockdata[20]) );
  MXI4X1 U1537 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n1440), .S1(n1406), .Y(n1263) );
  MXI4X1 U1538 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n1440), .S1(n1406), .Y(n1262) );
  MXI2X1 U1539 ( .A(n1260), .B(n1261), .S0(n1371), .Y(blockdata[21]) );
  MXI4X1 U1540 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n1440), .S1(n1405), .Y(n1261) );
  MXI4X1 U1541 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n1440), .S1(n1405), .Y(n1260) );
  MXI2X1 U1542 ( .A(n1258), .B(n1259), .S0(n1371), .Y(blockdata[22]) );
  MXI4X1 U1543 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n1440), .S1(n1405), .Y(n1259) );
  MXI4X1 U1544 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n1440), .S1(n1405), .Y(n1258) );
  MXI2X1 U1545 ( .A(n1256), .B(n1257), .S0(n1371), .Y(blockdata[23]) );
  MXI4X1 U1546 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n1440), .S1(n1405), .Y(n1257) );
  MXI4X1 U1547 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n1440), .S1(n1405), .Y(n1256) );
  MXI2X1 U1548 ( .A(n1254), .B(n1255), .S0(n1371), .Y(blockdata[24]) );
  MXI4X1 U1549 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n1440), .S1(n1405), .Y(n1255) );
  MXI4X1 U1550 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n1440), .S1(n1405), .Y(n1254) );
  MXI2X1 U1551 ( .A(n1276), .B(n1277), .S0(n1372), .Y(blockdata[13]) );
  MXI4X1 U1552 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n1441), .S1(n1407), .Y(n1277) );
  MXI4X1 U1553 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n1441), .S1(n1407), .Y(n1276) );
  MXI2X1 U1554 ( .A(n1274), .B(n1275), .S0(n1372), .Y(blockdata[14]) );
  MXI4X1 U1555 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n1441), .S1(n1407), .Y(n1275) );
  MXI4X1 U1556 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n1441), .S1(n1407), .Y(n1274) );
  MXI2X1 U1557 ( .A(n1272), .B(n1273), .S0(n1372), .Y(blockdata[15]) );
  MXI4X1 U1558 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n1441), .S1(n1406), .Y(n1273) );
  MXI4X1 U1559 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n1441), .S1(n1406), .Y(n1272) );
  MXI2X1 U1560 ( .A(n1270), .B(n1271), .S0(n1372), .Y(blockdata[16]) );
  MXI4X1 U1561 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n1441), .S1(n1406), .Y(n1271) );
  MXI4X1 U1562 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n1441), .S1(n1406), .Y(n1270) );
  MXI2X1 U1563 ( .A(n1268), .B(n1269), .S0(n1372), .Y(blockdata[17]) );
  MXI4X1 U1564 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n1441), .S1(n1406), .Y(n1269) );
  MXI4X1 U1565 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n1441), .S1(n1406), .Y(n1268) );
  MXI2X1 U1566 ( .A(n1266), .B(n1267), .S0(n1372), .Y(blockdata[18]) );
  MXI4X1 U1567 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n1440), .S1(n1406), .Y(n1267) );
  MXI4X1 U1568 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n1441), .S1(n1406), .Y(n1266) );
  MXI2X1 U1569 ( .A(n1264), .B(n1265), .S0(n1372), .Y(blockdata[19]) );
  MXI4X1 U1570 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n1440), .S1(n1406), .Y(n1265) );
  MXI4X1 U1571 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n1440), .S1(n1406), .Y(n1264) );
  MXI2X1 U1572 ( .A(n1252), .B(n1253), .S0(n1371), .Y(blockdata[25]) );
  MXI4X1 U1573 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n1439), .S1(n1405), .Y(n1253) );
  MXI4X1 U1574 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n1439), .S1(n1405), .Y(n1252) );
  MXI2X1 U1575 ( .A(n1250), .B(n1251), .S0(n1371), .Y(blockdata[26]) );
  MXI4X1 U1576 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n1439), .S1(n1405), .Y(n1251) );
  MXI4X1 U1577 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n1439), .S1(n1405), .Y(n1250) );
  MXI2X1 U1578 ( .A(n1248), .B(n1249), .S0(n1371), .Y(blockdata[27]) );
  MXI4X1 U1579 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n1439), .S1(n1404), .Y(n1249) );
  MXI4X1 U1580 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n1439), .S1(n1404), .Y(n1248) );
  MXI2X1 U1581 ( .A(n1246), .B(n1247), .S0(n1371), .Y(blockdata[28]) );
  MXI4X1 U1582 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n1439), .S1(n1404), .Y(n1247) );
  MXI4X1 U1583 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n1439), .S1(n1404), .Y(n1246) );
  MXI2X1 U1584 ( .A(n1244), .B(n1245), .S0(n1371), .Y(blockdata[29]) );
  MXI4X1 U1585 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n1439), .S1(n1404), .Y(n1245) );
  MXI4X1 U1586 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n1439), .S1(n1404), .Y(n1244) );
  MXI2X1 U1587 ( .A(n1242), .B(n1243), .S0(n1371), .Y(blockdata[30]) );
  MXI4X1 U1588 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n1439), .S1(n1404), .Y(n1243) );
  MXI4X1 U1589 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n1439), .S1(n1404), .Y(n1242) );
  MXI2X1 U1590 ( .A(n1240), .B(n1241), .S0(n1371), .Y(blockdata[31]) );
  MXI4X1 U1591 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n1438), .S1(n1404), .Y(n1241) );
  MXI4X1 U1592 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n1439), .S1(n1404), .Y(n1240) );
  MXI2X1 U1593 ( .A(n1282), .B(n1283), .S0(n1372), .Y(blockdata[10]) );
  MXI2X1 U1594 ( .A(n1280), .B(n1281), .S0(n1372), .Y(blockdata[11]) );
  MXI2X1 U1595 ( .A(n1278), .B(n1279), .S0(n1372), .Y(blockdata[12]) );
  MXI4X1 U1596 ( .A(\block[4][12] ), .B(\block[5][12] ), .C(\block[6][12] ), 
        .D(\block[7][12] ), .S0(n1441), .S1(n1407), .Y(n1279) );
  MXI4X1 U1597 ( .A(\block[0][12] ), .B(\block[1][12] ), .C(\block[2][12] ), 
        .D(\block[3][12] ), .S0(n1441), .S1(n1407), .Y(n1278) );
  MXI4XL U1598 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n1443), .S1(n1409), .Y(n1301) );
  MXI4XL U1599 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n1443), .S1(n1409), .Y(n1300) );
  MXI4XL U1600 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n1443), .S1(n1409), .Y(n1299) );
  MXI4XL U1601 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n1443), .S1(n1409), .Y(n1298) );
  MXI4XL U1602 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n1443), .S1(n1408), .Y(n1297) );
  MXI4XL U1603 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n1443), .S1(n1408), .Y(n1296) );
  MXI4XL U1604 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n1443), .S1(n1408), .Y(n1295) );
  MXI4XL U1605 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n1443), .S1(n1408), .Y(n1294) );
  MXI4X1 U1606 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n1442), .S1(n1408), .Y(n1293) );
  MXI4XL U1607 ( .A(\block[0][5] ), .B(\block[1][5] ), .C(\block[2][5] ), .D(
        \block[3][5] ), .S0(n1443), .S1(n1408), .Y(n1292) );
  MXI4X1 U1608 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n1442), .S1(n1408), .Y(n1291) );
  MXI4X1 U1609 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n1442), .S1(n1408), .Y(n1290) );
  MXI2XL U1610 ( .A(n1288), .B(n1289), .S0(n1373), .Y(blockdata[7]) );
  MXI4X1 U1611 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n1442), .S1(n1408), .Y(n1289) );
  MXI4X1 U1612 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n1442), .S1(n1408), .Y(n1288) );
  MXI2X1 U1613 ( .A(n1094), .B(n1095), .S0(n1367), .Y(blockdata[104]) );
  MXI4X1 U1614 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n1427), .S1(n1392), .Y(n1095) );
  MXI4X1 U1615 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n1427), .S1(n1392), .Y(n1094) );
  MXI2X1 U1616 ( .A(n1092), .B(n1093), .S0(n1366), .Y(blockdata[105]) );
  MXI4X1 U1617 ( .A(\block[4][105] ), .B(\block[5][105] ), .C(\block[6][105] ), 
        .D(\block[7][105] ), .S0(n1427), .S1(n1391), .Y(n1093) );
  MXI4X1 U1618 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n1427), .S1(n1391), .Y(n1092) );
  MXI2X1 U1619 ( .A(n1090), .B(n1091), .S0(n1366), .Y(blockdata[106]) );
  MXI4X1 U1620 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n1427), .S1(n1391), .Y(n1091) );
  MXI4X1 U1621 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n1427), .S1(n1391), .Y(n1090) );
  MXI2X1 U1622 ( .A(n1088), .B(n1089), .S0(n1366), .Y(blockdata[107]) );
  MXI4X1 U1623 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n1427), .S1(n1391), .Y(n1089) );
  MXI4X1 U1624 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n1427), .S1(n1391), .Y(n1088) );
  MXI2X1 U1625 ( .A(n1086), .B(n1087), .S0(n1366), .Y(blockdata[108]) );
  MXI4X1 U1626 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n1427), .S1(n1391), .Y(n1087) );
  MXI4X1 U1627 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n1427), .S1(n1391), .Y(n1086) );
  MXI2X1 U1628 ( .A(n1210), .B(n1211), .S0(n1366), .Y(blockdata[46]) );
  MXI4X1 U1629 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n1436), .S1(n1401), .Y(n1211) );
  MXI4X1 U1630 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n1436), .S1(n1401), .Y(n1210) );
  MXI2X1 U1631 ( .A(n1208), .B(n1209), .S0(n1366), .Y(blockdata[47]) );
  MXI4X1 U1632 ( .A(\block[4][47] ), .B(\block[5][47] ), .C(\block[6][47] ), 
        .D(\block[7][47] ), .S0(n1436), .S1(n1401), .Y(n1209) );
  MXI4X1 U1633 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n1436), .S1(n1401), .Y(n1208) );
  MXI2X1 U1634 ( .A(n1206), .B(n1207), .S0(n1366), .Y(blockdata[48]) );
  MXI4X1 U1635 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n1436), .S1(n1401), .Y(n1207) );
  MXI4X1 U1636 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n1436), .S1(n1401), .Y(n1206) );
  MXI2X1 U1637 ( .A(n1204), .B(n1205), .S0(n1366), .Y(blockdata[49]) );
  MXI4X1 U1638 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n1436), .S1(n1401), .Y(n1205) );
  MXI4X1 U1639 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n1436), .S1(n1401), .Y(n1204) );
  MXI2X1 U1640 ( .A(n1202), .B(n1203), .S0(n1366), .Y(blockdata[50]) );
  MXI4X1 U1641 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n1436), .S1(n1401), .Y(n1203) );
  MXI4X1 U1642 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n1436), .S1(n1401), .Y(n1202) );
  MXI2X1 U1643 ( .A(n1200), .B(n1201), .S0(n1366), .Y(blockdata[51]) );
  MXI4X1 U1644 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n1435), .S1(n1400), .Y(n1201) );
  MXI4X1 U1645 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n1435), .S1(n1400), .Y(n1200) );
  MXI2X1 U1646 ( .A(n1198), .B(n1199), .S0(n1366), .Y(blockdata[52]) );
  MXI4X1 U1647 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n1435), .S1(n1400), .Y(n1199) );
  MXI4X1 U1648 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n1435), .S1(n1400), .Y(n1198) );
  MXI2X1 U1649 ( .A(n1196), .B(n1197), .S0(n1366), .Y(blockdata[53]) );
  MXI4X1 U1650 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n1435), .S1(n1400), .Y(n1197) );
  MXI4X1 U1651 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n1435), .S1(n1400), .Y(n1196) );
  MXI2X1 U1652 ( .A(n1194), .B(n1195), .S0(n1366), .Y(blockdata[54]) );
  MXI4X1 U1653 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n1435), .S1(n1400), .Y(n1195) );
  MXI4X1 U1654 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n1435), .S1(n1400), .Y(n1194) );
  MXI2X1 U1655 ( .A(n1192), .B(n1193), .S0(n1366), .Y(blockdata[55]) );
  MXI4X1 U1656 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n1435), .S1(n1400), .Y(n1193) );
  MXI4X1 U1657 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n1435), .S1(n1400), .Y(n1192) );
  MXI2X1 U1658 ( .A(n1238), .B(n1239), .S0(n1371), .Y(blockdata[32]) );
  MXI4X1 U1659 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n1438), .S1(n1404), .Y(n1239) );
  MXI4X1 U1660 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n1438), .S1(n1404), .Y(n1238) );
  MXI2X1 U1661 ( .A(n1228), .B(n1229), .S0(n1370), .Y(blockdata[37]) );
  MXI4X1 U1662 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n1438), .S1(n1403), .Y(n1229) );
  MXI4X1 U1663 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n1438), .S1(n1403), .Y(n1228) );
  MXI2X1 U1664 ( .A(n1136), .B(n1137), .S0(n1368), .Y(blockdata[83]) );
  MXI4X1 U1665 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n1430), .S1(n1395), .Y(n1137) );
  MXI4X1 U1666 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n1431), .S1(n1395), .Y(n1136) );
  MXI2X1 U1667 ( .A(n1134), .B(n1135), .S0(n1368), .Y(blockdata[84]) );
  MXI4X1 U1668 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n1430), .S1(n1395), .Y(n1135) );
  MXI4X1 U1669 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n1430), .S1(n1395), .Y(n1134) );
  MXI2X1 U1670 ( .A(n1132), .B(n1133), .S0(n1368), .Y(blockdata[85]) );
  MXI4X1 U1671 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n1430), .S1(n1395), .Y(n1133) );
  MXI4X1 U1672 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n1430), .S1(n1395), .Y(n1132) );
  MXI2X1 U1673 ( .A(n1130), .B(n1131), .S0(n1368), .Y(blockdata[86]) );
  MXI4X1 U1674 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n1430), .S1(n1395), .Y(n1131) );
  MXI4X1 U1675 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n1430), .S1(n1395), .Y(n1130) );
  MXI2X1 U1676 ( .A(n1128), .B(n1129), .S0(n1368), .Y(blockdata[87]) );
  MXI4X1 U1677 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n1430), .S1(n1394), .Y(n1129) );
  MXI4X1 U1678 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n1430), .S1(n1394), .Y(n1128) );
  MXI2X1 U1679 ( .A(n1174), .B(n1175), .S0(n1370), .Y(blockdata[64]) );
  MXI4X1 U1680 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n1433), .S1(n1398), .Y(n1175) );
  MXI4X1 U1681 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n1433), .S1(n1398), .Y(n1174) );
  MXI2X1 U1682 ( .A(n1172), .B(n1173), .S0(n1370), .Y(blockdata[65]) );
  MXI4X1 U1683 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n1433), .S1(n1398), .Y(n1173) );
  MXI4X1 U1684 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n1433), .S1(n1398), .Y(n1172) );
  MXI2X1 U1685 ( .A(n1170), .B(n1171), .S0(n1370), .Y(blockdata[66]) );
  MXI4X1 U1686 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n1433), .S1(n1398), .Y(n1171) );
  MXI4X1 U1687 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n1433), .S1(n1398), .Y(n1170) );
  MXI2X1 U1688 ( .A(n1168), .B(n1169), .S0(n1370), .Y(blockdata[67]) );
  MXI4X1 U1689 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n1433), .S1(n1398), .Y(n1169) );
  MXI4X1 U1690 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n1433), .S1(n1398), .Y(n1168) );
  MXI2X1 U1691 ( .A(n1166), .B(n1167), .S0(n1370), .Y(blockdata[68]) );
  MXI4X1 U1692 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n1433), .S1(n1398), .Y(n1167) );
  MXI4X1 U1693 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n1433), .S1(n1398), .Y(n1166) );
  MXI2X1 U1694 ( .A(n1164), .B(n1165), .S0(n1369), .Y(blockdata[69]) );
  MXI4X1 U1695 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n1433), .S1(n1397), .Y(n1165) );
  MXI4X1 U1696 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n1433), .S1(n1397), .Y(n1164) );
  MXI2X1 U1697 ( .A(n1162), .B(n1163), .S0(n1369), .Y(blockdata[70]) );
  MXI4X1 U1698 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n1432), .S1(n1397), .Y(n1163) );
  MXI4X1 U1699 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n1433), .S1(n1397), .Y(n1162) );
  MXI2X1 U1700 ( .A(n1110), .B(n1111), .S0(n1367), .Y(blockdata[96]) );
  MXI4X1 U1701 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n1428), .S1(n1393), .Y(n1111) );
  MXI4X1 U1702 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n1429), .S1(n1393), .Y(n1110) );
  MXI2X1 U1703 ( .A(n1108), .B(n1109), .S0(n1367), .Y(blockdata[97]) );
  MXI4X1 U1704 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n1428), .S1(n1393), .Y(n1109) );
  MXI4X1 U1705 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n1428), .S1(n1393), .Y(n1108) );
  MXI2X1 U1706 ( .A(n1106), .B(n1107), .S0(n1367), .Y(blockdata[98]) );
  MXI4X1 U1707 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n1428), .S1(n1393), .Y(n1107) );
  MXI4X1 U1708 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n1428), .S1(n1393), .Y(n1106) );
  MXI2X1 U1709 ( .A(n1104), .B(n1105), .S0(n1367), .Y(blockdata[99]) );
  MXI4X1 U1710 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n1428), .S1(n1392), .Y(n1105) );
  MXI4X1 U1711 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n1428), .S1(n1392), .Y(n1104) );
  MXI2X1 U1712 ( .A(n1102), .B(n1103), .S0(n1367), .Y(blockdata[100]) );
  MXI4X1 U1713 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n1428), .S1(n1392), .Y(n1103) );
  MXI4X1 U1714 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n1428), .S1(n1392), .Y(n1102) );
  MXI2X1 U1715 ( .A(n1100), .B(n1101), .S0(n1367), .Y(blockdata[101]) );
  MXI4X1 U1716 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n1428), .S1(n1392), .Y(n1101) );
  MXI4X1 U1717 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n1428), .S1(n1392), .Y(n1100) );
  MXI2X1 U1718 ( .A(n1098), .B(n1099), .S0(n1367), .Y(blockdata[102]) );
  MXI4X1 U1719 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n1428), .S1(n1392), .Y(n1099) );
  MXI4X1 U1720 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n1428), .S1(n1392), .Y(n1098) );
  MXI2X1 U1721 ( .A(n1096), .B(n1097), .S0(n1367), .Y(blockdata[103]) );
  MXI4X1 U1722 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n1427), .S1(n1392), .Y(n1097) );
  MXI4X1 U1723 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n1427), .S1(n1392), .Y(n1096) );
  MXI2X1 U1724 ( .A(n1190), .B(n1191), .S0(n1366), .Y(blockdata[56]) );
  MXI4X1 U1725 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n1435), .S1(n1400), .Y(n1191) );
  MXI4X1 U1726 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n1435), .S1(n1400), .Y(n1190) );
  MXI2X1 U1727 ( .A(n1188), .B(n1189), .S0(n1370), .Y(blockdata[57]) );
  MXI4X1 U1728 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n1434), .S1(n1399), .Y(n1189) );
  MXI4X1 U1729 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n1435), .S1(n1399), .Y(n1188) );
  MXI2X1 U1730 ( .A(n1186), .B(n1187), .S0(n1370), .Y(blockdata[58]) );
  MXI4X1 U1731 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n1434), .S1(n1399), .Y(n1187) );
  MXI4X1 U1732 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n1434), .S1(n1399), .Y(n1186) );
  MXI2X1 U1733 ( .A(n1184), .B(n1185), .S0(n1370), .Y(blockdata[59]) );
  MXI4X1 U1734 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n1434), .S1(n1399), .Y(n1185) );
  MXI4X1 U1735 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n1434), .S1(n1399), .Y(n1184) );
  MXI2X1 U1736 ( .A(n1182), .B(n1183), .S0(n1370), .Y(blockdata[60]) );
  MXI4X1 U1737 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n1434), .S1(n1399), .Y(n1183) );
  MXI4X1 U1738 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n1434), .S1(n1399), .Y(n1182) );
  MXI2X1 U1739 ( .A(n1180), .B(n1181), .S0(n1370), .Y(blockdata[61]) );
  MXI4X1 U1740 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n1434), .S1(n1399), .Y(n1181) );
  MXI4X1 U1741 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n1434), .S1(n1399), .Y(n1180) );
  MXI2X1 U1742 ( .A(n1178), .B(n1179), .S0(n1370), .Y(blockdata[62]) );
  MXI4X1 U1743 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n1434), .S1(n1399), .Y(n1179) );
  MXI4X1 U1744 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n1434), .S1(n1399), .Y(n1178) );
  MXI2X1 U1745 ( .A(n1176), .B(n1177), .S0(n1370), .Y(blockdata[63]) );
  MXI4X1 U1746 ( .A(\block[4][63] ), .B(\block[5][63] ), .C(\block[6][63] ), 
        .D(\block[7][63] ), .S0(n1434), .S1(n1398), .Y(n1177) );
  MXI4X1 U1747 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n1434), .S1(n1398), .Y(n1176) );
  MXI2X1 U1748 ( .A(n1126), .B(n1127), .S0(n1368), .Y(blockdata[88]) );
  MXI4X1 U1749 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n1430), .S1(n1394), .Y(n1127) );
  MXI4X1 U1750 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n1430), .S1(n1394), .Y(n1126) );
  MXI2X1 U1751 ( .A(n1124), .B(n1125), .S0(n1368), .Y(blockdata[89]) );
  MXI4X1 U1752 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n1430), .S1(n1394), .Y(n1125) );
  MXI4X1 U1753 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n1430), .S1(n1394), .Y(n1124) );
  MXI2X1 U1754 ( .A(n1122), .B(n1123), .S0(n1368), .Y(blockdata[90]) );
  MXI4X1 U1755 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n1429), .S1(n1394), .Y(n1123) );
  MXI4X1 U1756 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n1429), .S1(n1394), .Y(n1122) );
  MXI2X1 U1757 ( .A(n1120), .B(n1121), .S0(n1368), .Y(blockdata[91]) );
  MXI4X1 U1758 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n1429), .S1(n1394), .Y(n1121) );
  MXI4X1 U1759 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n1429), .S1(n1394), .Y(n1120) );
  MXI2X1 U1760 ( .A(n1118), .B(n1119), .S0(n1368), .Y(blockdata[92]) );
  MXI4X1 U1761 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n1429), .S1(n1394), .Y(n1119) );
  MXI4X1 U1762 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n1429), .S1(n1394), .Y(n1118) );
  MXI2X1 U1763 ( .A(n1116), .B(n1117), .S0(n1367), .Y(blockdata[93]) );
  MXI4X1 U1764 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n1429), .S1(n1393), .Y(n1117) );
  MXI4X1 U1765 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n1429), .S1(n1393), .Y(n1116) );
  MXI2X1 U1766 ( .A(n1114), .B(n1115), .S0(n1367), .Y(blockdata[94]) );
  MXI4X1 U1767 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), 
        .D(\block[7][94] ), .S0(n1429), .S1(n1393), .Y(n1115) );
  MXI4X1 U1768 ( .A(\block[0][94] ), .B(\block[1][94] ), .C(\block[2][94] ), 
        .D(\block[3][94] ), .S0(n1429), .S1(n1393), .Y(n1114) );
  MXI2X1 U1769 ( .A(n1112), .B(n1113), .S0(n1367), .Y(blockdata[95]) );
  MXI4X1 U1770 ( .A(\block[4][95] ), .B(\block[5][95] ), .C(\block[6][95] ), 
        .D(\block[7][95] ), .S0(n1429), .S1(n1393), .Y(n1113) );
  MXI4X1 U1771 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n1429), .S1(n1393), .Y(n1112) );
  MXI2XL U1772 ( .A(n1286), .B(n1287), .S0(n1373), .Y(blockdata[8]) );
  MXI4X1 U1773 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n1442), .S1(n1408), .Y(n1287) );
  MXI4X1 U1774 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n1442), .S1(n1408), .Y(n1286) );
  MXI2X1 U1775 ( .A(n1284), .B(n1285), .S0(n1372), .Y(blockdata[9]) );
  MXI2XL U1776 ( .A(n1302), .B(n1303), .S0(n1373), .Y(blockdata[0]) );
  MXI4XL U1777 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n1443), .S1(n1409), .Y(n1302) );
  MXI4XL U1778 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n1443), .S1(n1409), .Y(n1303) );
  MXI2X1 U1779 ( .A(n1066), .B(n1067), .S0(n1365), .Y(blockdata[118]) );
  MXI2X1 U1780 ( .A(n1064), .B(n1065), .S0(n1365), .Y(blockdata[119]) );
  MXI2X1 U1781 ( .A(n1062), .B(n1063), .S0(n1365), .Y(blockdata[120]) );
  MXI2X1 U1782 ( .A(n1060), .B(n1061), .S0(n1365), .Y(blockdata[121]) );
  MXI2XL U1783 ( .A(n1084), .B(n1085), .S0(n1366), .Y(blockdata[109]) );
  MXI4XL U1784 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n1427), .S1(n1391), .Y(n1084) );
  MXI4XL U1785 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n1426), .S1(n1391), .Y(n1085) );
  MXI2XL U1786 ( .A(n1082), .B(n1083), .S0(n1366), .Y(blockdata[110]) );
  MXI4XL U1787 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n1426), .S1(n1391), .Y(n1082) );
  MXI4XL U1788 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n1426), .S1(n1391), .Y(n1083) );
  MXI2XL U1789 ( .A(n1080), .B(n1081), .S0(n1366), .Y(blockdata[111]) );
  MXI4X1 U1790 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n1426), .S1(n1390), .Y(n1080) );
  MXI4X1 U1791 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n1426), .S1(n1390), .Y(n1081) );
  MXI2XL U1792 ( .A(n1078), .B(n1079), .S0(n1366), .Y(blockdata[112]) );
  MXI4X1 U1793 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n1426), .S1(n1390), .Y(n1078) );
  MXI4X1 U1794 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n1426), .S1(n1390), .Y(n1079) );
  MXI2XL U1795 ( .A(n1076), .B(n1077), .S0(n1366), .Y(blockdata[113]) );
  MXI4X1 U1796 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n1426), .S1(n1390), .Y(n1076) );
  MXI4X1 U1797 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n1426), .S1(n1390), .Y(n1077) );
  MXI2XL U1798 ( .A(n1074), .B(n1075), .S0(n1366), .Y(blockdata[114]) );
  MXI4X1 U1799 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n1426), .S1(n1390), .Y(n1074) );
  MXI4X1 U1800 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n1426), .S1(n1390), .Y(n1075) );
  MXI2XL U1801 ( .A(n1072), .B(n1073), .S0(n1366), .Y(blockdata[115]) );
  MXI4X1 U1802 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n1426), .S1(n1390), .Y(n1072) );
  MXI4X1 U1803 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n1426), .S1(n1390), .Y(n1073) );
  MXI2XL U1804 ( .A(n1070), .B(n1071), .S0(n1366), .Y(blockdata[116]) );
  MXI4X1 U1805 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n1430), .S1(n1390), .Y(n1070) );
  MXI4X1 U1806 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n1442), .S1(n1390), .Y(n1071) );
  MXI2X1 U1807 ( .A(n1068), .B(n1069), .S0(n1365), .Y(blockdata[117]) );
  MXI2X1 U1808 ( .A(n1058), .B(n1059), .S0(n1365), .Y(blockdata[122]) );
  MXI4X1 U1809 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n1425), .S1(n1389), .Y(n1059) );
  MXI2XL U1810 ( .A(n1222), .B(n1223), .S0(n1366), .Y(blockdata[40]) );
  MXI4X1 U1811 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n1437), .S1(n1402), .Y(n1222) );
  MXI4X1 U1812 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n1437), .S1(n1402), .Y(n1223) );
  MXI2XL U1813 ( .A(n1220), .B(n1221), .S0(n1366), .Y(blockdata[41]) );
  MXI4X1 U1814 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n1437), .S1(n1402), .Y(n1220) );
  MXI4X1 U1815 ( .A(\block[4][41] ), .B(\block[5][41] ), .C(\block[6][41] ), 
        .D(\block[7][41] ), .S0(n1437), .S1(n1402), .Y(n1221) );
  MXI2XL U1816 ( .A(n1218), .B(n1219), .S0(n1366), .Y(blockdata[42]) );
  MXI4X1 U1817 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n1437), .S1(n1402), .Y(n1218) );
  MXI4X1 U1818 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n1437), .S1(n1402), .Y(n1219) );
  MXI2XL U1819 ( .A(n1216), .B(n1217), .S0(n1366), .Y(blockdata[43]) );
  MXI4X1 U1820 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n1437), .S1(n1402), .Y(n1216) );
  MXI4X1 U1821 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n1437), .S1(n1402), .Y(n1217) );
  MXI4XL U1822 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n1436), .S1(n1402), .Y(n1215) );
  MXI2XL U1823 ( .A(n1212), .B(n1213), .S0(n1366), .Y(blockdata[45]) );
  MXI4XL U1824 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n1436), .S1(n1401), .Y(n1212) );
  MXI4XL U1825 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n1436), .S1(n1401), .Y(n1213) );
  MXI2XL U1826 ( .A(n1236), .B(n1237), .S0(n1366), .Y(blockdata[33]) );
  MXI4XL U1827 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n1438), .S1(n1403), .Y(n1236) );
  MXI4XL U1828 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n1438), .S1(n1403), .Y(n1237) );
  MXI2XL U1829 ( .A(n1234), .B(n1235), .S0(n1366), .Y(blockdata[34]) );
  MXI4XL U1830 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n1438), .S1(n1403), .Y(n1234) );
  MXI4XL U1831 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n1438), .S1(n1403), .Y(n1235) );
  MXI2XL U1832 ( .A(n1232), .B(n1233), .S0(n1366), .Y(blockdata[35]) );
  MXI4XL U1833 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n1438), .S1(n1403), .Y(n1232) );
  MXI4XL U1834 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n1438), .S1(n1403), .Y(n1233) );
  MXI2XL U1835 ( .A(n1230), .B(n1231), .S0(n1366), .Y(blockdata[36]) );
  MXI4XL U1836 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n1438), .S1(n1403), .Y(n1230) );
  MXI4XL U1837 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n1438), .S1(n1403), .Y(n1231) );
  MXI2XL U1838 ( .A(n1226), .B(n1227), .S0(n1366), .Y(blockdata[38]) );
  MXI4XL U1839 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n1437), .S1(n1403), .Y(n1226) );
  MXI4XL U1840 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n1437), .S1(n1403), .Y(n1227) );
  MXI2XL U1841 ( .A(n1224), .B(n1225), .S0(n1370), .Y(blockdata[39]) );
  MXI2XL U1842 ( .A(n1158), .B(n1159), .S0(n1369), .Y(blockdata[72]) );
  MXI4XL U1843 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n1432), .S1(n1397), .Y(n1158) );
  MXI4XL U1844 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n1432), .S1(n1397), .Y(n1159) );
  MXI2XL U1845 ( .A(n1156), .B(n1157), .S0(n1369), .Y(blockdata[73]) );
  MXI4XL U1846 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n1432), .S1(n1397), .Y(n1156) );
  MXI4XL U1847 ( .A(\block[4][73] ), .B(\block[5][73] ), .C(\block[6][73] ), 
        .D(\block[7][73] ), .S0(n1432), .S1(n1397), .Y(n1157) );
  MXI2XL U1848 ( .A(n1154), .B(n1155), .S0(n1369), .Y(blockdata[74]) );
  MXI4XL U1849 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n1432), .S1(n1397), .Y(n1154) );
  MXI4XL U1850 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n1432), .S1(n1397), .Y(n1155) );
  MXI2XL U1851 ( .A(n1152), .B(n1153), .S0(n1369), .Y(blockdata[75]) );
  MXI4XL U1852 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n1432), .S1(n1396), .Y(n1152) );
  MXI4XL U1853 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n1432), .S1(n1396), .Y(n1153) );
  MXI2XL U1854 ( .A(n1150), .B(n1151), .S0(n1369), .Y(blockdata[76]) );
  MXI4XL U1855 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n1432), .S1(n1396), .Y(n1150) );
  MXI4XL U1856 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n1432), .S1(n1396), .Y(n1151) );
  MXI2XL U1857 ( .A(n1148), .B(n1149), .S0(n1369), .Y(blockdata[77]) );
  MXI4XL U1858 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n1431), .S1(n1396), .Y(n1148) );
  MXI4XL U1859 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n1431), .S1(n1396), .Y(n1149) );
  MXI2XL U1860 ( .A(n1146), .B(n1147), .S0(n1369), .Y(blockdata[78]) );
  MXI4XL U1861 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n1431), .S1(n1396), .Y(n1146) );
  MXI4XL U1862 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n1431), .S1(n1396), .Y(n1147) );
  MXI2XL U1863 ( .A(n1144), .B(n1145), .S0(n1369), .Y(blockdata[79]) );
  MXI4XL U1864 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n1431), .S1(n1396), .Y(n1144) );
  MXI4XL U1865 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n1431), .S1(n1396), .Y(n1145) );
  MXI2XL U1866 ( .A(n1142), .B(n1143), .S0(n1369), .Y(blockdata[80]) );
  MXI4XL U1867 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n1431), .S1(n1396), .Y(n1142) );
  MXI4XL U1868 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n1431), .S1(n1396), .Y(n1143) );
  MXI2XL U1869 ( .A(n1140), .B(n1141), .S0(n1368), .Y(blockdata[81]) );
  MXI4XL U1870 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n1431), .S1(n1395), .Y(n1140) );
  MXI4XL U1871 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n1431), .S1(n1395), .Y(n1141) );
  MXI2XL U1872 ( .A(n1138), .B(n1139), .S0(n1368), .Y(blockdata[82]) );
  MXI4XL U1873 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n1431), .S1(n1395), .Y(n1138) );
  MXI4XL U1874 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n1431), .S1(n1395), .Y(n1139) );
  MXI2XL U1875 ( .A(n1160), .B(n1161), .S0(n1369), .Y(blockdata[71]) );
  MXI4XL U1876 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n1432), .S1(n1397), .Y(n1160) );
  MXI4XL U1877 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n1432), .S1(n1397), .Y(n1161) );
  MXI2X1 U1878 ( .A(n1056), .B(n1057), .S0(n1365), .Y(blockdata[123]) );
  MXI4X1 U1879 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n1425), .S1(n1388), .Y(n1056) );
  MXI4X1 U1880 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n1425), .S1(n1388), .Y(n1057) );
  MXI2X1 U1881 ( .A(n1054), .B(n1055), .S0(n1365), .Y(blockdata[124]) );
  MXI4X1 U1882 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n1425), .S1(n1388), .Y(n1054) );
  MXI4X1 U1883 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n1425), .S1(n1388), .Y(n1055) );
  MXI2X1 U1884 ( .A(n1052), .B(n1053), .S0(n1365), .Y(blockdata[125]) );
  MXI4X1 U1885 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n1425), .S1(n1388), .Y(n1052) );
  MXI4X1 U1886 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n1425), .S1(n1388), .Y(n1053) );
  MXI2X1 U1887 ( .A(n1050), .B(n1051), .S0(n1365), .Y(blockdata[126]) );
  MXI4X1 U1888 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n1425), .S1(n1388), .Y(n1050) );
  MXI4X1 U1889 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n1425), .S1(n1388), .Y(n1051) );
  MXI2X1 U1890 ( .A(n1048), .B(n1049), .S0(n1365), .Y(blockdata[127]) );
  MXI4X1 U1891 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n1425), .S1(n1388), .Y(n1048) );
  MXI4X1 U1892 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n1425), .S1(n1388), .Y(n1049) );
  AO21XL U1893 ( .A0(mem_ready), .A1(n1948), .B0(valid), .Y(n1852) );
  MXI2X4 U1894 ( .A(n1304), .B(n1305), .S0(n1373), .Y(valid) );
  MXI2X4 U1895 ( .A(n1308), .B(n1309), .S0(n1373), .Y(tag[24]) );
  MXI2X4 U1896 ( .A(n1312), .B(n1313), .S0(n1374), .Y(tag[22]) );
  MXI2X4 U1897 ( .A(n1322), .B(n1323), .S0(n1374), .Y(tag[17]) );
  MXI2X4 U1898 ( .A(n1324), .B(n1325), .S0(n1374), .Y(tag[16]) );
  MXI2X4 U1899 ( .A(n1332), .B(n1333), .S0(n1374), .Y(tag[12]) );
  MXI2X4 U1900 ( .A(n1338), .B(n1339), .S0(n1375), .Y(tag[9]) );
  MXI2X4 U1901 ( .A(n1344), .B(n1345), .S0(n1375), .Y(tag[6]) );
  MXI2X4 U1902 ( .A(n1346), .B(n1347), .S0(n1375), .Y(tag[5]) );
  MXI2X4 U1903 ( .A(n1350), .B(n1351), .S0(n1375), .Y(tag[3]) );
  MXI2X4 U1904 ( .A(n1354), .B(n1355), .S0(n1375), .Y(tag[1]) );
  MXI2X4 U1905 ( .A(n1356), .B(n1357), .S0(n1375), .Y(tag[0]) );
  MXI4X4 U1906 ( .A(\blocktag[4][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[7][22] ), .S0(n1444), .S1(n1410), .Y(
        n1313) );
  MXI4X4 U1907 ( .A(\blocktag[0][22] ), .B(\blocktag[1][22] ), .C(
        \blocktag[2][22] ), .D(\blocktag[3][22] ), .S0(n1444), .S1(n118), .Y(
        n1312) );
  MXI4X4 U1908 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n119), .S1(n1411), .Y(
        n1322) );
  MXI4X4 U1909 ( .A(\blocktag[4][7] ), .B(\blocktag[5][7] ), .C(
        \blocktag[6][7] ), .D(\blocktag[7][7] ), .S0(n120), .S1(n1412), .Y(
        n1343) );
  MXI4X4 U1910 ( .A(\blocktag[0][7] ), .B(\blocktag[1][7] ), .C(
        \blocktag[2][7] ), .D(\blocktag[3][7] ), .S0(n120), .S1(n1412), .Y(
        n1342) );
  MXI4X4 U1911 ( .A(\blocktag[4][0] ), .B(\blocktag[5][0] ), .C(
        \blocktag[6][0] ), .D(\blocktag[7][0] ), .S0(n1447), .S1(n1413), .Y(
        n1357) );
  MXI4X4 U1912 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(
        \blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n1618), .S1(n1413), .Y(
        n1356) );
  AND2XL U1913 ( .A(n1626), .B(blockdata[33]), .Y(mem_wdata[33]) );
  AND2XL U1914 ( .A(n1625), .B(blockdata[71]), .Y(mem_wdata[71]) );
  AND2XL U1915 ( .A(n1624), .B(blockdata[109]), .Y(mem_wdata[109]) );
  AND2XL U1916 ( .A(n1626), .B(blockdata[34]), .Y(mem_wdata[34]) );
  AND2XL U1917 ( .A(n1625), .B(blockdata[72]), .Y(mem_wdata[72]) );
  AND2XL U1918 ( .A(n1624), .B(blockdata[110]), .Y(mem_wdata[110]) );
  AND2XL U1919 ( .A(n1626), .B(blockdata[35]), .Y(mem_wdata[35]) );
  AND2XL U1920 ( .A(n1625), .B(blockdata[73]), .Y(mem_wdata[73]) );
  AND2XL U1921 ( .A(n1624), .B(blockdata[111]), .Y(mem_wdata[111]) );
  AND2XL U1922 ( .A(n1626), .B(blockdata[36]), .Y(mem_wdata[36]) );
  AND2XL U1923 ( .A(n1625), .B(blockdata[74]), .Y(mem_wdata[74]) );
  AND2XL U1924 ( .A(n1624), .B(blockdata[112]), .Y(mem_wdata[112]) );
  AND2XL U1925 ( .A(mem_write), .B(blockdata[0]), .Y(mem_wdata[0]) );
  AND2XL U1926 ( .A(n1626), .B(blockdata[38]), .Y(mem_wdata[38]) );
  AND2XL U1927 ( .A(n1625), .B(blockdata[75]), .Y(mem_wdata[75]) );
  AND2XL U1928 ( .A(n1624), .B(blockdata[113]), .Y(mem_wdata[113]) );
  AND2XL U1929 ( .A(mem_write), .B(blockdata[121]), .Y(mem_wdata[121]) );
  AND2XL U1930 ( .A(n1626), .B(blockdata[39]), .Y(mem_wdata[39]) );
  AND2XL U1931 ( .A(n1625), .B(blockdata[76]), .Y(mem_wdata[76]) );
  AND2XL U1932 ( .A(n1624), .B(blockdata[114]), .Y(mem_wdata[114]) );
  AND2XL U1933 ( .A(mem_write), .B(blockdata[122]), .Y(mem_wdata[122]) );
  AND2XL U1934 ( .A(n1626), .B(blockdata[40]), .Y(mem_wdata[40]) );
  AND2XL U1935 ( .A(n1625), .B(blockdata[77]), .Y(mem_wdata[77]) );
  AND2XL U1936 ( .A(n1624), .B(blockdata[115]), .Y(mem_wdata[115]) );
  AND2XL U1937 ( .A(mem_write), .B(blockdata[123]), .Y(mem_wdata[123]) );
  AND2XL U1938 ( .A(n1626), .B(blockdata[41]), .Y(mem_wdata[41]) );
  AND2XL U1939 ( .A(n1625), .B(blockdata[78]), .Y(mem_wdata[78]) );
  AND2XL U1940 ( .A(n1624), .B(blockdata[116]), .Y(mem_wdata[116]) );
  AND2XL U1941 ( .A(mem_write), .B(blockdata[124]), .Y(mem_wdata[124]) );
  AND2XL U1942 ( .A(n1626), .B(blockdata[42]), .Y(mem_wdata[42]) );
  AND2XL U1943 ( .A(n1625), .B(blockdata[79]), .Y(mem_wdata[79]) );
  AND2XL U1944 ( .A(n1624), .B(blockdata[117]), .Y(mem_wdata[117]) );
  AND2XL U1945 ( .A(mem_write), .B(blockdata[125]), .Y(mem_wdata[125]) );
  AND2XL U1946 ( .A(n1626), .B(blockdata[43]), .Y(mem_wdata[43]) );
  AND2XL U1947 ( .A(n1625), .B(blockdata[80]), .Y(mem_wdata[80]) );
  AND2XL U1948 ( .A(n1624), .B(blockdata[118]), .Y(mem_wdata[118]) );
  AND2XL U1949 ( .A(mem_write), .B(blockdata[126]), .Y(mem_wdata[126]) );
  AND2XL U1950 ( .A(n1626), .B(blockdata[44]), .Y(mem_wdata[44]) );
  AND2XL U1951 ( .A(n1625), .B(blockdata[81]), .Y(mem_wdata[81]) );
  AND2XL U1952 ( .A(n1624), .B(blockdata[119]), .Y(mem_wdata[119]) );
  AND2XL U1953 ( .A(mem_write), .B(blockdata[127]), .Y(mem_wdata[127]) );
  AND2XL U1954 ( .A(n1626), .B(blockdata[45]), .Y(mem_wdata[45]) );
  AND2XL U1955 ( .A(n1625), .B(blockdata[82]), .Y(mem_wdata[82]) );
  AND2XL U1956 ( .A(n1624), .B(blockdata[120]), .Y(mem_wdata[120]) );
  AND3X8 U1957 ( .A(n1657), .B(n1656), .C(n1655), .Y(n1658) );
  CLKXOR2X2 U1958 ( .A(n1869), .B(proc_addr[25]), .Y(n1654) );
  OAI221X4 U1959 ( .A0(n1472), .A1(n1831), .B0(n1849), .B1(n2009), .C0(n1830), 
        .Y(block_next[9]) );
  NAND3BXL U1960 ( .AN(proc_addr[0]), .B(n1955), .C(n1958), .Y(n2123) );
  NAND3BXL U1961 ( .AN(n1959), .B(proc_addr[0]), .C(n1958), .Y(n2116) );
  NAND2X1 U1962 ( .A(proc_addr[0]), .B(proc_addr[1]), .Y(n1672) );
  OAI221X4 U1963 ( .A0(n1472), .A1(n1833), .B0(n1849), .B1(n2004), .C0(n1832), 
        .Y(block_next[8]) );
  XOR2X2 U1964 ( .A(n1905), .B(proc_addr[12]), .Y(n1647) );
  AOI2BB1X2 U1965 ( .A0N(n1666), .A1N(n8), .B0(n11), .Y(n1667) );
  CLKINVX3 U1966 ( .A(proc_read), .Y(n1669) );
  NAND2X2 U1967 ( .A(n1669), .B(n1954), .Y(n1948) );
  NAND4BBX4 U1968 ( .AN(n1676), .BN(n1675), .C(valid), .D(n1674), .Y(n1677) );
  OAI21X4 U1969 ( .A0(n1677), .A1(n16), .B0(n1948), .Y(n1853) );
  OAI221X2 U1970 ( .A0(n1464), .A1(n1985), .B0(n1839), .B1(n1465), .C0(n1779), 
        .Y(block_next[37]) );
  OAI221X2 U1971 ( .A0(n1472), .A1(n1835), .B0(n1849), .B1(n1999), .C0(n1834), 
        .Y(block_next[7]) );
  CLKINVX3 U1972 ( .A(n1852), .Y(n1944) );
  CLKINVX3 U1973 ( .A(n1856), .Y(n1946) );
  CLKINVX3 U1974 ( .A(n1858), .Y(blocktag_next[24]) );
  CLKINVX3 U1975 ( .A(n1861), .Y(blocktag_next[23]) );
  CLKINVX3 U1976 ( .A(n1864), .Y(blocktag_next[22]) );
  CLKINVX3 U1977 ( .A(n1867), .Y(blocktag_next[21]) );
  CLKINVX3 U1978 ( .A(n1870), .Y(blocktag_next[20]) );
  CLKINVX3 U1979 ( .A(n1873), .Y(blocktag_next[19]) );
  CLKINVX3 U1980 ( .A(n1875), .Y(blocktag_next[18]) );
  CLKINVX3 U1981 ( .A(n1878), .Y(blocktag_next[17]) );
  CLKINVX3 U1982 ( .A(n1881), .Y(blocktag_next[16]) );
  CLKINVX3 U1983 ( .A(n1883), .Y(blocktag_next[15]) );
  CLKINVX3 U1984 ( .A(n1885), .Y(blocktag_next[14]) );
  CLKINVX3 U1985 ( .A(n1888), .Y(blocktag_next[13]) );
  CLKINVX3 U1986 ( .A(n1891), .Y(blocktag_next[12]) );
  CLKINVX3 U1987 ( .A(n1894), .Y(blocktag_next[11]) );
  CLKINVX3 U1988 ( .A(n1897), .Y(blocktag_next[10]) );
  CLKINVX3 U1989 ( .A(n1900), .Y(blocktag_next[9]) );
  CLKINVX3 U1990 ( .A(n1903), .Y(blocktag_next[8]) );
  CLKINVX3 U1991 ( .A(n1906), .Y(blocktag_next[7]) );
  CLKINVX3 U1992 ( .A(n1909), .Y(blocktag_next[6]) );
  CLKINVX3 U1993 ( .A(n1912), .Y(blocktag_next[5]) );
  CLKINVX3 U1994 ( .A(n1915), .Y(blocktag_next[4]) );
  CLKINVX3 U1995 ( .A(n1918), .Y(blocktag_next[3]) );
  CLKINVX3 U1996 ( .A(n1920), .Y(blocktag_next[2]) );
  CLKINVX3 U1997 ( .A(n1923), .Y(blocktag_next[1]) );
  CLKINVX3 U1998 ( .A(n1927), .Y(blocktag_next[0]) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, \blocktag[7][24] , \blocktag[7][22] , \blocktag[7][21] ,
         \blocktag[7][20] , \blocktag[7][19] , \blocktag[7][17] ,
         \blocktag[7][12] , \blocktag[7][8] , \blocktag[7][3] ,
         \blocktag[7][0] , \blocktag[6][24] , \blocktag[6][22] ,
         \blocktag[6][21] , \blocktag[6][20] , \blocktag[6][19] ,
         \blocktag[6][17] , \blocktag[6][12] , \blocktag[6][8] ,
         \blocktag[6][3] , \blocktag[6][0] , \blocktag[5][24] ,
         \blocktag[5][22] , \blocktag[5][21] , \blocktag[5][20] ,
         \blocktag[5][19] , \blocktag[5][17] , \blocktag[5][12] ,
         \blocktag[5][8] , \blocktag[5][3] , \blocktag[5][0] ,
         \blocktag[4][24] , \blocktag[4][22] , \blocktag[4][21] ,
         \blocktag[4][20] , \blocktag[4][19] , \blocktag[4][17] ,
         \blocktag[4][12] , \blocktag[4][8] , \blocktag[4][3] ,
         \blocktag[4][0] , \blocktag[3][24] , \blocktag[3][21] ,
         \blocktag[3][20] , \blocktag[3][19] , \blocktag[3][18] ,
         \blocktag[3][17] , \blocktag[3][16] , \blocktag[3][13] ,
         \blocktag[3][12] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][7] , \blocktag[3][4] , \blocktag[3][3] ,
         \blocktag[3][1] , \blocktag[3][0] , \blocktag[2][24] ,
         \blocktag[2][21] , \blocktag[2][20] , \blocktag[2][19] ,
         \blocktag[2][18] , \blocktag[2][17] , \blocktag[2][16] ,
         \blocktag[2][13] , \blocktag[2][12] , \blocktag[2][11] ,
         \blocktag[2][10] , \blocktag[2][7] , \blocktag[2][4] ,
         \blocktag[2][3] , \blocktag[2][1] , \blocktag[2][0] ,
         \blocktag[1][24] , \blocktag[1][21] , \blocktag[1][20] ,
         \blocktag[1][19] , \blocktag[1][18] , \blocktag[1][17] ,
         \blocktag[1][16] , \blocktag[1][13] , \blocktag[1][12] ,
         \blocktag[1][11] , \blocktag[1][10] , \blocktag[1][7] ,
         \blocktag[1][4] , \blocktag[1][3] , \blocktag[1][1] ,
         \blocktag[1][0] , \blocktag[0][24] , \blocktag[0][21] ,
         \blocktag[0][20] , \blocktag[0][19] , \blocktag[0][18] ,
         \blocktag[0][17] , \blocktag[0][16] , \blocktag[0][13] ,
         \blocktag[0][12] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][7] , \blocktag[0][4] , \blocktag[0][3] ,
         \blocktag[0][1] , \blocktag[0][0] , \block[7][127] , \block[7][126] ,
         \block[7][125] , \block[7][124] , \block[7][123] , \block[7][122] ,
         \block[7][121] , \block[7][120] , \block[7][119] , \block[7][118] ,
         \block[7][117] , \block[7][116] , \block[7][115] , \block[7][114] ,
         \block[7][113] , \block[7][112] , \block[7][111] , \block[7][110] ,
         \block[7][109] , \block[7][108] , \block[7][107] , \block[7][106] ,
         \block[7][105] , \block[7][104] , \block[7][103] , \block[7][102] ,
         \block[7][101] , \block[7][100] , \block[7][99] , \block[7][98] ,
         \block[7][97] , \block[7][96] , \block[7][95] , \block[7][94] ,
         \block[7][93] , \block[7][92] , \block[7][91] , \block[7][90] ,
         \block[7][89] , \block[7][88] , \block[7][87] , \block[7][86] ,
         \block[7][85] , \block[7][84] , \block[7][83] , \block[7][82] ,
         \block[7][81] , \block[7][80] , \block[7][79] , \block[7][78] ,
         \block[7][77] , \block[7][76] , \block[7][75] , \block[7][74] ,
         \block[7][73] , \block[7][72] , \block[7][71] , \block[7][70] ,
         \block[7][69] , \block[7][68] , \block[7][67] , \block[7][66] ,
         \block[7][65] , \block[7][64] , \block[7][63] , \block[7][62] ,
         \block[7][61] , \block[7][60] , \block[7][59] , \block[7][58] ,
         \block[7][57] , \block[7][56] , \block[7][55] , \block[7][54] ,
         \block[7][53] , \block[7][52] , \block[7][51] , \block[7][50] ,
         \block[7][49] , \block[7][48] , \block[7][47] , \block[7][46] ,
         \block[7][45] , \block[7][44] , \block[7][43] , \block[7][42] ,
         \block[7][41] , \block[7][40] , \block[7][39] , \block[7][38] ,
         \block[7][37] , \block[7][36] , \block[7][35] , \block[7][34] ,
         \block[7][33] , \block[7][32] , \block[7][31] , \block[7][30] ,
         \block[7][29] , \block[7][28] , \block[7][27] , \block[7][26] ,
         \block[7][25] , \block[7][24] , \block[7][23] , \block[7][22] ,
         \block[7][21] , \block[7][20] , \block[7][19] , \block[7][18] ,
         \block[7][17] , \block[7][16] , \block[7][15] , \block[7][14] ,
         \block[7][13] , \block[7][12] , \block[7][11] , \block[7][10] ,
         \block[7][9] , \block[7][8] , \block[7][7] , \block[7][6] ,
         \block[7][5] , \block[7][4] , \block[7][3] , \block[7][2] ,
         \block[7][1] , \block[7][0] , \block[6][127] , \block[6][126] ,
         \block[6][125] , \block[6][124] , \block[6][123] , \block[6][122] ,
         \block[6][121] , \block[6][120] , \block[6][119] , \block[6][118] ,
         \block[6][117] , \block[6][116] , \block[6][115] , \block[6][114] ,
         \block[6][113] , \block[6][112] , \block[6][111] , \block[6][110] ,
         \block[6][109] , \block[6][108] , \block[6][107] , \block[6][106] ,
         \block[6][105] , \block[6][104] , \block[6][103] , \block[6][102] ,
         \block[6][101] , \block[6][100] , \block[6][99] , \block[6][98] ,
         \block[6][97] , \block[6][96] , \block[6][95] , \block[6][94] ,
         \block[6][93] , \block[6][92] , \block[6][91] , \block[6][90] ,
         \block[6][89] , \block[6][88] , \block[6][87] , \block[6][86] ,
         \block[6][85] , \block[6][84] , \block[6][83] , \block[6][82] ,
         \block[6][81] , \block[6][80] , \block[6][79] , \block[6][78] ,
         \block[6][77] , \block[6][76] , \block[6][75] , \block[6][74] ,
         \block[6][73] , \block[6][72] , \block[6][71] , \block[6][70] ,
         \block[6][69] , \block[6][68] , \block[6][67] , \block[6][66] ,
         \block[6][65] , \block[6][64] , \block[6][63] , \block[6][62] ,
         \block[6][61] , \block[6][60] , \block[6][59] , \block[6][58] ,
         \block[6][57] , \block[6][56] , \block[6][55] , \block[6][54] ,
         \block[6][53] , \block[6][52] , \block[6][51] , \block[6][50] ,
         \block[6][49] , \block[6][48] , \block[6][47] , \block[6][46] ,
         \block[6][45] , \block[6][44] , \block[6][43] , \block[6][42] ,
         \block[6][41] , \block[6][40] , \block[6][39] , \block[6][38] ,
         \block[6][37] , \block[6][36] , \block[6][35] , \block[6][34] ,
         \block[6][33] , \block[6][32] , \block[6][31] , \block[6][30] ,
         \block[6][29] , \block[6][28] , \block[6][27] , \block[6][26] ,
         \block[6][25] , \block[6][24] , \block[6][23] , \block[6][22] ,
         \block[6][21] , \block[6][20] , \block[6][19] , \block[6][18] ,
         \block[6][17] , \block[6][16] , \block[6][15] , \block[6][14] ,
         \block[6][13] , \block[6][12] , \block[6][11] , \block[6][10] ,
         \block[6][9] , \block[6][8] , \block[6][7] , \block[6][6] ,
         \block[6][5] , \block[6][4] , \block[6][3] , \block[6][2] ,
         \block[6][1] , \block[6][0] , \block[5][127] , \block[5][126] ,
         \block[5][125] , \block[5][124] , \block[5][123] , \block[5][122] ,
         \block[5][121] , \block[5][120] , \block[5][119] , \block[5][118] ,
         \block[5][117] , \block[5][116] , \block[5][115] , \block[5][114] ,
         \block[5][113] , \block[5][112] , \block[5][111] , \block[5][110] ,
         \block[5][109] , \block[5][108] , \block[5][107] , \block[5][106] ,
         \block[5][105] , \block[5][104] , \block[5][103] , \block[5][102] ,
         \block[5][101] , \block[5][100] , \block[5][99] , \block[5][98] ,
         \block[5][97] , \block[5][96] , \block[5][95] , \block[5][94] ,
         \block[5][93] , \block[5][92] , \block[5][91] , \block[5][90] ,
         \block[5][89] , \block[5][88] , \block[5][87] , \block[5][86] ,
         \block[5][85] , \block[5][84] , \block[5][83] , \block[5][82] ,
         \block[5][81] , \block[5][80] , \block[5][79] , \block[5][78] ,
         \block[5][77] , \block[5][76] , \block[5][75] , \block[5][74] ,
         \block[5][73] , \block[5][72] , \block[5][71] , \block[5][70] ,
         \block[5][69] , \block[5][68] , \block[5][67] , \block[5][66] ,
         \block[5][65] , \block[5][64] , \block[5][63] , \block[5][62] ,
         \block[5][61] , \block[5][60] , \block[5][59] , \block[5][58] ,
         \block[5][57] , \block[5][56] , \block[5][55] , \block[5][54] ,
         \block[5][53] , \block[5][52] , \block[5][51] , \block[5][50] ,
         \block[5][49] , \block[5][48] , \block[5][47] , \block[5][46] ,
         \block[5][45] , \block[5][44] , \block[5][43] , \block[5][42] ,
         \block[5][41] , \block[5][40] , \block[5][39] , \block[5][38] ,
         \block[5][37] , \block[5][36] , \block[5][35] , \block[5][34] ,
         \block[5][33] , \block[5][32] , \block[5][31] , \block[5][30] ,
         \block[5][29] , \block[5][28] , \block[5][27] , \block[5][26] ,
         \block[5][25] , \block[5][24] , \block[5][23] , \block[5][22] ,
         \block[5][21] , \block[5][20] , \block[5][19] , \block[5][18] ,
         \block[5][17] , \block[5][16] , \block[5][15] , \block[5][14] ,
         \block[5][13] , \block[5][12] , \block[5][11] , \block[5][10] ,
         \block[5][9] , \block[5][8] , \block[5][7] , \block[5][6] ,
         \block[5][5] , \block[5][4] , \block[5][3] , \block[5][2] ,
         \block[5][1] , \block[5][0] , \block[4][127] , \block[4][126] ,
         \block[4][125] , \block[4][124] , \block[4][123] , \block[4][122] ,
         \block[4][121] , \block[4][120] , \block[4][119] , \block[4][118] ,
         \block[4][117] , \block[4][116] , \block[4][115] , \block[4][114] ,
         \block[4][113] , \block[4][112] , \block[4][111] , \block[4][110] ,
         \block[4][109] , \block[4][108] , \block[4][107] , \block[4][106] ,
         \block[4][105] , \block[4][104] , \block[4][103] , \block[4][102] ,
         \block[4][101] , \block[4][100] , \block[4][99] , \block[4][98] ,
         \block[4][97] , \block[4][96] , \block[4][95] , \block[4][94] ,
         \block[4][93] , \block[4][92] , \block[4][91] , \block[4][90] ,
         \block[4][89] , \block[4][88] , \block[4][87] , \block[4][86] ,
         \block[4][85] , \block[4][84] , \block[4][83] , \block[4][82] ,
         \block[4][81] , \block[4][80] , \block[4][79] , \block[4][78] ,
         \block[4][77] , \block[4][76] , \block[4][75] , \block[4][74] ,
         \block[4][73] , \block[4][72] , \block[4][71] , \block[4][70] ,
         \block[4][69] , \block[4][68] , \block[4][67] , \block[4][66] ,
         \block[4][65] , \block[4][64] , \block[4][63] , \block[4][62] ,
         \block[4][61] , \block[4][60] , \block[4][59] , \block[4][58] ,
         \block[4][57] , \block[4][56] , \block[4][55] , \block[4][54] ,
         \block[4][53] , \block[4][52] , \block[4][51] , \block[4][50] ,
         \block[4][49] , \block[4][48] , \block[4][47] , \block[4][46] ,
         \block[4][45] , \block[4][44] , \block[4][43] , \block[4][42] ,
         \block[4][41] , \block[4][40] , \block[4][39] , \block[4][38] ,
         \block[4][37] , \block[4][36] , \block[4][35] , \block[4][34] ,
         \block[4][33] , \block[4][32] , \block[4][31] , \block[4][30] ,
         \block[4][29] , \block[4][28] , \block[4][27] , \block[4][26] ,
         \block[4][25] , \block[4][24] , \block[4][23] , \block[4][22] ,
         \block[4][21] , \block[4][20] , \block[4][19] , \block[4][18] ,
         \block[4][17] , \block[4][16] , \block[4][15] , \block[4][14] ,
         \block[4][13] , \block[4][12] , \block[4][11] , \block[4][10] ,
         \block[4][9] , \block[4][8] , \block[4][7] , \block[4][6] ,
         \block[4][5] , \block[4][4] , \block[4][3] , \block[4][2] ,
         \block[4][1] , \block[4][0] , \block[3][127] , \block[3][126] ,
         \block[3][125] , \block[3][124] , \block[3][123] , \block[3][122] ,
         \block[3][121] , \block[3][120] , \block[3][119] , \block[3][118] ,
         \block[3][117] , \block[3][116] , \block[3][115] , \block[3][114] ,
         \block[3][113] , \block[3][112] , \block[3][111] , \block[3][110] ,
         \block[3][109] , \block[3][108] , \block[3][107] , \block[3][106] ,
         \block[3][105] , \block[3][104] , \block[3][103] , \block[3][102] ,
         \block[3][101] , \block[3][100] , \block[3][99] , \block[3][98] ,
         \block[3][97] , \block[3][96] , \block[3][95] , \block[3][94] ,
         \block[3][93] , \block[3][92] , \block[3][91] , \block[3][90] ,
         \block[3][89] , \block[3][88] , \block[3][87] , \block[3][86] ,
         \block[3][85] , \block[3][84] , \block[3][83] , \block[3][82] ,
         \block[3][81] , \block[3][80] , \block[3][79] , \block[3][78] ,
         \block[3][77] , \block[3][76] , \block[3][75] , \block[3][74] ,
         \block[3][73] , \block[3][72] , \block[3][71] , \block[3][70] ,
         \block[3][69] , \block[3][68] , \block[3][67] , \block[3][66] ,
         \block[3][65] , \block[3][64] , \block[3][63] , \block[3][62] ,
         \block[3][61] , \block[3][60] , \block[3][59] , \block[3][58] ,
         \block[3][57] , \block[3][56] , \block[3][55] , \block[3][54] ,
         \block[3][53] , \block[3][52] , \block[3][51] , \block[3][50] ,
         \block[3][49] , \block[3][48] , \block[3][47] , \block[3][46] ,
         \block[3][45] , \block[3][44] , \block[3][43] , \block[3][42] ,
         \block[3][41] , \block[3][40] , \block[3][39] , \block[3][38] ,
         \block[3][37] , \block[3][36] , \block[3][35] , \block[3][34] ,
         \block[3][33] , \block[3][32] , \block[3][31] , \block[3][30] ,
         \block[3][29] , \block[3][28] , \block[3][27] , \block[3][26] ,
         \block[3][25] , \block[3][24] , \block[3][23] , \block[3][22] ,
         \block[3][21] , \block[3][20] , \block[3][19] , \block[3][18] ,
         \block[3][17] , \block[3][16] , \block[3][15] , \block[3][14] ,
         \block[3][13] , \block[3][12] , \block[3][11] , \block[3][10] ,
         \block[3][9] , \block[3][8] , \block[3][7] , \block[3][6] ,
         \block[3][5] , \block[3][4] , \block[3][3] , \block[3][2] ,
         \block[3][1] , \block[3][0] , \block[2][127] , \block[2][126] ,
         \block[2][125] , \block[2][124] , \block[2][123] , \block[2][122] ,
         \block[2][121] , \block[2][120] , \block[2][119] , \block[2][118] ,
         \block[2][117] , \block[2][116] , \block[2][115] , \block[2][114] ,
         \block[2][113] , \block[2][112] , \block[2][111] , \block[2][110] ,
         \block[2][109] , \block[2][108] , \block[2][107] , \block[2][106] ,
         \block[2][105] , \block[2][104] , \block[2][103] , \block[2][102] ,
         \block[2][101] , \block[2][100] , \block[2][99] , \block[2][98] ,
         \block[2][97] , \block[2][96] , \block[2][95] , \block[2][94] ,
         \block[2][93] , \block[2][92] , \block[2][91] , \block[2][90] ,
         \block[2][89] , \block[2][88] , \block[2][87] , \block[2][86] ,
         \block[2][85] , \block[2][84] , \block[2][83] , \block[2][82] ,
         \block[2][81] , \block[2][80] , \block[2][79] , \block[2][78] ,
         \block[2][77] , \block[2][76] , \block[2][75] , \block[2][74] ,
         \block[2][73] , \block[2][72] , \block[2][71] , \block[2][70] ,
         \block[2][69] , \block[2][68] , \block[2][67] , \block[2][66] ,
         \block[2][65] , \block[2][64] , \block[2][63] , \block[2][62] ,
         \block[2][61] , \block[2][60] , \block[2][59] , \block[2][58] ,
         \block[2][57] , \block[2][56] , \block[2][55] , \block[2][54] ,
         \block[2][53] , \block[2][52] , \block[2][51] , \block[2][50] ,
         \block[2][49] , \block[2][48] , \block[2][47] , \block[2][46] ,
         \block[2][45] , \block[2][44] , \block[2][43] , \block[2][42] ,
         \block[2][41] , \block[2][40] , \block[2][39] , \block[2][38] ,
         \block[2][37] , \block[2][36] , \block[2][35] , \block[2][34] ,
         \block[2][33] , \block[2][32] , \block[2][31] , \block[2][30] ,
         \block[2][29] , \block[2][28] , \block[2][27] , \block[2][26] ,
         \block[2][25] , \block[2][24] , \block[2][23] , \block[2][22] ,
         \block[2][21] , \block[2][20] , \block[2][19] , \block[2][18] ,
         \block[2][17] , \block[2][16] , \block[2][15] , \block[2][14] ,
         \block[2][13] , \block[2][12] , \block[2][11] , \block[2][10] ,
         \block[2][9] , \block[2][8] , \block[2][7] , \block[2][6] ,
         \block[2][5] , \block[2][4] , \block[2][3] , \block[2][2] ,
         \block[2][1] , \block[2][0] , \block[1][127] , \block[1][126] ,
         \block[1][125] , \block[1][124] , \block[1][123] , \block[1][122] ,
         \block[1][121] , \block[1][120] , \block[1][119] , \block[1][118] ,
         \block[1][117] , \block[1][116] , \block[1][115] , \block[1][114] ,
         \block[1][113] , \block[1][112] , \block[1][111] , \block[1][110] ,
         \block[1][109] , \block[1][108] , \block[1][107] , \block[1][106] ,
         \block[1][105] , \block[1][104] , \block[1][103] , \block[1][102] ,
         \block[1][101] , \block[1][100] , \block[1][99] , \block[1][98] ,
         \block[1][97] , \block[1][96] , \block[1][95] , \block[1][94] ,
         \block[1][93] , \block[1][92] , \block[1][91] , \block[1][90] ,
         \block[1][89] , \block[1][88] , \block[1][87] , \block[1][86] ,
         \block[1][85] , \block[1][84] , \block[1][83] , \block[1][82] ,
         \block[1][81] , \block[1][80] , \block[1][79] , \block[1][78] ,
         \block[1][77] , \block[1][76] , \block[1][75] , \block[1][74] ,
         \block[1][73] , \block[1][72] , \block[1][71] , \block[1][70] ,
         \block[1][69] , \block[1][68] , \block[1][67] , \block[1][66] ,
         \block[1][65] , \block[1][64] , \block[1][63] , \block[1][62] ,
         \block[1][61] , \block[1][60] , \block[1][59] , \block[1][58] ,
         \block[1][57] , \block[1][56] , \block[1][55] , \block[1][54] ,
         \block[1][53] , \block[1][52] , \block[1][51] , \block[1][50] ,
         \block[1][49] , \block[1][48] , \block[1][47] , \block[1][46] ,
         \block[1][45] , \block[1][44] , \block[1][43] , \block[1][42] ,
         \block[1][41] , \block[1][40] , \block[1][39] , \block[1][38] ,
         \block[1][37] , \block[1][36] , \block[1][35] , \block[1][34] ,
         \block[1][33] , \block[1][32] , \block[1][31] , \block[1][30] ,
         \block[1][29] , \block[1][28] , \block[1][27] , \block[1][26] ,
         \block[1][25] , \block[1][24] , \block[1][23] , \block[1][22] ,
         \block[1][21] , \block[1][20] , \block[1][19] , \block[1][18] ,
         \block[1][17] , \block[1][16] , \block[1][15] , \block[1][14] ,
         \block[1][13] , \block[1][12] , \block[1][11] , \block[1][10] ,
         \block[1][9] , \block[1][8] , \block[1][7] , \block[1][6] ,
         \block[1][5] , \block[1][4] , \block[1][3] , \block[1][2] ,
         \block[1][1] , \block[1][0] , \block[0][127] , \block[0][126] ,
         \block[0][125] , \block[0][124] , \block[0][123] , \block[0][122] ,
         \block[0][121] , \block[0][120] , \block[0][119] , \block[0][118] ,
         \block[0][117] , \block[0][116] , \block[0][115] , \block[0][114] ,
         \block[0][113] , \block[0][112] , \block[0][111] , \block[0][110] ,
         \block[0][109] , \block[0][108] , \block[0][107] , \block[0][106] ,
         \block[0][105] , \block[0][104] , \block[0][103] , \block[0][102] ,
         \block[0][101] , \block[0][100] , \block[0][99] , \block[0][98] ,
         \block[0][97] , \block[0][96] , \block[0][95] , \block[0][94] ,
         \block[0][93] , \block[0][92] , \block[0][91] , \block[0][90] ,
         \block[0][89] , \block[0][88] , \block[0][87] , \block[0][86] ,
         \block[0][85] , \block[0][84] , \block[0][83] , \block[0][82] ,
         \block[0][81] , \block[0][80] , \block[0][79] , \block[0][78] ,
         \block[0][77] , \block[0][76] , \block[0][75] , \block[0][74] ,
         \block[0][73] , \block[0][72] , \block[0][71] , \block[0][70] ,
         \block[0][69] , \block[0][68] , \block[0][67] , \block[0][66] ,
         \block[0][65] , \block[0][64] , \block[0][63] , \block[0][62] ,
         \block[0][61] , \block[0][60] , \block[0][59] , \block[0][58] ,
         \block[0][57] , \block[0][56] , \block[0][55] , \block[0][54] ,
         \block[0][53] , \block[0][52] , \block[0][51] , \block[0][50] ,
         \block[0][49] , \block[0][48] , \block[0][47] , \block[0][46] ,
         \block[0][45] , \block[0][44] , \block[0][43] , \block[0][42] ,
         \block[0][41] , \block[0][40] , \block[0][39] , \block[0][38] ,
         \block[0][37] , \block[0][36] , \block[0][35] , \block[0][34] ,
         \block[0][33] , \block[0][32] , \block[0][31] , \block[0][30] ,
         \block[0][29] , \block[0][28] , \block[0][27] , \block[0][26] ,
         \block[0][25] , \block[0][24] , \block[0][23] , \block[0][22] ,
         \block[0][21] , \block[0][20] , \block[0][19] , \block[0][18] ,
         \block[0][17] , \block[0][16] , \block[0][15] , \block[0][14] ,
         \block[0][13] , \block[0][12] , \block[0][11] , \block[0][10] ,
         \block[0][9] , \block[0][8] , \block[0][7] , \block[0][6] ,
         \block[0][5] , \block[0][4] , \block[0][3] , \block[0][2] ,
         \block[0][1] , \block[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n120, n122, n124, n126, n128, n130, n132, n134, n136, n138,
         n140, n142, n144, n146, n148, n150, n152, n154, n156, n158, n160,
         n162, n164, n166, n168, n170, n172, n174, n176, n178, n180, n182,
         n184, n186, n188, n190, n192, n194, n196, n198, n200, n202, n204,
         n206, n208, n210, n212, n214, n216, n218, n220, n222, n224, n226,
         n228, n230, n232, n234, n236, n238, n240, n242, n244, n246, n248,
         n250, n252, n254, n256, n258, n260, n262, n264, n266, n268, n270,
         n272, n274, n276, n278, n280, n282, n284, n286, n288, n290, n292,
         n294, n296, n298, n300, n302, n304, n306, n308, n310, n312, n314,
         n316, n318, n320, n322, n324, n326, n328, n330, n332, n334, n336,
         n338, n340, n342, n344, n346, n348, n350, n352, n354, n356, n358,
         n360, n362, n364, n366, n368, n370, n372, n374, n376, n378, n380,
         n382, n384, n386, n388, n390, n392, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n502, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n789, n790, n791, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  DFFRX4 \blockvalid_reg[7]  ( .D(n1712), .CK(clk), .RN(n794), .Q(
        blockvalid[7]), .QN(n1728) );
  DFFRX4 \blockvalid_reg[6]  ( .D(n1713), .CK(clk), .RN(n794), .Q(
        blockvalid[6]), .QN(n1729) );
  DFFRX4 \blockvalid_reg[4]  ( .D(n1715), .CK(clk), .RN(n794), .Q(
        blockvalid[4]), .QN(n1731) );
  DFFRX4 \blockvalid_reg[3]  ( .D(n1716), .CK(clk), .RN(n794), .Q(
        blockvalid[3]), .QN(n1732) );
  DFFRX4 \blockvalid_reg[2]  ( .D(n1717), .CK(clk), .RN(n794), .Q(
        blockvalid[2]), .QN(n1733) );
  EDFFXL \block_reg[2][113]  ( .D(block_next[113]), .E(n668), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFXL \block_reg[2][112]  ( .D(block_next[112]), .E(n668), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFXL \block_reg[2][90]  ( .D(block_next[90]), .E(n669), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFXL \block_reg[2][89]  ( .D(block_next[89]), .E(n669), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFXL \block_reg[2][88]  ( .D(block_next[88]), .E(n670), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFXL \block_reg[2][87]  ( .D(block_next[87]), .E(n670), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFXL \block_reg[2][84]  ( .D(block_next[84]), .E(n670), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFXL \block_reg[2][82]  ( .D(block_next[82]), .E(n670), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFXL \block_reg[2][81]  ( .D(block_next[81]), .E(n670), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFXL \block_reg[2][80]  ( .D(block_next[80]), .E(n670), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFX1 \block_reg[2][58]  ( .D(block_next[58]), .E(n672), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFX1 \block_reg[2][57]  ( .D(block_next[57]), .E(n672), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFX1 \block_reg[2][56]  ( .D(block_next[56]), .E(n672), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFX1 \block_reg[2][55]  ( .D(block_next[55]), .E(n672), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFX1 \block_reg[2][52]  ( .D(block_next[52]), .E(n672), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFX1 \block_reg[2][50]  ( .D(block_next[50]), .E(n672), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFX1 \block_reg[2][49]  ( .D(block_next[49]), .E(n673), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFX1 \block_reg[2][48]  ( .D(block_next[48]), .E(n673), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFX1 \block_reg[2][26]  ( .D(block_next[26]), .E(n674), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFX1 \block_reg[2][25]  ( .D(block_next[25]), .E(n674), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFX1 \block_reg[2][24]  ( .D(block_next[24]), .E(n674), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFX1 \block_reg[2][20]  ( .D(block_next[20]), .E(n675), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFXL \block_reg[2][122]  ( .D(block_next[122]), .E(n667), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFXL \block_reg[2][121]  ( .D(block_next[121]), .E(n667), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFXL \block_reg[2][120]  ( .D(block_next[120]), .E(n667), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFXL \block_reg[2][119]  ( .D(block_next[119]), .E(n667), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFXL \block_reg[2][118]  ( .D(block_next[118]), .E(n667), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFXL \block_reg[2][116]  ( .D(block_next[116]), .E(n667), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFXL \block_reg[2][114]  ( .D(block_next[114]), .E(n668), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFXL \block_reg[6][113]  ( .D(block_next[113]), .E(n603), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFXL \block_reg[6][112]  ( .D(block_next[112]), .E(n603), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFXL \block_reg[6][90]  ( .D(block_next[90]), .E(n604), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFXL \block_reg[6][89]  ( .D(block_next[89]), .E(n604), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFXL \block_reg[6][88]  ( .D(block_next[88]), .E(n605), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFXL \block_reg[6][87]  ( .D(block_next[87]), .E(n605), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFXL \block_reg[6][84]  ( .D(block_next[84]), .E(n605), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFXL \block_reg[6][82]  ( .D(block_next[82]), .E(n605), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFXL \block_reg[6][81]  ( .D(block_next[81]), .E(n605), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFXL \block_reg[6][80]  ( .D(block_next[80]), .E(n605), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFX1 \block_reg[6][58]  ( .D(block_next[58]), .E(n607), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFX1 \block_reg[6][57]  ( .D(block_next[57]), .E(n607), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFX1 \block_reg[6][56]  ( .D(block_next[56]), .E(n607), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFX1 \block_reg[6][55]  ( .D(block_next[55]), .E(n607), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n607), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[6][50]  ( .D(block_next[50]), .E(n607), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFX1 \block_reg[6][49]  ( .D(block_next[49]), .E(n608), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFX1 \block_reg[6][48]  ( .D(block_next[48]), .E(n608), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n610), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFXL \block_reg[6][122]  ( .D(block_next[122]), .E(n602), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFXL \block_reg[6][121]  ( .D(block_next[121]), .E(n602), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFXL \block_reg[6][120]  ( .D(block_next[120]), .E(n602), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFXL \block_reg[6][119]  ( .D(block_next[119]), .E(n602), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFXL \block_reg[6][118]  ( .D(block_next[118]), .E(n602), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFXL \block_reg[6][116]  ( .D(block_next[116]), .E(n602), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFXL \block_reg[6][114]  ( .D(block_next[114]), .E(n603), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFX1 \block_reg[2][54]  ( .D(block_next[54]), .E(n672), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFXL \block_reg[2][86]  ( .D(block_next[86]), .E(n670), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFX1 \block_reg[6][54]  ( .D(block_next[54]), .E(n607), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFXL \block_reg[6][86]  ( .D(block_next[86]), .E(n605), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFXL \block_reg[2][117]  ( .D(block_next[117]), .E(n667), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFX1 \block_reg[2][51]  ( .D(block_next[51]), .E(n672), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFX1 \block_reg[2][53]  ( .D(block_next[53]), .E(n672), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFXL \block_reg[6][117]  ( .D(block_next[117]), .E(n602), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFXL \block_reg[2][115]  ( .D(block_next[115]), .E(n667), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFX1 \block_reg[6][51]  ( .D(block_next[51]), .E(n607), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n607), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFXL \block_reg[6][115]  ( .D(block_next[115]), .E(n602), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFXL \block_reg[2][85]  ( .D(block_next[85]), .E(n670), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFXL \block_reg[6][85]  ( .D(block_next[85]), .E(n605), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFXL \block_reg[2][83]  ( .D(block_next[83]), .E(n670), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFXL \block_reg[6][83]  ( .D(block_next[83]), .E(n605), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFXL \block_reg[2][109]  ( .D(block_next[109]), .E(n668), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFXL \block_reg[6][109]  ( .D(block_next[109]), .E(n603), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFXL \block_reg[6][108]  ( .D(block_next[108]), .E(n603), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFXL \block_reg[2][108]  ( .D(block_next[108]), .E(n668), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFX1 \block_reg[6][45]  ( .D(block_next[45]), .E(n608), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFXL \block_reg[6][76]  ( .D(block_next[76]), .E(n605), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFX1 \block_reg[2][45]  ( .D(block_next[45]), .E(n673), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFXL \block_reg[2][76]  ( .D(block_next[76]), .E(n670), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFXL \block_reg[6][68]  ( .D(block_next[68]), .E(n606), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFXL \block_reg[2][110]  ( .D(block_next[110]), .E(n668), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFXL \block_reg[2][68]  ( .D(block_next[68]), .E(n671), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFXL \block_reg[6][110]  ( .D(block_next[110]), .E(n603), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFXL \block_reg[2][77]  ( .D(block_next[77]), .E(n670), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFXL \block_reg[6][77]  ( .D(block_next[77]), .E(n605), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFXL \block_reg[6][104]  ( .D(block_next[104]), .E(n603), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFXL \block_reg[2][104]  ( .D(block_next[104]), .E(n668), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFX1 \block_reg[6][44]  ( .D(block_next[44]), .E(n608), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFX1 \block_reg[2][44]  ( .D(block_next[44]), .E(n673), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFXL \block_reg[2][106]  ( .D(block_next[106]), .E(n668), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFXL \block_reg[6][106]  ( .D(block_next[106]), .E(n603), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFXL \block_reg[6][100]  ( .D(block_next[100]), .E(n604), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFXL \block_reg[2][100]  ( .D(block_next[100]), .E(n669), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFXL \block_reg[6][73]  ( .D(block_next[73]), .E(n606), .CK(clk), .Q(
        \block[6][73] ) );
  EDFFXL \block_reg[2][73]  ( .D(block_next[73]), .E(n671), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFXL \block_reg[2][74]  ( .D(block_next[74]), .E(n671), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFXL \block_reg[6][102]  ( .D(block_next[102]), .E(n603), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFXL \block_reg[6][72]  ( .D(block_next[72]), .E(n606), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFX1 \block_reg[6][6]  ( .D(block_next[6]), .E(n611), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFXL \block_reg[2][102]  ( .D(block_next[102]), .E(n668), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFXL \block_reg[6][105]  ( .D(block_next[105]), .E(n603), .CK(clk), .Q(
        \block[6][105] ) );
  EDFFXL \block_reg[2][72]  ( .D(block_next[72]), .E(n671), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFXL \block_reg[2][105]  ( .D(block_next[105]), .E(n668), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFX1 \block_reg[2][6]  ( .D(block_next[6]), .E(n676), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFXL \block_reg[2][78]  ( .D(block_next[78]), .E(n670), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFXL \block_reg[6][74]  ( .D(block_next[74]), .E(n606), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFXL \block_reg[2][79]  ( .D(block_next[79]), .E(n670), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n609), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFXL \block_reg[6][78]  ( .D(block_next[78]), .E(n605), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFX1 \block_reg[2][36]  ( .D(block_next[36]), .E(n674), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFXL \block_reg[6][70]  ( .D(block_next[70]), .E(n606), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFXL \block_reg[6][79]  ( .D(block_next[79]), .E(n605), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFXL \block_reg[2][70]  ( .D(block_next[70]), .E(n671), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFX1 \block_reg[2][46]  ( .D(block_next[46]), .E(n673), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFX1 \block_reg[6][40]  ( .D(block_next[40]), .E(n608), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFX1 \block_reg[6][46]  ( .D(block_next[46]), .E(n608), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFX1 \block_reg[2][40]  ( .D(block_next[40]), .E(n673), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFXL \block_reg[2][111]  ( .D(block_next[111]), .E(n668), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFXL \block_reg[6][111]  ( .D(block_next[111]), .E(n603), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFX1 \block_reg[2][42]  ( .D(block_next[42]), .E(n673), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFX1 \block_reg[6][42]  ( .D(block_next[42]), .E(n608), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n608), .CK(clk), .Q(
        \block[6][41] ) );
  EDFFX1 \block_reg[2][41]  ( .D(block_next[41]), .E(n673), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n608), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[2][38]  ( .D(block_next[38]), .E(n673), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFXL \block_reg[6][107]  ( .D(block_next[107]), .E(n603), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFXL \block_reg[2][107]  ( .D(block_next[107]), .E(n668), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFX1 \block_reg[2][47]  ( .D(block_next[47]), .E(n673), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFX1 \block_reg[6][47]  ( .D(block_next[47]), .E(n608), .CK(clk), .Q(
        \block[6][47] ) );
  EDFFXL \block_reg[6][98]  ( .D(block_next[98]), .E(n604), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFXL \block_reg[2][98]  ( .D(block_next[98]), .E(n669), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFXL \block_reg[6][97]  ( .D(block_next[97]), .E(n604), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFXL \block_reg[2][97]  ( .D(block_next[97]), .E(n669), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFXL \block_reg[2][75]  ( .D(block_next[75]), .E(n671), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFX1 \block_reg[6][33]  ( .D(block_next[33]), .E(n609), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFX1 \block_reg[2][33]  ( .D(block_next[33]), .E(n674), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFXL \block_reg[6][75]  ( .D(block_next[75]), .E(n606), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFXL \block_reg[2][66]  ( .D(block_next[66]), .E(n671), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFXL \block_reg[6][66]  ( .D(block_next[66]), .E(n606), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFX1 \block_reg[6][43]  ( .D(block_next[43]), .E(n608), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFXL \block_reg[2][65]  ( .D(block_next[65]), .E(n671), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFX1 \block_reg[2][43]  ( .D(block_next[43]), .E(n673), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFXL \block_reg[6][65]  ( .D(block_next[65]), .E(n606), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFX1 \block_reg[2][34]  ( .D(block_next[34]), .E(n674), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFX1 \block_reg[6][34]  ( .D(block_next[34]), .E(n609), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFXL \block_reg[6][103]  ( .D(block_next[103]), .E(n603), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFXL \block_reg[2][103]  ( .D(block_next[103]), .E(n668), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFXL \block_reg[2][67]  ( .D(block_next[67]), .E(n671), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFX1 \block_reg[6][39]  ( .D(block_next[39]), .E(n608), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFX1 \block_reg[2][39]  ( .D(block_next[39]), .E(n673), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFXL \block_reg[6][67]  ( .D(block_next[67]), .E(n606), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFXL \block_reg[6][99]  ( .D(block_next[99]), .E(n604), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFXL \block_reg[2][99]  ( .D(block_next[99]), .E(n669), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFXL \block_reg[6][71]  ( .D(block_next[71]), .E(n606), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFXL \block_reg[2][71]  ( .D(block_next[71]), .E(n671), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFXL \block_reg[6][101]  ( .D(block_next[101]), .E(n604), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFXL \block_reg[2][101]  ( .D(block_next[101]), .E(n669), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFXL \block_reg[6][69]  ( .D(block_next[69]), .E(n606), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFXL \block_reg[2][69]  ( .D(block_next[69]), .E(n671), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n608), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[2][37]  ( .D(block_next[37]), .E(n673), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFX1 \block_reg[2][35]  ( .D(block_next[35]), .E(n674), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n609), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFXL \block_reg[6][96]  ( .D(block_next[96]), .E(n604), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFXL \block_reg[2][96]  ( .D(block_next[96]), .E(n669), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFXL \block_reg[6][64]  ( .D(block_next[64]), .E(n606), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFXL \block_reg[2][64]  ( .D(block_next[64]), .E(n671), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n609), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[2][32]  ( .D(block_next[32]), .E(n674), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFX1 \block_reg[6][27]  ( .D(block_next[27]), .E(n609), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFX1 \block_reg[2][27]  ( .D(block_next[27]), .E(n674), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFXL \block_reg[6][127]  ( .D(block_next[127]), .E(n602), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFXL \block_reg[2][127]  ( .D(block_next[127]), .E(n667), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFXL \block_reg[6][124]  ( .D(block_next[124]), .E(n602), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFXL \block_reg[2][124]  ( .D(block_next[124]), .E(n667), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFXL \block_reg[6][125]  ( .D(block_next[125]), .E(n602), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFXL \block_reg[2][125]  ( .D(block_next[125]), .E(n667), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFXL \block_reg[6][126]  ( .D(block_next[126]), .E(n602), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFXL \block_reg[2][126]  ( .D(block_next[126]), .E(n667), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFXL \block_reg[6][123]  ( .D(block_next[123]), .E(n602), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFXL \block_reg[2][123]  ( .D(block_next[123]), .E(n667), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFX1 \block_reg[2][28]  ( .D(block_next[28]), .E(n674), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFX1 \block_reg[6][28]  ( .D(block_next[28]), .E(n609), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFX1 \block_reg[6][30]  ( .D(block_next[30]), .E(n609), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFX1 \block_reg[2][30]  ( .D(block_next[30]), .E(n674), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFX1 \block_reg[2][29]  ( .D(block_next[29]), .E(n674), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFX1 \block_reg[6][29]  ( .D(block_next[29]), .E(n609), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFX1 \block_reg[6][31]  ( .D(block_next[31]), .E(n609), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFX1 \block_reg[2][31]  ( .D(block_next[31]), .E(n674), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFXL \block_reg[3][113]  ( .D(block_next[113]), .E(n652), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFXL \block_reg[3][112]  ( .D(block_next[112]), .E(n652), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFXL \block_reg[3][90]  ( .D(block_next[90]), .E(n653), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFXL \block_reg[3][89]  ( .D(block_next[89]), .E(n653), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFXL \block_reg[3][88]  ( .D(block_next[88]), .E(n654), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFXL \block_reg[3][87]  ( .D(block_next[87]), .E(n654), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFXL \block_reg[3][84]  ( .D(block_next[84]), .E(n654), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFXL \block_reg[3][82]  ( .D(block_next[82]), .E(n654), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFXL \block_reg[3][81]  ( .D(block_next[81]), .E(n654), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFXL \block_reg[3][80]  ( .D(block_next[80]), .E(n654), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFX1 \block_reg[3][58]  ( .D(block_next[58]), .E(n656), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFX1 \block_reg[3][57]  ( .D(block_next[57]), .E(n656), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFX1 \block_reg[3][56]  ( .D(block_next[56]), .E(n656), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFX1 \block_reg[3][55]  ( .D(block_next[55]), .E(n656), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n656), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[3][50]  ( .D(block_next[50]), .E(n656), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n657), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[3][48]  ( .D(block_next[48]), .E(n657), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFX1 \block_reg[3][26]  ( .D(block_next[26]), .E(n658), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFX1 \block_reg[3][25]  ( .D(block_next[25]), .E(n658), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFX1 \block_reg[3][24]  ( .D(block_next[24]), .E(n658), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n659), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFXL \block_reg[3][122]  ( .D(block_next[122]), .E(n651), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFXL \block_reg[3][121]  ( .D(block_next[121]), .E(n651), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFXL \block_reg[3][120]  ( .D(block_next[120]), .E(n651), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFXL \block_reg[3][119]  ( .D(block_next[119]), .E(n651), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFXL \block_reg[3][118]  ( .D(block_next[118]), .E(n651), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFXL \block_reg[3][116]  ( .D(block_next[116]), .E(n651), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFXL \block_reg[3][114]  ( .D(block_next[114]), .E(n652), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFXL \block_reg[7][113]  ( .D(block_next[113]), .E(n588), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFXL \block_reg[7][112]  ( .D(block_next[112]), .E(n588), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFXL \block_reg[7][90]  ( .D(block_next[90]), .E(n589), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFXL \block_reg[7][89]  ( .D(block_next[89]), .E(n589), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFXL \block_reg[7][88]  ( .D(block_next[88]), .E(n590), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFXL \block_reg[7][87]  ( .D(block_next[87]), .E(n590), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFXL \block_reg[7][84]  ( .D(block_next[84]), .E(n590), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFXL \block_reg[7][82]  ( .D(block_next[82]), .E(n590), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFXL \block_reg[7][81]  ( .D(block_next[81]), .E(n590), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFXL \block_reg[7][80]  ( .D(block_next[80]), .E(n590), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFX1 \block_reg[7][58]  ( .D(block_next[58]), .E(n592), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFX1 \block_reg[7][57]  ( .D(block_next[57]), .E(n592), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFX1 \block_reg[7][56]  ( .D(block_next[56]), .E(n592), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFX1 \block_reg[7][55]  ( .D(block_next[55]), .E(n592), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n592), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[7][50]  ( .D(block_next[50]), .E(n592), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n593), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[7][48]  ( .D(block_next[48]), .E(n593), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFXL \block_reg[7][122]  ( .D(block_next[122]), .E(n587), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFXL \block_reg[7][121]  ( .D(block_next[121]), .E(n587), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFXL \block_reg[7][120]  ( .D(block_next[120]), .E(n587), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFXL \block_reg[7][119]  ( .D(block_next[119]), .E(n587), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFXL \block_reg[7][118]  ( .D(block_next[118]), .E(n587), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFXL \block_reg[7][116]  ( .D(block_next[116]), .E(n587), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFXL \block_reg[7][114]  ( .D(block_next[114]), .E(n588), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFX1 \block_reg[3][54]  ( .D(block_next[54]), .E(n656), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFXL \block_reg[3][86]  ( .D(block_next[86]), .E(n654), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFX1 \block_reg[7][54]  ( .D(block_next[54]), .E(n592), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFXL \block_reg[7][86]  ( .D(block_next[86]), .E(n590), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFXL \block_reg[3][117]  ( .D(block_next[117]), .E(n651), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFX1 \block_reg[3][51]  ( .D(block_next[51]), .E(n656), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n656), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFXL \block_reg[7][117]  ( .D(block_next[117]), .E(n587), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFXL \block_reg[3][115]  ( .D(block_next[115]), .E(n651), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFX1 \block_reg[7][51]  ( .D(block_next[51]), .E(n592), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n592), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFXL \block_reg[7][115]  ( .D(block_next[115]), .E(n587), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFXL \block_reg[3][85]  ( .D(block_next[85]), .E(n654), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFXL \block_reg[7][85]  ( .D(block_next[85]), .E(n590), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFXL \block_reg[3][83]  ( .D(block_next[83]), .E(n654), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFXL \block_reg[7][83]  ( .D(block_next[83]), .E(n590), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFXL \block_reg[3][109]  ( .D(block_next[109]), .E(n652), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFXL \block_reg[7][108]  ( .D(block_next[108]), .E(n588), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFXL \block_reg[3][108]  ( .D(block_next[108]), .E(n652), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFXL \block_reg[7][109]  ( .D(block_next[109]), .E(n588), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFX1 \block_reg[7][45]  ( .D(block_next[45]), .E(n593), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFXL \block_reg[7][76]  ( .D(block_next[76]), .E(n590), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFX1 \block_reg[3][45]  ( .D(block_next[45]), .E(n657), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFXL \block_reg[3][76]  ( .D(block_next[76]), .E(n654), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFXL \block_reg[7][68]  ( .D(block_next[68]), .E(n591), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFXL \block_reg[3][68]  ( .D(block_next[68]), .E(n655), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFXL \block_reg[3][110]  ( .D(block_next[110]), .E(n652), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFXL \block_reg[7][110]  ( .D(block_next[110]), .E(n588), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFXL \block_reg[3][77]  ( .D(block_next[77]), .E(n654), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFXL \block_reg[7][104]  ( .D(block_next[104]), .E(n588), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFXL \block_reg[3][104]  ( .D(block_next[104]), .E(n652), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFX1 \block_reg[7][44]  ( .D(block_next[44]), .E(n593), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFXL \block_reg[7][77]  ( .D(block_next[77]), .E(n590), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFX1 \block_reg[3][44]  ( .D(block_next[44]), .E(n657), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFXL \block_reg[7][100]  ( .D(block_next[100]), .E(n589), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFXL \block_reg[3][100]  ( .D(block_next[100]), .E(n653), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFXL \block_reg[3][106]  ( .D(block_next[106]), .E(n652), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFXL \block_reg[7][106]  ( .D(block_next[106]), .E(n588), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFXL \block_reg[7][73]  ( .D(block_next[73]), .E(n591), .CK(clk), .Q(
        \block[7][73] ) );
  EDFFXL \block_reg[3][73]  ( .D(block_next[73]), .E(n655), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFXL \block_reg[7][102]  ( .D(block_next[102]), .E(n588), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFXL \block_reg[7][72]  ( .D(block_next[72]), .E(n591), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFXL \block_reg[3][102]  ( .D(block_next[102]), .E(n652), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFXL \block_reg[7][105]  ( .D(block_next[105]), .E(n588), .CK(clk), .Q(
        \block[7][105] ) );
  EDFFXL \block_reg[3][72]  ( .D(block_next[72]), .E(n655), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFXL \block_reg[3][105]  ( .D(block_next[105]), .E(n652), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFX1 \block_reg[3][6]  ( .D(block_next[6]), .E(n660), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFXL \block_reg[3][74]  ( .D(block_next[74]), .E(n655), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n594), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n658), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFXL \block_reg[7][74]  ( .D(block_next[74]), .E(n591), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFXL \block_reg[3][78]  ( .D(block_next[78]), .E(n654), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFXL \block_reg[7][70]  ( .D(block_next[70]), .E(n591), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFXL \block_reg[3][70]  ( .D(block_next[70]), .E(n655), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFXL \block_reg[7][78]  ( .D(block_next[78]), .E(n590), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFXL \block_reg[3][79]  ( .D(block_next[79]), .E(n654), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFX1 \block_reg[7][40]  ( .D(block_next[40]), .E(n593), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFX1 \block_reg[3][40]  ( .D(block_next[40]), .E(n657), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFX1 \block_reg[3][46]  ( .D(block_next[46]), .E(n657), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFXL \block_reg[7][79]  ( .D(block_next[79]), .E(n590), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFX1 \block_reg[7][46]  ( .D(block_next[46]), .E(n593), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFXL \block_reg[3][111]  ( .D(block_next[111]), .E(n652), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n593), .CK(clk), .Q(
        \block[7][41] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n657), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[3][42]  ( .D(block_next[42]), .E(n657), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n593), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n657), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFXL \block_reg[7][107]  ( .D(block_next[107]), .E(n588), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFXL \block_reg[7][111]  ( .D(block_next[111]), .E(n588), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFXL \block_reg[3][107]  ( .D(block_next[107]), .E(n652), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFX1 \block_reg[7][42]  ( .D(block_next[42]), .E(n593), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFX1 \block_reg[3][47]  ( .D(block_next[47]), .E(n657), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFXL \block_reg[7][98]  ( .D(block_next[98]), .E(n589), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFXL \block_reg[3][98]  ( .D(block_next[98]), .E(n653), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFX1 \block_reg[7][47]  ( .D(block_next[47]), .E(n593), .CK(clk), .Q(
        \block[7][47] ) );
  EDFFXL \block_reg[7][97]  ( .D(block_next[97]), .E(n589), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFXL \block_reg[3][97]  ( .D(block_next[97]), .E(n653), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFX1 \block_reg[7][33]  ( .D(block_next[33]), .E(n594), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFX1 \block_reg[3][33]  ( .D(block_next[33]), .E(n658), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFXL \block_reg[3][75]  ( .D(block_next[75]), .E(n655), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFXL \block_reg[7][75]  ( .D(block_next[75]), .E(n591), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFXL \block_reg[3][66]  ( .D(block_next[66]), .E(n655), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFX1 \block_reg[7][43]  ( .D(block_next[43]), .E(n593), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFX1 \block_reg[3][43]  ( .D(block_next[43]), .E(n657), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFXL \block_reg[7][66]  ( .D(block_next[66]), .E(n591), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFXL \block_reg[3][65]  ( .D(block_next[65]), .E(n655), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFXL \block_reg[7][65]  ( .D(block_next[65]), .E(n591), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n658), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n594), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFXL \block_reg[7][103]  ( .D(block_next[103]), .E(n588), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFXL \block_reg[3][103]  ( .D(block_next[103]), .E(n652), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFX1 \block_reg[7][39]  ( .D(block_next[39]), .E(n593), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFX1 \block_reg[3][39]  ( .D(block_next[39]), .E(n657), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFXL \block_reg[3][67]  ( .D(block_next[67]), .E(n655), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFXL \block_reg[7][67]  ( .D(block_next[67]), .E(n591), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFXL \block_reg[7][99]  ( .D(block_next[99]), .E(n589), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFXL \block_reg[3][99]  ( .D(block_next[99]), .E(n653), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFXL \block_reg[7][71]  ( .D(block_next[71]), .E(n591), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFXL \block_reg[3][71]  ( .D(block_next[71]), .E(n655), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFXL \block_reg[7][101]  ( .D(block_next[101]), .E(n589), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFXL \block_reg[3][101]  ( .D(block_next[101]), .E(n653), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFXL \block_reg[7][69]  ( .D(block_next[69]), .E(n591), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFXL \block_reg[3][69]  ( .D(block_next[69]), .E(n655), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n593), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n657), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n658), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n594), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFXL \block_reg[7][96]  ( .D(block_next[96]), .E(n589), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFXL \block_reg[3][96]  ( .D(block_next[96]), .E(n653), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFXL \block_reg[7][64]  ( .D(block_next[64]), .E(n591), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFXL \block_reg[3][64]  ( .D(block_next[64]), .E(n655), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n594), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n658), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[7][27]  ( .D(block_next[27]), .E(n594), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFX1 \block_reg[3][27]  ( .D(block_next[27]), .E(n658), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFXL \block_reg[7][127]  ( .D(block_next[127]), .E(n587), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFXL \block_reg[3][127]  ( .D(block_next[127]), .E(n651), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFXL \block_reg[7][124]  ( .D(block_next[124]), .E(n587), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFXL \block_reg[3][124]  ( .D(block_next[124]), .E(n651), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFXL \block_reg[7][125]  ( .D(block_next[125]), .E(n587), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFXL \block_reg[3][125]  ( .D(block_next[125]), .E(n651), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFXL \block_reg[7][126]  ( .D(block_next[126]), .E(n587), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFXL \block_reg[3][126]  ( .D(block_next[126]), .E(n651), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFXL \block_reg[7][123]  ( .D(block_next[123]), .E(n587), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFXL \block_reg[3][123]  ( .D(block_next[123]), .E(n651), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFX1 \block_reg[3][28]  ( .D(block_next[28]), .E(n658), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFX1 \block_reg[7][30]  ( .D(block_next[30]), .E(n594), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFX1 \block_reg[3][30]  ( .D(block_next[30]), .E(n658), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFX1 \block_reg[7][28]  ( .D(block_next[28]), .E(n594), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFX1 \block_reg[3][29]  ( .D(block_next[29]), .E(n658), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFX1 \block_reg[7][29]  ( .D(block_next[29]), .E(n594), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFX1 \block_reg[7][31]  ( .D(block_next[31]), .E(n594), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFX1 \block_reg[3][31]  ( .D(block_next[31]), .E(n658), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFXL \block_reg[0][113]  ( .D(block_next[113]), .E(n698), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFXL \block_reg[0][112]  ( .D(block_next[112]), .E(n698), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFXL \block_reg[0][90]  ( .D(block_next[90]), .E(n699), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFXL \block_reg[0][89]  ( .D(block_next[89]), .E(n699), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFXL \block_reg[0][88]  ( .D(block_next[88]), .E(n700), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFXL \block_reg[0][87]  ( .D(block_next[87]), .E(n700), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFXL \block_reg[0][84]  ( .D(block_next[84]), .E(n700), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFXL \block_reg[0][82]  ( .D(block_next[82]), .E(n700), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFXL \block_reg[0][81]  ( .D(block_next[81]), .E(n700), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFXL \block_reg[0][80]  ( .D(block_next[80]), .E(n700), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFX1 \block_reg[0][58]  ( .D(block_next[58]), .E(n702), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFX1 \block_reg[0][57]  ( .D(block_next[57]), .E(n702), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFX1 \block_reg[0][56]  ( .D(block_next[56]), .E(n702), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFX1 \block_reg[0][55]  ( .D(block_next[55]), .E(n702), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n702), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[0][50]  ( .D(block_next[50]), .E(n702), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n703), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[0][48]  ( .D(block_next[48]), .E(n703), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFX1 \block_reg[0][26]  ( .D(block_next[26]), .E(n704), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFX1 \block_reg[0][25]  ( .D(block_next[25]), .E(n704), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFX1 \block_reg[0][24]  ( .D(block_next[24]), .E(n704), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n705), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFXL \block_reg[0][122]  ( .D(block_next[122]), .E(n697), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFXL \block_reg[0][121]  ( .D(block_next[121]), .E(n697), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFXL \block_reg[0][120]  ( .D(block_next[120]), .E(n697), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFXL \block_reg[0][119]  ( .D(block_next[119]), .E(n697), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFXL \block_reg[0][118]  ( .D(block_next[118]), .E(n697), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFXL \block_reg[0][116]  ( .D(block_next[116]), .E(n697), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFXL \block_reg[0][114]  ( .D(block_next[114]), .E(n698), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFXL \block_reg[4][113]  ( .D(block_next[113]), .E(n634), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFXL \block_reg[4][112]  ( .D(block_next[112]), .E(n634), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFXL \block_reg[4][90]  ( .D(block_next[90]), .E(n635), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFXL \block_reg[4][89]  ( .D(block_next[89]), .E(n635), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFXL \block_reg[4][88]  ( .D(block_next[88]), .E(n636), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFXL \block_reg[4][87]  ( .D(block_next[87]), .E(n636), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFXL \block_reg[4][84]  ( .D(block_next[84]), .E(n636), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFXL \block_reg[4][82]  ( .D(block_next[82]), .E(n636), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFXL \block_reg[4][81]  ( .D(block_next[81]), .E(n636), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFXL \block_reg[4][80]  ( .D(block_next[80]), .E(n636), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFX1 \block_reg[4][58]  ( .D(block_next[58]), .E(n638), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFX1 \block_reg[4][57]  ( .D(block_next[57]), .E(n638), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFX1 \block_reg[4][56]  ( .D(block_next[56]), .E(n638), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFX1 \block_reg[4][55]  ( .D(block_next[55]), .E(n638), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n638), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[4][50]  ( .D(block_next[50]), .E(n638), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n639), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[4][48]  ( .D(block_next[48]), .E(n639), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFX1 \block_reg[4][26]  ( .D(block_next[26]), .E(n640), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFX1 \block_reg[4][25]  ( .D(block_next[25]), .E(n640), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFX1 \block_reg[4][24]  ( .D(block_next[24]), .E(n640), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n641), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFXL \block_reg[4][122]  ( .D(block_next[122]), .E(n633), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFXL \block_reg[4][121]  ( .D(block_next[121]), .E(n633), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFXL \block_reg[4][120]  ( .D(block_next[120]), .E(n633), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFXL \block_reg[4][119]  ( .D(block_next[119]), .E(n633), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFXL \block_reg[4][118]  ( .D(block_next[118]), .E(n633), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFXL \block_reg[4][116]  ( .D(block_next[116]), .E(n633), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFXL \block_reg[4][114]  ( .D(block_next[114]), .E(n634), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFX1 \block_reg[0][54]  ( .D(block_next[54]), .E(n702), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFXL \block_reg[0][86]  ( .D(block_next[86]), .E(n700), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFX1 \block_reg[4][54]  ( .D(block_next[54]), .E(n638), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFXL \block_reg[4][86]  ( .D(block_next[86]), .E(n636), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFXL \block_reg[0][117]  ( .D(block_next[117]), .E(n697), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFX1 \block_reg[0][51]  ( .D(block_next[51]), .E(n702), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n702), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFXL \block_reg[4][117]  ( .D(block_next[117]), .E(n633), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFXL \block_reg[0][115]  ( .D(block_next[115]), .E(n697), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFX1 \block_reg[4][51]  ( .D(block_next[51]), .E(n638), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n638), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFXL \block_reg[4][115]  ( .D(block_next[115]), .E(n633), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFXL \block_reg[0][85]  ( .D(block_next[85]), .E(n700), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFXL \block_reg[4][85]  ( .D(block_next[85]), .E(n636), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFXL \block_reg[0][83]  ( .D(block_next[83]), .E(n700), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFXL \block_reg[4][83]  ( .D(block_next[83]), .E(n636), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFXL \block_reg[0][109]  ( .D(block_next[109]), .E(n698), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFXL \block_reg[4][109]  ( .D(block_next[109]), .E(n634), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFXL \block_reg[4][108]  ( .D(block_next[108]), .E(n634), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFXL \block_reg[0][108]  ( .D(block_next[108]), .E(n698), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFX1 \block_reg[4][45]  ( .D(block_next[45]), .E(n639), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFXL \block_reg[4][76]  ( .D(block_next[76]), .E(n636), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFX1 \block_reg[0][45]  ( .D(block_next[45]), .E(n703), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFXL \block_reg[0][76]  ( .D(block_next[76]), .E(n700), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFXL \block_reg[0][110]  ( .D(block_next[110]), .E(n698), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFXL \block_reg[4][68]  ( .D(block_next[68]), .E(n637), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFXL \block_reg[0][68]  ( .D(block_next[68]), .E(n701), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFXL \block_reg[4][110]  ( .D(block_next[110]), .E(n634), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFXL \block_reg[0][77]  ( .D(block_next[77]), .E(n700), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFXL \block_reg[4][77]  ( .D(block_next[77]), .E(n636), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFXL \block_reg[4][104]  ( .D(block_next[104]), .E(n634), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFXL \block_reg[0][104]  ( .D(block_next[104]), .E(n698), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFX1 \block_reg[4][44]  ( .D(block_next[44]), .E(n639), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFX1 \block_reg[0][44]  ( .D(block_next[44]), .E(n703), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFXL \block_reg[0][106]  ( .D(block_next[106]), .E(n698), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFXL \block_reg[4][106]  ( .D(block_next[106]), .E(n634), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFXL \block_reg[4][100]  ( .D(block_next[100]), .E(n635), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFXL \block_reg[0][100]  ( .D(block_next[100]), .E(n699), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFXL \block_reg[4][73]  ( .D(block_next[73]), .E(n637), .CK(clk), .Q(
        \block[4][73] ) );
  EDFFXL \block_reg[0][73]  ( .D(block_next[73]), .E(n701), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFXL \block_reg[0][74]  ( .D(block_next[74]), .E(n701), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFXL \block_reg[4][102]  ( .D(block_next[102]), .E(n634), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFXL \block_reg[4][72]  ( .D(block_next[72]), .E(n637), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFXL \block_reg[0][78]  ( .D(block_next[78]), .E(n700), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFXL \block_reg[0][102]  ( .D(block_next[102]), .E(n698), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFX1 \block_reg[4][6]  ( .D(block_next[6]), .E(n642), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFXL \block_reg[4][105]  ( .D(block_next[105]), .E(n634), .CK(clk), .Q(
        \block[4][105] ) );
  EDFFXL \block_reg[0][72]  ( .D(block_next[72]), .E(n701), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFXL \block_reg[4][74]  ( .D(block_next[74]), .E(n637), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFXL \block_reg[0][105]  ( .D(block_next[105]), .E(n698), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFX1 \block_reg[0][6]  ( .D(block_next[6]), .E(n706), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFXL \block_reg[0][79]  ( .D(block_next[79]), .E(n700), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFXL \block_reg[4][78]  ( .D(block_next[78]), .E(n636), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n640), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n704), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFXL \block_reg[4][79]  ( .D(block_next[79]), .E(n636), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFX1 \block_reg[0][46]  ( .D(block_next[46]), .E(n703), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFXL \block_reg[4][70]  ( .D(block_next[70]), .E(n637), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFXL \block_reg[0][70]  ( .D(block_next[70]), .E(n701), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFX1 \block_reg[4][46]  ( .D(block_next[46]), .E(n639), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFX1 \block_reg[4][40]  ( .D(block_next[40]), .E(n639), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFX1 \block_reg[0][40]  ( .D(block_next[40]), .E(n703), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFXL \block_reg[0][111]  ( .D(block_next[111]), .E(n698), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFXL \block_reg[4][111]  ( .D(block_next[111]), .E(n634), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFX1 \block_reg[0][42]  ( .D(block_next[42]), .E(n703), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFX1 \block_reg[4][42]  ( .D(block_next[42]), .E(n639), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n639), .CK(clk), .Q(
        \block[4][41] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n703), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n639), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n703), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFXL \block_reg[4][107]  ( .D(block_next[107]), .E(n634), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFXL \block_reg[0][107]  ( .D(block_next[107]), .E(n698), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFX1 \block_reg[0][47]  ( .D(block_next[47]), .E(n703), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFX1 \block_reg[4][47]  ( .D(block_next[47]), .E(n639), .CK(clk), .Q(
        \block[4][47] ) );
  EDFFXL \block_reg[4][98]  ( .D(block_next[98]), .E(n635), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFXL \block_reg[0][98]  ( .D(block_next[98]), .E(n699), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFXL \block_reg[4][97]  ( .D(block_next[97]), .E(n635), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFXL \block_reg[0][97]  ( .D(block_next[97]), .E(n699), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFXL \block_reg[0][75]  ( .D(block_next[75]), .E(n701), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFXL \block_reg[4][75]  ( .D(block_next[75]), .E(n637), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFX1 \block_reg[4][33]  ( .D(block_next[33]), .E(n640), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFX1 \block_reg[0][33]  ( .D(block_next[33]), .E(n704), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFXL \block_reg[0][66]  ( .D(block_next[66]), .E(n701), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFXL \block_reg[4][66]  ( .D(block_next[66]), .E(n637), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFXL \block_reg[0][65]  ( .D(block_next[65]), .E(n701), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFX1 \block_reg[4][43]  ( .D(block_next[43]), .E(n639), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFX1 \block_reg[0][43]  ( .D(block_next[43]), .E(n703), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFXL \block_reg[4][65]  ( .D(block_next[65]), .E(n637), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFX1 \block_reg[0][34]  ( .D(block_next[34]), .E(n704), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFX1 \block_reg[4][34]  ( .D(block_next[34]), .E(n640), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFXL \block_reg[4][103]  ( .D(block_next[103]), .E(n634), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFXL \block_reg[0][103]  ( .D(block_next[103]), .E(n698), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFXL \block_reg[0][67]  ( .D(block_next[67]), .E(n701), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFX1 \block_reg[4][39]  ( .D(block_next[39]), .E(n639), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFXL \block_reg[4][67]  ( .D(block_next[67]), .E(n637), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFX1 \block_reg[0][39]  ( .D(block_next[39]), .E(n703), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFXL \block_reg[4][99]  ( .D(block_next[99]), .E(n635), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFXL \block_reg[0][99]  ( .D(block_next[99]), .E(n699), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFXL \block_reg[4][71]  ( .D(block_next[71]), .E(n637), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFXL \block_reg[0][71]  ( .D(block_next[71]), .E(n701), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFXL \block_reg[4][101]  ( .D(block_next[101]), .E(n635), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFXL \block_reg[0][101]  ( .D(block_next[101]), .E(n699), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFXL \block_reg[4][69]  ( .D(block_next[69]), .E(n637), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFXL \block_reg[0][69]  ( .D(block_next[69]), .E(n701), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n639), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n703), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n704), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n640), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFXL \block_reg[4][96]  ( .D(block_next[96]), .E(n635), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFXL \block_reg[0][96]  ( .D(block_next[96]), .E(n699), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFXL \block_reg[4][64]  ( .D(block_next[64]), .E(n637), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFXL \block_reg[0][64]  ( .D(block_next[64]), .E(n701), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n640), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n704), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[4][27]  ( .D(block_next[27]), .E(n640), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFX1 \block_reg[0][27]  ( .D(block_next[27]), .E(n704), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFXL \block_reg[4][127]  ( .D(block_next[127]), .E(n633), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFXL \block_reg[0][127]  ( .D(block_next[127]), .E(n697), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFXL \block_reg[4][124]  ( .D(block_next[124]), .E(n633), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFXL \block_reg[0][124]  ( .D(block_next[124]), .E(n697), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFXL \block_reg[4][125]  ( .D(block_next[125]), .E(n633), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFXL \block_reg[0][125]  ( .D(block_next[125]), .E(n697), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFXL \block_reg[4][126]  ( .D(block_next[126]), .E(n633), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFXL \block_reg[0][126]  ( .D(block_next[126]), .E(n697), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFXL \block_reg[4][123]  ( .D(block_next[123]), .E(n633), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFXL \block_reg[0][123]  ( .D(block_next[123]), .E(n697), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFX1 \block_reg[0][28]  ( .D(block_next[28]), .E(n704), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFX1 \block_reg[4][28]  ( .D(block_next[28]), .E(n640), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFX1 \block_reg[4][30]  ( .D(block_next[30]), .E(n640), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFX1 \block_reg[0][29]  ( .D(block_next[29]), .E(n704), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFX1 \block_reg[0][30]  ( .D(block_next[30]), .E(n704), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFX1 \block_reg[4][29]  ( .D(block_next[29]), .E(n640), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFX1 \block_reg[4][31]  ( .D(block_next[31]), .E(n640), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFX1 \block_reg[0][31]  ( .D(block_next[31]), .E(n704), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFXL \block_reg[1][113]  ( .D(block_next[113]), .E(n683), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFXL \block_reg[1][112]  ( .D(block_next[112]), .E(n683), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFXL \block_reg[1][90]  ( .D(block_next[90]), .E(n684), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFXL \block_reg[1][89]  ( .D(block_next[89]), .E(n684), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFXL \block_reg[1][88]  ( .D(block_next[88]), .E(n685), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFXL \block_reg[1][87]  ( .D(block_next[87]), .E(n685), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFXL \block_reg[1][84]  ( .D(block_next[84]), .E(n685), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFXL \block_reg[1][82]  ( .D(block_next[82]), .E(n685), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFXL \block_reg[1][81]  ( .D(block_next[81]), .E(n685), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFXL \block_reg[1][80]  ( .D(block_next[80]), .E(n685), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFX1 \block_reg[1][58]  ( .D(block_next[58]), .E(n687), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFX1 \block_reg[1][57]  ( .D(block_next[57]), .E(n687), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFX1 \block_reg[1][56]  ( .D(block_next[56]), .E(n687), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFX1 \block_reg[1][55]  ( .D(block_next[55]), .E(n687), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n687), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[1][50]  ( .D(block_next[50]), .E(n687), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n688), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[1][48]  ( .D(block_next[48]), .E(n688), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFX1 \block_reg[1][26]  ( .D(block_next[26]), .E(n689), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFX1 \block_reg[1][25]  ( .D(block_next[25]), .E(n689), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFX1 \block_reg[1][24]  ( .D(block_next[24]), .E(n689), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n690), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFXL \block_reg[1][122]  ( .D(block_next[122]), .E(n682), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFXL \block_reg[1][121]  ( .D(block_next[121]), .E(n682), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFXL \block_reg[1][120]  ( .D(block_next[120]), .E(n682), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFXL \block_reg[1][119]  ( .D(block_next[119]), .E(n682), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFXL \block_reg[1][118]  ( .D(block_next[118]), .E(n682), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFXL \block_reg[1][116]  ( .D(block_next[116]), .E(n682), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFXL \block_reg[1][114]  ( .D(block_next[114]), .E(n683), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFXL \block_reg[5][113]  ( .D(block_next[113]), .E(n616), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFXL \block_reg[5][112]  ( .D(block_next[112]), .E(n616), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFXL \block_reg[5][90]  ( .D(block_next[90]), .E(n617), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFXL \block_reg[5][89]  ( .D(block_next[89]), .E(n617), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFXL \block_reg[5][88]  ( .D(block_next[88]), .E(n618), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFXL \block_reg[5][87]  ( .D(block_next[87]), .E(n618), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFXL \block_reg[5][84]  ( .D(block_next[84]), .E(n618), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFXL \block_reg[5][82]  ( .D(block_next[82]), .E(n618), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFXL \block_reg[5][81]  ( .D(block_next[81]), .E(n618), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFXL \block_reg[5][80]  ( .D(block_next[80]), .E(n618), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFXL \block_reg[5][58]  ( .D(block_next[58]), .E(n620), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFXL \block_reg[5][57]  ( .D(block_next[57]), .E(n620), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFXL \block_reg[5][56]  ( .D(block_next[56]), .E(n620), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFXL \block_reg[5][55]  ( .D(block_next[55]), .E(n620), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFXL \block_reg[5][52]  ( .D(block_next[52]), .E(n620), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFXL \block_reg[5][50]  ( .D(block_next[50]), .E(n620), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFXL \block_reg[5][49]  ( .D(block_next[49]), .E(n621), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFXL \block_reg[5][48]  ( .D(block_next[48]), .E(n621), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFXL \block_reg[5][26]  ( .D(block_next[26]), .E(n622), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFXL \block_reg[5][25]  ( .D(block_next[25]), .E(n622), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFXL \block_reg[5][24]  ( .D(block_next[24]), .E(n622), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFXL \block_reg[5][23]  ( .D(block_next[23]), .E(n623), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFXL \block_reg[5][22]  ( .D(block_next[22]), .E(n623), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFXL \block_reg[5][20]  ( .D(block_next[20]), .E(n623), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFXL \block_reg[5][18]  ( .D(block_next[18]), .E(n623), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFXL \block_reg[5][17]  ( .D(block_next[17]), .E(n623), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFXL \block_reg[5][16]  ( .D(block_next[16]), .E(n623), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFXL \block_reg[5][122]  ( .D(block_next[122]), .E(n615), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFXL \block_reg[5][121]  ( .D(block_next[121]), .E(n615), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFXL \block_reg[5][120]  ( .D(block_next[120]), .E(n615), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFXL \block_reg[5][119]  ( .D(block_next[119]), .E(n615), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFXL \block_reg[5][118]  ( .D(block_next[118]), .E(n615), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFXL \block_reg[5][116]  ( .D(block_next[116]), .E(n615), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFXL \block_reg[5][114]  ( .D(block_next[114]), .E(n616), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFXL \block_reg[5][21]  ( .D(block_next[21]), .E(n623), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[1][54]  ( .D(block_next[54]), .E(n687), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFXL \block_reg[1][86]  ( .D(block_next[86]), .E(n685), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFXL \block_reg[5][54]  ( .D(block_next[54]), .E(n620), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFXL \block_reg[5][86]  ( .D(block_next[86]), .E(n618), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFXL \block_reg[1][117]  ( .D(block_next[117]), .E(n682), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFX1 \block_reg[1][51]  ( .D(block_next[51]), .E(n687), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n687), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFXL \block_reg[5][117]  ( .D(block_next[117]), .E(n615), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFXL \block_reg[1][115]  ( .D(block_next[115]), .E(n682), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFXL \block_reg[5][51]  ( .D(block_next[51]), .E(n620), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFXL \block_reg[5][53]  ( .D(block_next[53]), .E(n620), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFXL \block_reg[5][115]  ( .D(block_next[115]), .E(n615), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFXL \block_reg[1][85]  ( .D(block_next[85]), .E(n685), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFXL \block_reg[5][85]  ( .D(block_next[85]), .E(n618), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFXL \block_reg[5][19]  ( .D(block_next[19]), .E(n623), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFXL \block_reg[1][83]  ( .D(block_next[83]), .E(n685), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFXL \block_reg[5][83]  ( .D(block_next[83]), .E(n618), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFXL \block_reg[5][12]  ( .D(block_next[12]), .E(n623), .CK(clk), .Q(
        \block[5][12] ) );
  EDFFXL \block_reg[5][13]  ( .D(block_next[13]), .E(n623), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFXL \block_reg[1][109]  ( .D(block_next[109]), .E(n683), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFXL \block_reg[5][108]  ( .D(block_next[108]), .E(n616), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFXL \block_reg[5][10]  ( .D(block_next[10]), .E(n624), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFXL \block_reg[1][108]  ( .D(block_next[108]), .E(n683), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFXL \block_reg[5][109]  ( .D(block_next[109]), .E(n616), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFXL \block_reg[5][15]  ( .D(block_next[15]), .E(n623), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[5][45]  ( .D(block_next[45]), .E(n621), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFXL \block_reg[1][45]  ( .D(block_next[45]), .E(n688), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFXL \block_reg[1][76]  ( .D(block_next[76]), .E(n685), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFXL \block_reg[1][68]  ( .D(block_next[68]), .E(n686), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFXL \block_reg[1][110]  ( .D(block_next[110]), .E(n683), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFXL \block_reg[1][9]  ( .D(block_next[9]), .E(n691), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFXL \block_reg[5][14]  ( .D(block_next[14]), .E(n623), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFXL \block_reg[5][110]  ( .D(block_next[110]), .E(n616), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFXL \block_reg[5][104]  ( .D(block_next[104]), .E(n616), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFXL \block_reg[1][104]  ( .D(block_next[104]), .E(n683), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFX1 \block_reg[5][44]  ( .D(block_next[44]), .E(n621), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFXL \block_reg[5][77]  ( .D(block_next[77]), .E(n618), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFXL \block_reg[1][44]  ( .D(block_next[44]), .E(n688), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFXL \block_reg[5][11]  ( .D(block_next[11]), .E(n623), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFXL \block_reg[5][100]  ( .D(block_next[100]), .E(n617), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFXL \block_reg[1][100]  ( .D(block_next[100]), .E(n684), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFXL \block_reg[1][106]  ( .D(block_next[106]), .E(n683), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFXL \block_reg[5][106]  ( .D(block_next[106]), .E(n616), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFXL \block_reg[1][4]  ( .D(block_next[4]), .E(n691), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFXL \block_reg[1][73]  ( .D(block_next[73]), .E(n686), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFXL \block_reg[1][8]  ( .D(block_next[8]), .E(n691), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFXL \block_reg[5][102]  ( .D(block_next[102]), .E(n616), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFXL \block_reg[1][102]  ( .D(block_next[102]), .E(n683), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFXL \block_reg[5][105]  ( .D(block_next[105]), .E(n616), .CK(clk), .Q(
        \block[5][105] ) );
  EDFFXL \block_reg[1][72]  ( .D(block_next[72]), .E(n686), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFXL \block_reg[1][105]  ( .D(block_next[105]), .E(n683), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFX1 \block_reg[1][6]  ( .D(block_next[6]), .E(n691), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFXL \block_reg[5][6]  ( .D(block_next[6]), .E(n624), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFXL \block_reg[1][2]  ( .D(block_next[2]), .E(n691), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n622), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFXL \block_reg[1][36]  ( .D(block_next[36]), .E(n689), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFXL \block_reg[5][74]  ( .D(block_next[74]), .E(n619), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFXL \block_reg[1][70]  ( .D(block_next[70]), .E(n686), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFXL \block_reg[5][78]  ( .D(block_next[78]), .E(n618), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFX1 \block_reg[5][40]  ( .D(block_next[40]), .E(n621), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFXL \block_reg[1][40]  ( .D(block_next[40]), .E(n688), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFX1 \block_reg[1][46]  ( .D(block_next[46]), .E(n688), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFXL \block_reg[5][79]  ( .D(block_next[79]), .E(n618), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFXL \block_reg[5][46]  ( .D(block_next[46]), .E(n621), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFXL \block_reg[1][111]  ( .D(block_next[111]), .E(n683), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n621), .CK(clk), .Q(
        \block[5][41] ) );
  EDFFXL \block_reg[1][41]  ( .D(block_next[41]), .E(n688), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[1][42]  ( .D(block_next[42]), .E(n688), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFXL \block_reg[1][1]  ( .D(block_next[1]), .E(n691), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n621), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFXL \block_reg[1][38]  ( .D(block_next[38]), .E(n688), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFXL \block_reg[5][111]  ( .D(block_next[111]), .E(n616), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFXL \block_reg[5][107]  ( .D(block_next[107]), .E(n616), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFXL \block_reg[1][107]  ( .D(block_next[107]), .E(n683), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFXL \block_reg[5][42]  ( .D(block_next[42]), .E(n621), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFX1 \block_reg[1][47]  ( .D(block_next[47]), .E(n688), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFXL \block_reg[5][98]  ( .D(block_next[98]), .E(n617), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFXL \block_reg[1][98]  ( .D(block_next[98]), .E(n684), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFXL \block_reg[5][47]  ( .D(block_next[47]), .E(n621), .CK(clk), .Q(
        \block[5][47] ) );
  EDFFXL \block_reg[5][97]  ( .D(block_next[97]), .E(n617), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFXL \block_reg[1][97]  ( .D(block_next[97]), .E(n684), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFX1 \block_reg[5][33]  ( .D(block_next[33]), .E(n622), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFXL \block_reg[1][33]  ( .D(block_next[33]), .E(n689), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFXL \block_reg[5][75]  ( .D(block_next[75]), .E(n619), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFX1 \block_reg[5][43]  ( .D(block_next[43]), .E(n621), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFXL \block_reg[1][43]  ( .D(block_next[43]), .E(n688), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFXL \block_reg[5][66]  ( .D(block_next[66]), .E(n619), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFX1 \block_reg[1][65]  ( .D(block_next[65]), .E(n686), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFXL \block_reg[5][65]  ( .D(block_next[65]), .E(n619), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFX1 \block_reg[1][34]  ( .D(block_next[34]), .E(n689), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFXL \block_reg[5][34]  ( .D(block_next[34]), .E(n622), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFXL \block_reg[5][3]  ( .D(block_next[3]), .E(n624), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFXL \block_reg[5][103]  ( .D(block_next[103]), .E(n616), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFXL \block_reg[1][103]  ( .D(block_next[103]), .E(n683), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFX1 \block_reg[5][39]  ( .D(block_next[39]), .E(n621), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFXL \block_reg[1][39]  ( .D(block_next[39]), .E(n688), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFXL \block_reg[5][67]  ( .D(block_next[67]), .E(n619), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFXL \block_reg[5][99]  ( .D(block_next[99]), .E(n617), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFXL \block_reg[1][99]  ( .D(block_next[99]), .E(n684), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFXL \block_reg[1][7]  ( .D(block_next[7]), .E(n691), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFXL \block_reg[1][71]  ( .D(block_next[71]), .E(n686), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFXL \block_reg[5][101]  ( .D(block_next[101]), .E(n617), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFXL \block_reg[1][101]  ( .D(block_next[101]), .E(n684), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFXL \block_reg[1][0]  ( .D(block_next[0]), .E(n691), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFXL \block_reg[1][69]  ( .D(block_next[69]), .E(n686), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFXL \block_reg[1][5]  ( .D(block_next[5]), .E(n691), .CK(clk), .Q(
        \block[1][5] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n621), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFXL \block_reg[1][37]  ( .D(block_next[37]), .E(n688), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(n689), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFXL \block_reg[5][35]  ( .D(block_next[35]), .E(n622), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFXL \block_reg[5][96]  ( .D(block_next[96]), .E(n617), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFXL \block_reg[1][96]  ( .D(block_next[96]), .E(n684), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFX1 \block_reg[5][64]  ( .D(block_next[64]), .E(n619), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFXL \block_reg[1][64]  ( .D(block_next[64]), .E(n686), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n622), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFXL \block_reg[1][32]  ( .D(block_next[32]), .E(n689), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[5][27]  ( .D(block_next[27]), .E(n622), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFXL \block_reg[1][27]  ( .D(block_next[27]), .E(n689), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFXL \block_reg[5][127]  ( .D(block_next[127]), .E(n615), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFXL \block_reg[1][127]  ( .D(block_next[127]), .E(n682), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFXL \block_reg[5][124]  ( .D(block_next[124]), .E(n615), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFXL \block_reg[1][124]  ( .D(block_next[124]), .E(n682), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFXL \block_reg[5][125]  ( .D(block_next[125]), .E(n615), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFXL \block_reg[1][125]  ( .D(block_next[125]), .E(n682), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFXL \block_reg[5][126]  ( .D(block_next[126]), .E(n615), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFXL \block_reg[1][126]  ( .D(block_next[126]), .E(n682), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFXL \block_reg[5][123]  ( .D(block_next[123]), .E(n615), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFXL \block_reg[1][123]  ( .D(block_next[123]), .E(n682), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFX1 \block_reg[1][28]  ( .D(block_next[28]), .E(n689), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFX1 \block_reg[5][30]  ( .D(block_next[30]), .E(n622), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFXL \block_reg[1][30]  ( .D(block_next[30]), .E(n689), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFXL \block_reg[5][28]  ( .D(block_next[28]), .E(n622), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFX1 \block_reg[1][29]  ( .D(block_next[29]), .E(n689), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFXL \block_reg[5][29]  ( .D(block_next[29]), .E(n622), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFX1 \block_reg[5][31]  ( .D(block_next[31]), .E(n622), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFXL \block_reg[1][31]  ( .D(block_next[31]), .E(n689), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n677), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n612), .CK(clk), .QN(
        n535) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(n75), .E(n677), .CK(clk), .Q(
        \blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(n75), .E(n612), .CK(clk), .QN(n420) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(n72), .E(n678), .CK(clk), .QN(n108) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(n677), .CK(clk), 
        .Q(\blocktag[2][16] ) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(n76), .E(n612), .CK(clk), .QN(n510) );
  EDFFXL \block_reg[6][91]  ( .D(block_next[91]), .E(n604), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFXL \block_reg[2][91]  ( .D(block_next[91]), .E(n669), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFXL \block_reg[2][92]  ( .D(block_next[92]), .E(n669), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFXL \block_reg[6][92]  ( .D(block_next[92]), .E(n604), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFX1 \block_reg[6][62]  ( .D(block_next[62]), .E(n607), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFX1 \block_reg[2][62]  ( .D(block_next[62]), .E(n672), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFX1 \block_reg[2][61]  ( .D(block_next[61]), .E(n672), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFX1 \block_reg[6][61]  ( .D(block_next[61]), .E(n607), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFXL \block_reg[6][94]  ( .D(block_next[94]), .E(n604), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFXL \block_reg[2][94]  ( .D(block_next[94]), .E(n669), .CK(clk), .Q(
        \block[2][94] ) );
  EDFFXL \block_reg[6][95]  ( .D(block_next[95]), .E(n604), .CK(clk), .Q(
        \block[6][95] ) );
  EDFFXL \block_reg[2][95]  ( .D(block_next[95]), .E(n669), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFX1 \block_reg[6][59]  ( .D(block_next[59]), .E(n607), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFX1 \block_reg[2][59]  ( .D(block_next[59]), .E(n672), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFX1 \block_reg[2][60]  ( .D(block_next[60]), .E(n672), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFXL \block_reg[2][93]  ( .D(block_next[93]), .E(n669), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFX1 \block_reg[6][60]  ( .D(block_next[60]), .E(n607), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFXL \block_reg[6][93]  ( .D(block_next[93]), .E(n604), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n677), .CK(clk), 
        .Q(\blocktag[2][20] ) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n612), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n677), .CK(clk), 
        .Q(\blocktag[2][19] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n613), .CK(clk), .QN(
        n460) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n612), .CK(clk), 
        .Q(\blocktag[6][19] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n678), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n677), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n612), .CK(clk), 
        .QN(n455) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(n68), .E(n677), .CK(clk), .QN(n410) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(n68), .E(n612), .CK(clk), .QN(n433) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n677), .CK(clk), 
        .Q(\blocktag[2][21] ) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n612), .CK(clk), 
        .Q(\blocktag[6][21] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(blocktag_next[7]), .E(n678), .CK(clk), .Q(
        \blocktag[2][7] ) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(blocktag_next[7]), .E(n613), .CK(clk), .QN(
        n50) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n678), .CK(clk), .Q(
        \blocktag[2][4] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n678), .CK(clk), .QN(
        n426) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n613), .CK(clk), .QN(
        n449) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n613), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(n69), .E(n676), .CK(clk), .QN(n507) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(n69), .E(n611), .CK(clk), .QN(n464) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n677), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n612), .CK(clk), .Q(
        \blocktag[6][0] ) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n676), .CK(clk), 
        .Q(\blocktag[2][24] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n611), .CK(clk), 
        .Q(\blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n678), .CK(clk), .QN(
        n517) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n661), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n595), .CK(clk), .QN(
        n537) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(n75), .E(n661), .CK(clk), .Q(
        \blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(n75), .E(n595), .CK(clk), .QN(n422) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(n72), .E(n662), .CK(clk), .QN(n110) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(n661), .CK(clk), 
        .Q(\blocktag[3][16] ) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(n76), .E(n595), .CK(clk), .QN(n512) );
  EDFFXL \block_reg[7][91]  ( .D(block_next[91]), .E(n589), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFXL \block_reg[3][91]  ( .D(block_next[91]), .E(n653), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFXL \block_reg[3][92]  ( .D(block_next[92]), .E(n653), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFX1 \block_reg[3][62]  ( .D(block_next[62]), .E(n656), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFXL \block_reg[7][92]  ( .D(block_next[92]), .E(n589), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFX1 \block_reg[3][61]  ( .D(block_next[61]), .E(n656), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFX1 \block_reg[7][61]  ( .D(block_next[61]), .E(n592), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFXL \block_reg[3][94]  ( .D(block_next[94]), .E(n653), .CK(clk), .Q(
        \block[3][94] ) );
  EDFFXL \block_reg[7][94]  ( .D(block_next[94]), .E(n589), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFXL \block_reg[3][95]  ( .D(block_next[95]), .E(n653), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFXL \block_reg[7][95]  ( .D(block_next[95]), .E(n589), .CK(clk), .Q(
        \block[7][95] ) );
  EDFFX1 \block_reg[7][59]  ( .D(block_next[59]), .E(n592), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFX1 \block_reg[3][59]  ( .D(block_next[59]), .E(n656), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFX1 \block_reg[3][60]  ( .D(block_next[60]), .E(n656), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFXL \block_reg[3][93]  ( .D(block_next[93]), .E(n653), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFX1 \block_reg[7][60]  ( .D(block_next[60]), .E(n592), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFXL \block_reg[7][93]  ( .D(block_next[93]), .E(n589), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n661), .CK(clk), 
        .Q(\blocktag[3][20] ) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n595), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n661), .CK(clk), 
        .Q(\blocktag[3][19] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n596), .CK(clk), .QN(
        n462) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n595), .CK(clk), 
        .Q(\blocktag[7][19] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n662), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n661), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n595), .CK(clk), 
        .QN(n457) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(n68), .E(n661), .CK(clk), .QN(n412) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(n68), .E(n595), .CK(clk), .QN(n431) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n661), .CK(clk), 
        .Q(\blocktag[3][21] ) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n595), .CK(clk), 
        .Q(\blocktag[7][21] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(blocktag_next[7]), .E(n662), .CK(clk), .Q(
        \blocktag[3][7] ) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(blocktag_next[7]), .E(n596), .CK(clk), .QN(
        n48) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(n662), .CK(clk), .Q(
        \blocktag[3][4] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(n662), .CK(clk), .QN(
        n428) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(n596), .CK(clk), .QN(
        n451) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(n596), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(n69), .E(n660), .CK(clk), .QN(n509) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(n69), .E(n597), .CK(clk), .QN(n466) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n661), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n595), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n660), .CK(clk), 
        .Q(\blocktag[3][24] ) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n597), .CK(clk), 
        .Q(\blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(n662), .CK(clk), .QN(
        n515) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n707), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n643), .CK(clk), .QN(
        n536) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(n75), .E(n707), .CK(clk), .Q(
        \blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(n75), .E(n643), .CK(clk), .QN(n421) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(n72), .E(n708), .CK(clk), .QN(n109) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(n707), .CK(clk), 
        .Q(\blocktag[0][16] ) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(n76), .E(n643), .CK(clk), .QN(n511) );
  EDFFXL \block_reg[4][91]  ( .D(block_next[91]), .E(n635), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFXL \block_reg[0][91]  ( .D(block_next[91]), .E(n699), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFXL \block_reg[0][92]  ( .D(block_next[92]), .E(n699), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFXL \block_reg[4][92]  ( .D(block_next[92]), .E(n635), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFX1 \block_reg[4][62]  ( .D(block_next[62]), .E(n638), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFX1 \block_reg[0][62]  ( .D(block_next[62]), .E(n702), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFX1 \block_reg[0][61]  ( .D(block_next[61]), .E(n702), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFX1 \block_reg[4][61]  ( .D(block_next[61]), .E(n638), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFXL \block_reg[4][94]  ( .D(block_next[94]), .E(n635), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFXL \block_reg[0][94]  ( .D(block_next[94]), .E(n699), .CK(clk), .Q(
        \block[0][94] ) );
  EDFFXL \block_reg[4][95]  ( .D(block_next[95]), .E(n635), .CK(clk), .Q(
        \block[4][95] ) );
  EDFFXL \block_reg[0][95]  ( .D(block_next[95]), .E(n699), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFX1 \block_reg[4][59]  ( .D(block_next[59]), .E(n638), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFX1 \block_reg[0][59]  ( .D(block_next[59]), .E(n702), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFX1 \block_reg[0][60]  ( .D(block_next[60]), .E(n702), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFXL \block_reg[0][93]  ( .D(block_next[93]), .E(n699), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFX1 \block_reg[4][60]  ( .D(block_next[60]), .E(n638), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFXL \block_reg[4][93]  ( .D(block_next[93]), .E(n635), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n707), .CK(clk), 
        .Q(\blocktag[0][20] ) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n643), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n707), .CK(clk), 
        .Q(\blocktag[0][19] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n644), .CK(clk), .QN(
        n459) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n643), .CK(clk), 
        .Q(\blocktag[4][19] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n708), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n707), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n643), .CK(clk), 
        .QN(n454) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(n68), .E(n707), .CK(clk), .QN(n411) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(n68), .E(n643), .CK(clk), .QN(n434) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n707), .CK(clk), 
        .Q(\blocktag[0][21] ) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n643), .CK(clk), 
        .Q(\blocktag[4][21] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(blocktag_next[7]), .E(n708), .CK(clk), .Q(
        \blocktag[0][7] ) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(blocktag_next[7]), .E(n644), .CK(clk), .QN(
        n51) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n708), .CK(clk), .Q(
        \blocktag[0][4] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n708), .CK(clk), .QN(
        n425) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n644), .CK(clk), .QN(
        n450) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n644), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(n69), .E(n706), .CK(clk), .QN(n506) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(n69), .E(n642), .CK(clk), .QN(n463) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n707), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n643), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n706), .CK(clk), 
        .Q(\blocktag[0][24] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n642), .CK(clk), 
        .Q(\blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n708), .CK(clk), .QN(
        n518) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n692), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n625), .CK(clk), .QN(
        n538) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(n75), .E(n692), .CK(clk), .Q(
        \blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(n75), .E(n625), .CK(clk), .QN(n423) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(n72), .E(n693), .CK(clk), .QN(n111) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n692), .CK(clk), 
        .Q(\blocktag[1][16] ) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(n76), .E(n625), .CK(clk), .QN(n513) );
  EDFFXL \block_reg[5][91]  ( .D(block_next[91]), .E(n617), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFXL \block_reg[1][91]  ( .D(block_next[91]), .E(n684), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFX1 \block_reg[5][62]  ( .D(block_next[62]), .E(n620), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFXL \block_reg[1][92]  ( .D(block_next[92]), .E(n684), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFXL \block_reg[1][62]  ( .D(block_next[62]), .E(n687), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFXL \block_reg[5][92]  ( .D(block_next[92]), .E(n617), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFX1 \block_reg[1][61]  ( .D(block_next[61]), .E(n687), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFXL \block_reg[5][61]  ( .D(block_next[61]), .E(n620), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFXL \block_reg[1][94]  ( .D(block_next[94]), .E(n684), .CK(clk), .Q(
        \block[1][94] ) );
  EDFFXL \block_reg[5][94]  ( .D(block_next[94]), .E(n617), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFXL \block_reg[1][95]  ( .D(block_next[95]), .E(n684), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFXL \block_reg[5][95]  ( .D(block_next[95]), .E(n617), .CK(clk), .Q(
        \block[5][95] ) );
  EDFFX1 \block_reg[5][59]  ( .D(block_next[59]), .E(n620), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFXL \block_reg[1][59]  ( .D(block_next[59]), .E(n687), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFX1 \block_reg[1][60]  ( .D(block_next[60]), .E(n687), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFXL \block_reg[1][93]  ( .D(block_next[93]), .E(n684), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFXL \block_reg[1][63]  ( .D(block_next[63]), .E(n686), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFXL \block_reg[5][60]  ( .D(block_next[60]), .E(n620), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFXL \block_reg[5][93]  ( .D(block_next[93]), .E(n617), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n692), .CK(clk), 
        .Q(\blocktag[1][20] ) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n625), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n692), .CK(clk), 
        .Q(\blocktag[1][19] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n626), .CK(clk), .QN(
        n461) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n625), .CK(clk), 
        .Q(\blocktag[5][19] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n693), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n692), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n625), .CK(clk), 
        .QN(n456) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(n68), .E(n692), .CK(clk), .QN(n413) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(n68), .E(n625), .CK(clk), .QN(n432) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n692), .CK(clk), 
        .Q(\blocktag[1][21] ) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n625), .CK(clk), 
        .Q(\blocktag[5][21] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(blocktag_next[7]), .E(n693), .CK(clk), .Q(
        \blocktag[1][7] ) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(blocktag_next[7]), .E(n626), .CK(clk), .QN(
        n49) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(n693), .CK(clk), .Q(
        \blocktag[1][4] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(n693), .CK(clk), .QN(
        n427) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n626), .CK(clk), .QN(
        n452) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n626), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(n69), .E(n691), .CK(clk), .QN(n508) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(n69), .E(n624), .CK(clk), .QN(n465) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n692), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(n625), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n691), .CK(clk), 
        .Q(\blocktag[1][24] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n624), .CK(clk), 
        .Q(\blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(n693), .CK(clk), .QN(
        n516) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n1725), .CK(clk), .RN(n794), .Q(
        blockdirty[2]), .QN(n1741) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n1721), .CK(clk), .RN(n794), .Q(
        blockdirty[6]), .QN(n1737) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n1724), .CK(clk), .RN(n794), .Q(
        blockdirty[3]), .QN(n1740) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n1720), .CK(clk), .RN(n794), .Q(
        blockdirty[7]), .QN(n1736) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n1727), .CK(clk), .RN(n794), .Q(
        blockdirty[0]), .QN(n1743) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n1723), .CK(clk), .RN(n794), .Q(
        blockdirty[4]), .QN(n1739) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n1726), .CK(clk), .RN(n794), .Q(
        blockdirty[1]), .QN(n1742) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n1722), .CK(clk), .RN(n794), .Q(
        blockdirty[5]), .QN(n1738) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n678), .CK(clk), .Q(
        \blocktag[2][3] ) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n613), .CK(clk), .Q(
        \blocktag[6][3] ) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(n678), .CK(clk), 
        .Q(\blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(n74), .E(n677), .CK(clk), .Q(
        \blocktag[2][12] ) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(n74), .E(n612), .CK(clk), .Q(
        \blocktag[6][12] ) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n662), .CK(clk), .Q(
        \blocktag[3][3] ) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n596), .CK(clk), .Q(
        \blocktag[7][3] ) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(n662), .CK(clk), 
        .Q(\blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(n74), .E(n661), .CK(clk), .Q(
        \blocktag[3][12] ) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(n74), .E(n595), .CK(clk), .Q(
        \blocktag[7][12] ) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n708), .CK(clk), .Q(
        \blocktag[0][3] ) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n644), .CK(clk), .Q(
        \blocktag[4][3] ) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(n708), .CK(clk), 
        .Q(\blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(n74), .E(n707), .CK(clk), .Q(
        \blocktag[0][12] ) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(n74), .E(n643), .CK(clk), .Q(
        \blocktag[4][12] ) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n693), .CK(clk), .Q(
        \blocktag[1][3] ) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n626), .CK(clk), .Q(
        \blocktag[5][3] ) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n693), .CK(clk), 
        .Q(\blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(n74), .E(n692), .CK(clk), .Q(
        \blocktag[1][12] ) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(n74), .E(n625), .CK(clk), .Q(
        \blocktag[5][12] ) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n707), .CK(clk), 
        .QN(n66) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n677), .CK(clk), 
        .QN(n77) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n643), .CK(clk), 
        .Q(\blocktag[4][22] ) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n612), .CK(clk), 
        .Q(\blocktag[6][22] ) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n661), .CK(clk), 
        .QN(n71) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n692), .CK(clk), 
        .QN(n62) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n595), .CK(clk), 
        .Q(\blocktag[7][22] ) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n625), .CK(clk), 
        .Q(\blocktag[5][22] ) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n1719), .CK(clk), .RN(n795), .Q(
        blockvalid[0]), .QN(n1735) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n1718), .CK(clk), .RN(n795), .Q(
        blockvalid[1]), .QN(n1734) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n1714), .CK(clk), .RN(n795), .Q(
        blockvalid[5]), .QN(n1730) );
  EDFFXL \block_reg[1][66]  ( .D(block_next[66]), .E(n686), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFXL \blocktag_reg[7][17]  ( .D(n73), .E(n56), .CK(clk), .Q(
        \blocktag[7][17] ) );
  EDFFXL \blocktag_reg[6][17]  ( .D(n73), .E(n55), .CK(clk), .Q(
        \blocktag[6][17] ) );
  EDFFXL \blocktag_reg[5][17]  ( .D(n73), .E(n64), .CK(clk), .Q(
        \blocktag[5][17] ) );
  EDFFXL \blocktag_reg[4][17]  ( .D(n73), .E(n61), .CK(clk), .Q(
        \blocktag[4][17] ) );
  EDFFXL \blocktag_reg[3][17]  ( .D(n73), .E(n54), .CK(clk), .Q(
        \blocktag[3][17] ) );
  EDFFXL \blocktag_reg[2][17]  ( .D(n73), .E(n52), .CK(clk), .Q(
        \blocktag[2][17] ) );
  EDFFXL \blocktag_reg[1][17]  ( .D(n73), .E(n53), .CK(clk), .Q(
        \blocktag[1][17] ) );
  EDFFXL \blocktag_reg[0][17]  ( .D(n73), .E(n1711), .CK(clk), .Q(
        \blocktag[0][17] ) );
  EDFFXL \block_reg[5][76]  ( .D(block_next[76]), .E(n64), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFXL \block_reg[5][73]  ( .D(block_next[73]), .E(n64), .CK(clk), .Q(
        \block[5][73] ) );
  EDFFXL \block_reg[5][72]  ( .D(block_next[72]), .E(n64), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFXL \block_reg[5][71]  ( .D(block_next[71]), .E(n64), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFXL \block_reg[5][70]  ( .D(block_next[70]), .E(n64), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFXL \block_reg[5][69]  ( .D(block_next[69]), .E(n64), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFXL \block_reg[5][68]  ( .D(block_next[68]), .E(n64), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFXL \block_reg[1][75]  ( .D(block_next[75]), .E(n53), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFXL \block_reg[1][74]  ( .D(block_next[74]), .E(n53), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFXL \block_reg[1][67]  ( .D(block_next[67]), .E(n53), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFXL \block_reg[7][63]  ( .D(block_next[63]), .E(n56), .CK(clk), .Q(
        \block[7][63] ) );
  EDFFXL \block_reg[6][63]  ( .D(block_next[63]), .E(n55), .CK(clk), .Q(
        \block[6][63] ) );
  EDFFXL \block_reg[5][63]  ( .D(block_next[63]), .E(n64), .CK(clk), .Q(
        \block[5][63] ) );
  EDFFXL \block_reg[4][63]  ( .D(block_next[63]), .E(n61), .CK(clk), .Q(
        \block[4][63] ) );
  EDFFXL \block_reg[3][63]  ( .D(block_next[63]), .E(n54), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFXL \block_reg[2][63]  ( .D(block_next[63]), .E(n52), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFXL \block_reg[0][63]  ( .D(block_next[63]), .E(n1711), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFXL \block_reg[1][79]  ( .D(block_next[79]), .E(n53), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFXL \block_reg[1][78]  ( .D(block_next[78]), .E(n53), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFXL \block_reg[1][77]  ( .D(block_next[77]), .E(n53), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFXL \block_reg[7][26]  ( .D(block_next[26]), .E(n56), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFXL \block_reg[7][25]  ( .D(block_next[25]), .E(n56), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFXL \block_reg[7][24]  ( .D(block_next[24]), .E(n56), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFXL \block_reg[7][23]  ( .D(block_next[23]), .E(n56), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFXL \block_reg[7][22]  ( .D(block_next[22]), .E(n56), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFXL \block_reg[7][21]  ( .D(block_next[21]), .E(n56), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFXL \block_reg[7][20]  ( .D(block_next[20]), .E(n56), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFXL \block_reg[7][19]  ( .D(block_next[19]), .E(n56), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFXL \block_reg[7][18]  ( .D(block_next[18]), .E(n56), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFXL \block_reg[7][17]  ( .D(block_next[17]), .E(n56), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFXL \block_reg[7][16]  ( .D(block_next[16]), .E(n56), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFXL \block_reg[7][15]  ( .D(block_next[15]), .E(n56), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFXL \block_reg[7][14]  ( .D(block_next[14]), .E(n56), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFXL \block_reg[7][13]  ( .D(block_next[13]), .E(n56), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFXL \block_reg[7][12]  ( .D(block_next[12]), .E(n56), .CK(clk), .Q(
        \block[7][12] ) );
  EDFFXL \block_reg[7][11]  ( .D(block_next[11]), .E(n56), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFXL \block_reg[7][10]  ( .D(block_next[10]), .E(n56), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFXL \block_reg[7][9]  ( .D(block_next[9]), .E(n56), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFXL \block_reg[7][8]  ( .D(block_next[8]), .E(n56), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFXL \block_reg[7][7]  ( .D(block_next[7]), .E(n56), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFXL \block_reg[7][6]  ( .D(block_next[6]), .E(n56), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFXL \block_reg[7][5]  ( .D(block_next[5]), .E(n56), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFXL \block_reg[7][4]  ( .D(block_next[4]), .E(n56), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFXL \block_reg[7][3]  ( .D(block_next[3]), .E(n56), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFXL \block_reg[7][2]  ( .D(block_next[2]), .E(n56), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFXL \block_reg[7][1]  ( .D(block_next[1]), .E(n56), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFXL \block_reg[6][26]  ( .D(block_next[26]), .E(n55), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFXL \block_reg[6][25]  ( .D(block_next[25]), .E(n55), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFXL \block_reg[6][24]  ( .D(block_next[24]), .E(n55), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFXL \block_reg[7][62]  ( .D(block_next[62]), .E(n592), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFX2 \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n644), .CK(clk), .QN(
        n117) );
  EDFFX2 \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n613), .CK(clk), .QN(
        n116) );
  EDFFX2 \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n626), .CK(clk), .QN(
        n115) );
  EDFFX2 \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n596), .CK(clk), .QN(
        n114) );
  EDFFX2 \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n626), .CK(clk), 
        .Q(n90) );
  EDFFX2 \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n596), .CK(clk), 
        .Q(n89) );
  EDFFX2 \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(n644), .CK(clk), 
        .Q(n88) );
  EDFFX2 \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n613), .CK(clk), 
        .Q(n87) );
  EDFFX4 \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(n595), .CK(clk), 
        .Q(n84) );
  EDFFX4 \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(n625), .CK(clk), 
        .Q(n83) );
  EDFFX4 \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n612), .CK(clk), 
        .Q(n82) );
  EDFFX4 \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(n643), .CK(clk), 
        .Q(n81) );
  EDFFXL \block_reg[6][7]  ( .D(block_next[7]), .E(n611), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFXL \block_reg[5][7]  ( .D(block_next[7]), .E(n624), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFXL \block_reg[4][7]  ( .D(block_next[7]), .E(n642), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFXL \block_reg[0][7]  ( .D(block_next[7]), .E(n706), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFXL \block_reg[3][7]  ( .D(block_next[7]), .E(n660), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFXL \block_reg[2][7]  ( .D(block_next[7]), .E(n676), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFXL \block_reg[6][22]  ( .D(block_next[22]), .E(n55), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFXL \block_reg[4][22]  ( .D(block_next[22]), .E(n641), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFXL \block_reg[3][22]  ( .D(block_next[22]), .E(n659), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFXL \block_reg[1][22]  ( .D(block_next[22]), .E(n690), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFXL \block_reg[0][22]  ( .D(block_next[22]), .E(n705), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFXL \block_reg[2][22]  ( .D(block_next[22]), .E(n675), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFXL \block_reg[6][11]  ( .D(block_next[11]), .E(n610), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFXL \block_reg[4][11]  ( .D(block_next[11]), .E(n641), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFXL \block_reg[1][11]  ( .D(block_next[11]), .E(n690), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFXL \block_reg[0][11]  ( .D(block_next[11]), .E(n705), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFXL \block_reg[3][11]  ( .D(block_next[11]), .E(n659), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFXL \block_reg[2][11]  ( .D(block_next[11]), .E(n675), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFXL \block_reg[6][23]  ( .D(block_next[23]), .E(n55), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFXL \block_reg[4][23]  ( .D(block_next[23]), .E(n641), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFXL \block_reg[3][23]  ( .D(block_next[23]), .E(n659), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFXL \block_reg[1][23]  ( .D(block_next[23]), .E(n690), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFXL \block_reg[0][23]  ( .D(block_next[23]), .E(n705), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFXL \block_reg[2][23]  ( .D(block_next[23]), .E(n675), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFXL \block_reg[6][10]  ( .D(block_next[10]), .E(n611), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFXL \block_reg[4][10]  ( .D(block_next[10]), .E(n642), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFXL \block_reg[1][10]  ( .D(block_next[10]), .E(n691), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFXL \block_reg[0][10]  ( .D(block_next[10]), .E(n706), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFXL \block_reg[3][10]  ( .D(block_next[10]), .E(n660), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFXL \block_reg[2][10]  ( .D(block_next[10]), .E(n676), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFXL \block_reg[6][19]  ( .D(block_next[19]), .E(n610), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFXL \block_reg[4][19]  ( .D(block_next[19]), .E(n641), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFXL \block_reg[3][19]  ( .D(block_next[19]), .E(n659), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFXL \block_reg[1][19]  ( .D(block_next[19]), .E(n690), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFXL \block_reg[0][19]  ( .D(block_next[19]), .E(n705), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFXL \block_reg[2][19]  ( .D(block_next[19]), .E(n675), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFXL \block_reg[6][3]  ( .D(block_next[3]), .E(n611), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFXL \block_reg[4][3]  ( .D(block_next[3]), .E(n642), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFXL \block_reg[1][3]  ( .D(block_next[3]), .E(n691), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFXL \block_reg[0][3]  ( .D(block_next[3]), .E(n706), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFXL \block_reg[3][3]  ( .D(block_next[3]), .E(n660), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFXL \block_reg[2][3]  ( .D(block_next[3]), .E(n676), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFXL \block_reg[6][13]  ( .D(block_next[13]), .E(n610), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFXL \block_reg[4][13]  ( .D(block_next[13]), .E(n641), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFXL \block_reg[1][13]  ( .D(block_next[13]), .E(n690), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFXL \block_reg[0][13]  ( .D(block_next[13]), .E(n705), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFXL \block_reg[3][13]  ( .D(block_next[13]), .E(n659), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFXL \block_reg[2][13]  ( .D(block_next[13]), .E(n675), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFXL \block_reg[6][8]  ( .D(block_next[8]), .E(n611), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFXL \block_reg[5][8]  ( .D(block_next[8]), .E(n624), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFXL \block_reg[4][8]  ( .D(block_next[8]), .E(n642), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFXL \block_reg[0][8]  ( .D(block_next[8]), .E(n706), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFXL \block_reg[3][8]  ( .D(block_next[8]), .E(n660), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFXL \block_reg[2][8]  ( .D(block_next[8]), .E(n676), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFXL \block_reg[6][12]  ( .D(block_next[12]), .E(n610), .CK(clk), .Q(
        \block[6][12] ) );
  EDFFXL \block_reg[4][12]  ( .D(block_next[12]), .E(n641), .CK(clk), .Q(
        \block[4][12] ) );
  EDFFXL \block_reg[1][12]  ( .D(block_next[12]), .E(n690), .CK(clk), .Q(
        \block[1][12] ) );
  EDFFXL \block_reg[0][12]  ( .D(block_next[12]), .E(n705), .CK(clk), .Q(
        \block[0][12] ) );
  EDFFXL \block_reg[3][12]  ( .D(block_next[12]), .E(n659), .CK(clk), .Q(
        \block[3][12] ) );
  EDFFXL \block_reg[2][12]  ( .D(block_next[12]), .E(n675), .CK(clk), .Q(
        \block[2][12] ) );
  EDFFXL \block_reg[6][2]  ( .D(block_next[2]), .E(n611), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFXL \block_reg[5][2]  ( .D(block_next[2]), .E(n624), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFXL \block_reg[4][2]  ( .D(block_next[2]), .E(n642), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFXL \block_reg[0][2]  ( .D(block_next[2]), .E(n706), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFXL \block_reg[3][2]  ( .D(block_next[2]), .E(n660), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFXL \block_reg[2][2]  ( .D(block_next[2]), .E(n676), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFXL \block_reg[6][17]  ( .D(block_next[17]), .E(n610), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFXL \block_reg[4][17]  ( .D(block_next[17]), .E(n641), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFXL \block_reg[3][17]  ( .D(block_next[17]), .E(n659), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFXL \block_reg[1][17]  ( .D(block_next[17]), .E(n690), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFXL \block_reg[0][17]  ( .D(block_next[17]), .E(n705), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFXL \block_reg[2][17]  ( .D(block_next[17]), .E(n675), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFXL \block_reg[6][4]  ( .D(block_next[4]), .E(n611), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFXL \block_reg[5][4]  ( .D(block_next[4]), .E(n624), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFXL \block_reg[4][4]  ( .D(block_next[4]), .E(n642), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFXL \block_reg[0][4]  ( .D(block_next[4]), .E(n706), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFXL \block_reg[3][4]  ( .D(block_next[4]), .E(n660), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFXL \block_reg[2][4]  ( .D(block_next[4]), .E(n676), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFXL \block_reg[6][15]  ( .D(block_next[15]), .E(n610), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFXL \block_reg[4][15]  ( .D(block_next[15]), .E(n641), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFXL \block_reg[1][15]  ( .D(block_next[15]), .E(n690), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFXL \block_reg[0][15]  ( .D(block_next[15]), .E(n705), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFXL \block_reg[3][15]  ( .D(block_next[15]), .E(n659), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFXL \block_reg[2][15]  ( .D(block_next[15]), .E(n675), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFXL \block_reg[6][9]  ( .D(block_next[9]), .E(n611), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFXL \block_reg[5][9]  ( .D(block_next[9]), .E(n624), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFXL \block_reg[4][9]  ( .D(block_next[9]), .E(n642), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFXL \block_reg[0][9]  ( .D(block_next[9]), .E(n706), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFXL \block_reg[3][9]  ( .D(block_next[9]), .E(n660), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFXL \block_reg[2][9]  ( .D(block_next[9]), .E(n676), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFXL \block_reg[6][14]  ( .D(block_next[14]), .E(n610), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFXL \block_reg[4][14]  ( .D(block_next[14]), .E(n641), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFXL \block_reg[1][14]  ( .D(block_next[14]), .E(n690), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFXL \block_reg[0][14]  ( .D(block_next[14]), .E(n705), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFXL \block_reg[3][14]  ( .D(block_next[14]), .E(n659), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFXL \block_reg[2][14]  ( .D(block_next[14]), .E(n675), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFXL \block_reg[6][5]  ( .D(block_next[5]), .E(n611), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFXL \block_reg[5][5]  ( .D(block_next[5]), .E(n624), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFXL \block_reg[4][5]  ( .D(block_next[5]), .E(n642), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFXL \block_reg[0][5]  ( .D(block_next[5]), .E(n706), .CK(clk), .Q(
        \block[0][5] ) );
  EDFFXL \block_reg[3][5]  ( .D(block_next[5]), .E(n660), .CK(clk), .Q(
        \block[3][5] ) );
  EDFFXL \block_reg[2][5]  ( .D(block_next[5]), .E(n676), .CK(clk), .Q(
        \block[2][5] ) );
  EDFFXL \block_reg[6][16]  ( .D(block_next[16]), .E(n610), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFXL \block_reg[4][16]  ( .D(block_next[16]), .E(n641), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFXL \block_reg[3][16]  ( .D(block_next[16]), .E(n659), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFXL \block_reg[1][16]  ( .D(block_next[16]), .E(n690), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFXL \block_reg[0][16]  ( .D(block_next[16]), .E(n705), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFXL \block_reg[2][16]  ( .D(block_next[16]), .E(n675), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFXL \block_reg[6][1]  ( .D(block_next[1]), .E(n611), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFXL \block_reg[5][1]  ( .D(block_next[1]), .E(n624), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFXL \block_reg[4][1]  ( .D(block_next[1]), .E(n642), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFXL \block_reg[0][1]  ( .D(block_next[1]), .E(n706), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFXL \block_reg[3][1]  ( .D(block_next[1]), .E(n660), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFXL \block_reg[2][1]  ( .D(block_next[1]), .E(n676), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFXL \block_reg[6][18]  ( .D(block_next[18]), .E(n610), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFXL \block_reg[4][18]  ( .D(block_next[18]), .E(n641), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFXL \block_reg[3][18]  ( .D(block_next[18]), .E(n659), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFXL \block_reg[1][18]  ( .D(block_next[18]), .E(n690), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFXL \block_reg[0][18]  ( .D(block_next[18]), .E(n705), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFXL \block_reg[2][18]  ( .D(block_next[18]), .E(n675), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFXL \block_reg[6][21]  ( .D(block_next[21]), .E(n55), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFXL \block_reg[4][21]  ( .D(block_next[21]), .E(n641), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFXL \block_reg[3][21]  ( .D(block_next[21]), .E(n659), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFXL \block_reg[1][21]  ( .D(block_next[21]), .E(n690), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFXL \block_reg[0][21]  ( .D(block_next[21]), .E(n705), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFXL \block_reg[2][21]  ( .D(block_next[21]), .E(n675), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFXL \block_reg[5][0]  ( .D(block_next[0]), .E(n624), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFXL \block_reg[0][0]  ( .D(block_next[0]), .E(n706), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFXL \block_reg[4][0]  ( .D(block_next[0]), .E(n642), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFXL \block_reg[3][0]  ( .D(block_next[0]), .E(n660), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFXL \block_reg[7][0]  ( .D(block_next[0]), .E(n597), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFXL \block_reg[2][0]  ( .D(block_next[0]), .E(n676), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFXL \block_reg[6][0]  ( .D(block_next[0]), .E(n611), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFX4 \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n693), .CK(clk), .Q(
        n47) );
  EDFFX4 \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n662), .CK(clk), .Q(
        n46) );
  EDFFX4 \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n708), .CK(clk), .Q(
        n45) );
  EDFFX4 \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n678), .CK(clk), .Q(
        n44) );
  EDFFX4 \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n626), .CK(clk), 
        .QN(n43) );
  EDFFX4 \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n596), .CK(clk), 
        .QN(n42) );
  EDFFX4 \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n644), .CK(clk), 
        .QN(n41) );
  EDFFX4 \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n613), .CK(clk), 
        .QN(n40) );
  EDFFX4 \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n662), .CK(clk), .Q(
        n37) );
  EDFFX4 \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n693), .CK(clk), .Q(
        n36) );
  EDFFX4 \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n678), .CK(clk), .Q(
        n35) );
  EDFFX4 \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n708), .CK(clk), .Q(
        n34) );
  EDFFX4 \blocktag_reg[5][5]  ( .D(n72), .E(n626), .CK(clk), .QN(n33) );
  EDFFX4 \blocktag_reg[7][5]  ( .D(n72), .E(n596), .CK(clk), .QN(n32) );
  EDFFX4 \blocktag_reg[4][5]  ( .D(n72), .E(n644), .CK(clk), .QN(n31) );
  EDFFX4 \blocktag_reg[6][5]  ( .D(n72), .E(n613), .CK(clk), .QN(n30) );
  EDFFX4 \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(n596), .CK(clk), .Q(
        n29) );
  EDFFX4 \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n626), .CK(clk), .Q(
        n28) );
  EDFFX4 \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n613), .CK(clk), .Q(
        n27) );
  EDFFX4 \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n644), .CK(clk), .Q(
        n26) );
  EDFFX4 \blocktag_reg[1][14]  ( .D(n76), .E(n692), .CK(clk), .QN(n9) );
  EDFFX4 \blocktag_reg[3][14]  ( .D(n76), .E(n661), .CK(clk), .QN(n8) );
  EDFFX4 \blocktag_reg[0][14]  ( .D(n76), .E(n707), .CK(clk), .QN(n7) );
  EDFFX4 \blocktag_reg[2][14]  ( .D(n76), .E(n677), .CK(clk), .QN(n6) );
  MX4X2 U3 ( .A(\blocktag[0][24] ), .B(\blocktag[2][24] ), .C(
        \blocktag[1][24] ), .D(\blocktag[3][24] ), .S0(n753), .S1(n725), .Y(
        n850) );
  MX4X2 U4 ( .A(\blocktag[4][17] ), .B(\blocktag[6][17] ), .C(
        \blocktag[5][17] ), .D(\blocktag[7][17] ), .S0(n753), .S1(n726), .Y(
        n863) );
  MX4X2 U5 ( .A(\blocktag[0][17] ), .B(\blocktag[2][17] ), .C(
        \blocktag[1][17] ), .D(\blocktag[3][17] ), .S0(n753), .S1(n726), .Y(
        n864) );
  MX4X2 U6 ( .A(\blocktag[0][1] ), .B(\blocktag[2][1] ), .C(\blocktag[1][1] ), 
        .D(\blocktag[3][1] ), .S0(n753), .S1(n726), .Y(n866) );
  MX4X2 U7 ( .A(n66), .B(n77), .C(n62), .D(n71), .S0(n753), .S1(n726), .Y(n862) );
  MX4XL U8 ( .A(\block[4][119] ), .B(\block[6][119] ), .C(\block[5][119] ), 
        .D(\block[7][119] ), .S0(n749), .S1(n721), .Y(n1471) );
  MX4X2 U9 ( .A(\blocktag[0][19] ), .B(\blocktag[2][19] ), .C(
        \blocktag[1][19] ), .D(\blocktag[3][19] ), .S0(n441), .S1(n724), .Y(
        n874) );
  OAI221X4 U10 ( .A0(n1599), .A1(n505), .B0(n1598), .B1(n582), .C0(n1597), .Y(
        proc_rdata[9]) );
  MX4X4 U11 ( .A(\blocktag[5][0] ), .B(\blocktag[7][0] ), .C(\blocktag[4][0] ), 
        .D(\blocktag[6][0] ), .S0(n752), .S1(n738), .Y(n851) );
  MXI4X2 U12 ( .A(n50), .B(n51), .C(n48), .D(n49), .S0(n763), .S1(n726), .Y(
        n839) );
  MX4X4 U13 ( .A(n34), .B(n35), .C(n36), .D(n37), .S0(n751), .S1(n724), .Y(
        n820) );
  AO22X1 U14 ( .A0(proc_addr[15]), .A1(mem_read), .B0(mem_write), .B1(n414), 
        .Y(n1763) );
  XOR2X4 U15 ( .A(n2), .B(n1), .Y(n869) );
  CLKINVX20 U16 ( .A(n4), .Y(n1) );
  MX2XL U17 ( .A(n842), .B(n841), .S0(n779), .Y(n430) );
  AO22X2 U18 ( .A0(proc_addr[26]), .A1(mem_read), .B0(mem_write), .B1(n1535), 
        .Y(n1752) );
  CLKINVX8 U19 ( .A(n1752), .Y(n164) );
  CLKMX2X6 U20 ( .A(n811), .B(n812), .S0(n106), .Y(n1523) );
  INVX20 U21 ( .A(n786), .Y(n780) );
  MXI2X4 U22 ( .A(n810), .B(n809), .S0(n772), .Y(n85) );
  INVX20 U23 ( .A(n784), .Y(n772) );
  CLKMX2X6 U24 ( .A(n862), .B(n861), .S0(n772), .Y(n2) );
  CLKBUFX2 U25 ( .A(n1537), .Y(n3) );
  CLKINVX20 U26 ( .A(proc_addr[27]), .Y(n4) );
  CLKINVX6 U27 ( .A(n398), .Y(n5) );
  CLKINVX6 U28 ( .A(n779), .Y(n398) );
  MX4X4 U29 ( .A(\blocktag[0][4] ), .B(\blocktag[2][4] ), .C(\blocktag[1][4] ), 
        .D(\blocktag[3][4] ), .S0(n752), .S1(n724), .Y(n824) );
  CLKINVX1 U30 ( .A(n1526), .Y(n906) );
  MXI4X4 U31 ( .A(n6), .B(n7), .C(n8), .D(n9), .S0(n502), .S1(n723), .Y(n834)
         );
  CLKINVX1 U32 ( .A(n906), .Y(n10) );
  XOR2X4 U33 ( .A(n11), .B(n19), .Y(n815) );
  MXI2X4 U34 ( .A(n813), .B(n814), .S0(n783), .Y(n11) );
  INVX3 U35 ( .A(n761), .Y(n757) );
  CLKINVX1 U36 ( .A(n96), .Y(n12) );
  INVX3 U37 ( .A(n12), .Y(n13) );
  BUFX20 U38 ( .A(n1709), .Y(n96) );
  MX4X4 U39 ( .A(\blocktag[5][12] ), .B(\blocktag[7][12] ), .C(
        \blocktag[4][12] ), .D(\blocktag[6][12] ), .S0(n415), .S1(n740), .Y(
        n831) );
  INVX20 U40 ( .A(n739), .Y(n724) );
  CLKMX2X6 U41 ( .A(n833), .B(n834), .S0(n106), .Y(n1530) );
  CLKINVX12 U42 ( .A(n780), .Y(n106) );
  CLKINVX1 U43 ( .A(n927), .Y(n414) );
  MXI2X2 U44 ( .A(n927), .B(n926), .S0(n565), .Y(n75) );
  MX4X4 U45 ( .A(n410), .B(n411), .C(n412), .D(n413), .S0(n762), .S1(n724), 
        .Y(n400) );
  XOR2X4 U46 ( .A(n1533), .B(n14), .Y(n875) );
  CLKINVX20 U47 ( .A(n930), .Y(n14) );
  XOR2X4 U48 ( .A(n95), .B(n916), .Y(n879) );
  CLKINVX3 U49 ( .A(proc_addr[18]), .Y(n916) );
  OR2X8 U50 ( .A(n1549), .B(n15), .Y(n541) );
  AND3X8 U51 ( .A(n1547), .B(n1546), .C(n523), .Y(n93) );
  AND3X6 U52 ( .A(n1546), .B(n1547), .C(n534), .Y(n521) );
  OR2X8 U53 ( .A(n1549), .B(n20), .Y(n97) );
  OR2X1 U54 ( .A(n394), .B(n1539), .Y(n15) );
  MX4X4 U55 ( .A(n87), .B(n89), .C(n88), .D(n90), .S0(n724), .S1(n532), .Y(
        n809) );
  INVX3 U56 ( .A(proc_addr[0]), .Y(n394) );
  CLKMX2X3 U57 ( .A(n810), .B(n809), .S0(n780), .Y(n437) );
  INVX3 U58 ( .A(n21), .Y(n22) );
  INVX1 U59 ( .A(n97), .Y(n539) );
  CLKINVX1 U60 ( .A(n1547), .Y(n21) );
  MXI2X4 U61 ( .A(n16), .B(n17), .S0(n781), .Y(n1536) );
  MX4X2 U62 ( .A(n465), .B(n466), .C(n463), .D(n464), .S0(n442), .S1(n738), 
        .Y(n16) );
  MX4X1 U63 ( .A(n506), .B(n507), .C(n508), .D(n509), .S0(n415), .S1(n725), 
        .Y(n17) );
  INVX20 U64 ( .A(n786), .Y(n779) );
  CLKBUFX8 U65 ( .A(n786), .Y(n781) );
  MX2XL U66 ( .A(n813), .B(n814), .S0(n783), .Y(n18) );
  CLKINVX20 U67 ( .A(n893), .Y(n19) );
  BUFX20 U68 ( .A(n743), .Y(n740) );
  NAND2X4 U69 ( .A(n958), .B(proc_stall), .Y(n883) );
  CLKINVX12 U70 ( .A(n948), .Y(proc_stall) );
  AOI2BB1X4 U71 ( .A0N(n948), .A1N(n965), .B0(n947), .Y(n949) );
  NAND2X8 U72 ( .A(n960), .B(n966), .Y(n948) );
  INVX20 U73 ( .A(n764), .Y(n415) );
  MX4X2 U74 ( .A(\blocktag[4][21] ), .B(\blocktag[6][21] ), .C(
        \blocktag[5][21] ), .D(\blocktag[7][21] ), .S0(n752), .S1(n726), .Y(
        n853) );
  MX2X6 U75 ( .A(n874), .B(n873), .S0(n779), .Y(n1533) );
  NAND3X8 U76 ( .A(n93), .B(n1548), .C(n92), .Y(n91) );
  CLKINVX20 U77 ( .A(n742), .Y(n713) );
  BUFX20 U78 ( .A(n744), .Y(n742) );
  OR2XL U79 ( .A(n394), .B(n1539), .Y(n20) );
  INVX16 U80 ( .A(n1541), .Y(n1546) );
  NAND2X4 U81 ( .A(n1518), .B(n1520), .Y(n1519) );
  OAI22X2 U82 ( .A0(n796), .A1(n960), .B0(n959), .B1(n958), .Y(n67) );
  MXI4X2 U83 ( .A(n535), .B(n536), .C(n537), .D(n538), .S0(n768), .S1(n726), 
        .Y(n865) );
  CLKAND2X3 U84 ( .A(n1519), .B(n760), .Y(n1774) );
  MX4XL U85 ( .A(\block[0][117] ), .B(\block[2][117] ), .C(\block[1][117] ), 
        .D(\block[3][117] ), .S0(n760), .S1(n721), .Y(n1462) );
  MX4X1 U86 ( .A(\block[4][30] ), .B(\block[6][30] ), .C(\block[5][30] ), .D(
        \block[7][30] ), .S0(n757), .S1(n731), .Y(n1085) );
  MX4X1 U87 ( .A(\block[4][31] ), .B(\block[6][31] ), .C(\block[5][31] ), .D(
        \block[7][31] ), .S0(n757), .S1(n731), .Y(n1089) );
  MX4X1 U88 ( .A(\block[4][29] ), .B(\block[6][29] ), .C(\block[5][29] ), .D(
        \block[7][29] ), .S0(n757), .S1(n731), .Y(n1081) );
  MX4X1 U89 ( .A(\block[0][29] ), .B(\block[2][29] ), .C(\block[1][29] ), .D(
        \block[3][29] ), .S0(n757), .S1(n731), .Y(n1082) );
  MX4X1 U90 ( .A(\block[0][30] ), .B(\block[2][30] ), .C(\block[1][30] ), .D(
        \block[3][30] ), .S0(n757), .S1(n731), .Y(n1086) );
  MX4X1 U91 ( .A(\block[0][28] ), .B(\block[2][28] ), .C(\block[1][28] ), .D(
        \block[3][28] ), .S0(n757), .S1(n731), .Y(n1078) );
  MX4X1 U92 ( .A(\block[4][27] ), .B(\block[6][27] ), .C(\block[5][27] ), .D(
        \block[7][27] ), .S0(n757), .S1(n731), .Y(n1073) );
  MX4X1 U93 ( .A(\block[4][28] ), .B(\block[6][28] ), .C(\block[5][28] ), .D(
        \block[7][28] ), .S0(n757), .S1(n731), .Y(n1077) );
  MX4XL U94 ( .A(\block[0][106] ), .B(\block[2][106] ), .C(\block[1][106] ), 
        .D(\block[3][106] ), .S0(n748), .S1(n719), .Y(n1407) );
  MX4XL U95 ( .A(\block[4][104] ), .B(\block[6][104] ), .C(\block[5][104] ), 
        .D(\block[7][104] ), .S0(n748), .S1(n719), .Y(n1396) );
  MX4XL U96 ( .A(\block[4][115] ), .B(\block[6][115] ), .C(\block[5][115] ), 
        .D(\block[7][115] ), .S0(n748), .S1(n721), .Y(n1451) );
  MX4XL U97 ( .A(\block[4][106] ), .B(\block[6][106] ), .C(\block[5][106] ), 
        .D(\block[7][106] ), .S0(n542), .S1(n719), .Y(n1406) );
  MX4XL U98 ( .A(\block[4][105] ), .B(\block[6][105] ), .C(\block[5][105] ), 
        .D(\block[7][105] ), .S0(n542), .S1(n719), .Y(n1401) );
  MX4XL U99 ( .A(\block[0][110] ), .B(\block[2][110] ), .C(\block[1][110] ), 
        .D(\block[3][110] ), .S0(n542), .S1(n720), .Y(n1427) );
  MX4XL U100 ( .A(\block[4][110] ), .B(\block[6][110] ), .C(\block[5][110] ), 
        .D(\block[7][110] ), .S0(n542), .S1(n720), .Y(n1426) );
  MX4XL U101 ( .A(\block[4][113] ), .B(\block[6][113] ), .C(\block[5][113] ), 
        .D(\block[7][113] ), .S0(n542), .S1(n720), .Y(n1441) );
  MX4XL U102 ( .A(\block[4][109] ), .B(\block[6][109] ), .C(\block[5][109] ), 
        .D(\block[7][109] ), .S0(n542), .S1(n720), .Y(n1421) );
  MX4XL U103 ( .A(\block[0][115] ), .B(\block[2][115] ), .C(\block[1][115] ), 
        .D(\block[3][115] ), .S0(n542), .S1(n720), .Y(n1452) );
  MX4X1 U104 ( .A(\block[4][61] ), .B(\block[6][61] ), .C(\block[5][61] ), .D(
        \block[7][61] ), .S0(n749), .S1(n713), .Y(n1210) );
  MX4XL U105 ( .A(\block[0][105] ), .B(\block[2][105] ), .C(\block[1][105] ), 
        .D(\block[3][105] ), .S0(n749), .S1(n719), .Y(n1402) );
  MX4XL U106 ( .A(\block[0][108] ), .B(\block[2][108] ), .C(\block[1][108] ), 
        .D(\block[3][108] ), .S0(n749), .S1(n719), .Y(n1417) );
  MX4XL U107 ( .A(\block[4][108] ), .B(\block[6][108] ), .C(\block[5][108] ), 
        .D(\block[7][108] ), .S0(n103), .S1(n719), .Y(n1416) );
  MX4XL U108 ( .A(\block[4][112] ), .B(\block[6][112] ), .C(\block[5][112] ), 
        .D(\block[7][112] ), .S0(n103), .S1(n720), .Y(n1436) );
  MX4XL U109 ( .A(\block[0][114] ), .B(\block[2][114] ), .C(\block[1][114] ), 
        .D(\block[3][114] ), .S0(n103), .S1(n720), .Y(n1447) );
  XOR2X4 U110 ( .A(n1536), .B(n23), .Y(n857) );
  CLKINVX20 U111 ( .A(proc_addr[28]), .Y(n23) );
  INVX8 U112 ( .A(n765), .Y(n103) );
  INVX16 U113 ( .A(n404), .Y(n758) );
  CLKBUFX2 U114 ( .A(n1524), .Y(n24) );
  BUFX8 U115 ( .A(n1522), .Y(n25) );
  INVX2 U116 ( .A(proc_addr[28]), .Y(n945) );
  MX4X4 U117 ( .A(n26), .B(n27), .C(n28), .D(n29), .S0(n439), .S1(n723), .Y(
        n821) );
  MXI4X4 U118 ( .A(n30), .B(n31), .C(n32), .D(n33), .S0(n763), .S1(n725), .Y(
        n813) );
  INVX8 U119 ( .A(n739), .Y(n725) );
  MX4X4 U120 ( .A(\blocktag[0][7] ), .B(\blocktag[2][7] ), .C(\blocktag[1][7] ), .D(\blocktag[3][7] ), .S0(n752), .S1(n724), .Y(n840) );
  XOR2X4 U121 ( .A(n1530), .B(n38), .Y(n835) );
  CLKINVX20 U122 ( .A(n39), .Y(n38) );
  CLKINVX20 U123 ( .A(n914), .Y(n39) );
  MXI4X4 U124 ( .A(n40), .B(n41), .C(n42), .D(n43), .S0(n761), .S1(n725), .Y(
        n837) );
  CLKINVX20 U125 ( .A(n771), .Y(n786) );
  MX4X2 U126 ( .A(n44), .B(n45), .C(n46), .D(n47), .S0(n502), .S1(n724), .Y(
        n812) );
  NAND4X8 U127 ( .A(n818), .B(n816), .C(n815), .D(n817), .Y(n828) );
  BUFX12 U128 ( .A(proc_read), .Y(n793) );
  CLKINVX4 U129 ( .A(n526), .Y(n524) );
  CLKINVX1 U130 ( .A(n891), .Y(n526) );
  INVX2 U131 ( .A(n533), .Y(n92) );
  INVX4 U132 ( .A(n1539), .Y(n1548) );
  NOR2X2 U133 ( .A(n1542), .B(n1539), .Y(n534) );
  MX4X1 U134 ( .A(\block[4][93] ), .B(\block[6][93] ), .C(\block[5][93] ), .D(
        \block[7][93] ), .S0(n103), .S1(n734), .Y(n1339) );
  MX4X1 U135 ( .A(\block[0][93] ), .B(\block[2][93] ), .C(\block[1][93] ), .D(
        \block[3][93] ), .S0(n542), .S1(n734), .Y(n1340) );
  MX4XL U136 ( .A(\block[0][124] ), .B(\block[2][124] ), .C(\block[1][124] ), 
        .D(\block[3][124] ), .S0(n750), .S1(n722), .Y(n1497) );
  BUFX20 U137 ( .A(n1748), .Y(mem_read) );
  CLKINVX3 U138 ( .A(n779), .Y(n86) );
  CLKINVX1 U139 ( .A(n397), .Y(n396) );
  CLKINVX1 U140 ( .A(n905), .Y(n446) );
  INVX3 U141 ( .A(n519), .Y(n403) );
  CLKINVX1 U142 ( .A(n902), .Y(n519) );
  CLKINVX1 U143 ( .A(n895), .Y(n514) );
  CLKINVX2 U144 ( .A(n780), .Y(n107) );
  CLKINVX1 U145 ( .A(n780), .Y(n435) );
  CLKINVX1 U146 ( .A(n919), .Y(n94) );
  INVX1 U147 ( .A(n933), .Y(n445) );
  INVX12 U148 ( .A(n793), .Y(n796) );
  MX4X1 U149 ( .A(blockdirty[0]), .B(blockdirty[2]), .C(blockdirty[1]), .D(
        blockdirty[3]), .S0(n748), .S1(n734), .Y(n807) );
  MX4XL U150 ( .A(\block[4][5] ), .B(\block[6][5] ), .C(\block[5][5] ), .D(
        \block[7][5] ), .S0(n444), .S1(n727), .Y(n985) );
  MX4XL U151 ( .A(\block[0][5] ), .B(\block[2][5] ), .C(\block[1][5] ), .D(
        \block[3][5] ), .S0(n754), .S1(n727), .Y(n986) );
  MX4XL U152 ( .A(\block[0][7] ), .B(\block[2][7] ), .C(\block[1][7] ), .D(
        \block[3][7] ), .S0(n755), .S1(n727), .Y(n994) );
  MX4XL U153 ( .A(\block[4][33] ), .B(\block[6][33] ), .C(\block[5][33] ), .D(
        \block[7][33] ), .S0(n758), .S1(n732), .Y(n1098) );
  MX4XL U154 ( .A(\block[0][34] ), .B(\block[2][34] ), .C(\block[1][34] ), .D(
        \block[3][34] ), .S0(n758), .S1(n732), .Y(n1103) );
  MX4XL U155 ( .A(\block[0][35] ), .B(\block[2][35] ), .C(\block[1][35] ), .D(
        \block[3][35] ), .S0(n758), .S1(n732), .Y(n1107) );
  MX4XL U156 ( .A(\block[4][37] ), .B(\block[6][37] ), .C(\block[5][37] ), .D(
        \block[7][37] ), .S0(n758), .S1(n732), .Y(n1114) );
  MX4XL U157 ( .A(\block[4][39] ), .B(\block[6][39] ), .C(\block[5][39] ), .D(
        \block[7][39] ), .S0(n759), .S1(n733), .Y(n1122) );
  MX4XL U158 ( .A(\block[0][42] ), .B(\block[2][42] ), .C(\block[1][42] ), .D(
        \block[3][42] ), .S0(n759), .S1(n733), .Y(n1135) );
  MX4XL U159 ( .A(\block[0][43] ), .B(\block[2][43] ), .C(\block[1][43] ), .D(
        \block[3][43] ), .S0(n759), .S1(n733), .Y(n1139) );
  MX4X1 U160 ( .A(\block[0][46] ), .B(\block[2][46] ), .C(\block[1][46] ), .D(
        \block[3][46] ), .S0(n760), .S1(n734), .Y(n1151) );
  MX4X1 U161 ( .A(\block[0][47] ), .B(\block[2][47] ), .C(\block[1][47] ), .D(
        \block[3][47] ), .S0(n760), .S1(n734), .Y(n1155) );
  MX4XL U162 ( .A(\block[4][69] ), .B(\block[6][69] ), .C(\block[5][69] ), .D(
        \block[7][69] ), .S0(n754), .S1(n714), .Y(n1243) );
  MX4XL U163 ( .A(\block[0][71] ), .B(\block[2][71] ), .C(\block[1][71] ), .D(
        \block[3][71] ), .S0(n754), .S1(n714), .Y(n1252) );
  MX4XL U164 ( .A(\block[0][74] ), .B(\block[2][74] ), .C(\block[1][74] ), .D(
        \block[3][74] ), .S0(n754), .S1(n715), .Y(n1264) );
  MX4XL U165 ( .A(\block[0][75] ), .B(\block[2][75] ), .C(\block[1][75] ), .D(
        \block[3][75] ), .S0(n749), .S1(n715), .Y(n1268) );
  MX4XL U166 ( .A(\block[0][78] ), .B(\block[2][78] ), .C(\block[1][78] ), .D(
        \block[3][78] ), .S0(n754), .S1(n715), .Y(n1280) );
  MX4XL U167 ( .A(\block[0][79] ), .B(\block[2][79] ), .C(\block[1][79] ), .D(
        \block[3][79] ), .S0(n754), .S1(n715), .Y(n1284) );
  MX4XL U168 ( .A(\block[0][94] ), .B(\block[2][94] ), .C(\block[1][94] ), .D(
        \block[3][94] ), .S0(n103), .S1(n734), .Y(n1344) );
  MX4XL U169 ( .A(\block[4][94] ), .B(\block[6][94] ), .C(\block[5][94] ), .D(
        \block[7][94] ), .S0(n542), .S1(n734), .Y(n1343) );
  MX4XL U170 ( .A(\block[4][98] ), .B(\block[6][98] ), .C(\block[5][98] ), .D(
        \block[7][98] ), .S0(n758), .S1(n718), .Y(n1366) );
  MX4XL U171 ( .A(\block[0][99] ), .B(\block[2][99] ), .C(\block[1][99] ), .D(
        \block[3][99] ), .S0(n747), .S1(n718), .Y(n1372) );
  MX4XL U172 ( .A(\block[4][101] ), .B(\block[6][101] ), .C(\block[5][101] ), 
        .D(\block[7][101] ), .S0(n747), .S1(n718), .Y(n1381) );
  MX4XL U173 ( .A(\block[4][103] ), .B(\block[6][103] ), .C(\block[5][103] ), 
        .D(\block[7][103] ), .S0(n747), .S1(n719), .Y(n1391) );
  MX4XL U174 ( .A(\block[0][107] ), .B(\block[2][107] ), .C(\block[1][107] ), 
        .D(\block[3][107] ), .S0(n748), .S1(n719), .Y(n1412) );
  MX4XL U175 ( .A(\block[0][111] ), .B(\block[2][111] ), .C(\block[1][111] ), 
        .D(\block[3][111] ), .S0(n542), .S1(n720), .Y(n1432) );
  MX4X1 U176 ( .A(\block[4][123] ), .B(\block[6][123] ), .C(\block[5][123] ), 
        .D(\block[7][123] ), .S0(n750), .S1(n722), .Y(n1491) );
  MX4X1 U177 ( .A(\block[0][123] ), .B(\block[2][123] ), .C(\block[1][123] ), 
        .D(\block[3][123] ), .S0(n750), .S1(n722), .Y(n1492) );
  MX4XL U178 ( .A(\block[0][126] ), .B(\block[2][126] ), .C(\block[1][126] ), 
        .D(\block[3][126] ), .S0(n750), .S1(n722), .Y(n1505) );
  MX4XL U179 ( .A(\block[4][126] ), .B(\block[6][126] ), .C(\block[5][126] ), 
        .D(\block[7][126] ), .S0(n750), .S1(n722), .Y(n1504) );
  CLKMX2X2 U180 ( .A(n1510), .B(n1509), .S0(n772), .Y(n1516) );
  NOR2X2 U181 ( .A(n100), .B(n945), .Y(n102) );
  MX2X2 U182 ( .A(n822), .B(n821), .S0(n780), .Y(n1525) );
  MX4X2 U183 ( .A(\blocktag[0][21] ), .B(\blocktag[2][21] ), .C(
        \blocktag[1][21] ), .D(\blocktag[3][21] ), .S0(n751), .S1(n438), .Y(
        n854) );
  INVX3 U184 ( .A(n1346), .Y(n1700) );
  BUFX4 U185 ( .A(n55), .Y(n601) );
  CLKINVX6 U186 ( .A(n1776), .Y(n390) );
  INVXL U187 ( .A(n527), .Y(n1503) );
  CLKBUFX12 U188 ( .A(n1751), .Y(mem_addr[25]) );
  CLKINVX1 U189 ( .A(n458), .Y(n920) );
  MXI2X4 U190 ( .A(n915), .B(n914), .S0(n558), .Y(n76) );
  CLKINVX1 U191 ( .A(n429), .Y(n915) );
  CLKAND2X12 U192 ( .A(n58), .B(n794), .Y(n52) );
  AND2X8 U193 ( .A(n57), .B(n794), .Y(n53) );
  AND2X4 U194 ( .A(n952), .B(n794), .Y(n54) );
  AND2X8 U195 ( .A(n953), .B(n794), .Y(n55) );
  BUFX16 U196 ( .A(n1511), .Y(n559) );
  BUFX16 U197 ( .A(n559), .Y(n569) );
  CLKINVX12 U198 ( .A(N31), .Y(n745) );
  BUFX16 U199 ( .A(n745), .Y(n739) );
  BUFX12 U200 ( .A(n745), .Y(n744) );
  CLKAND2X12 U201 ( .A(n60), .B(n794), .Y(n56) );
  AND2X2 U202 ( .A(n1744), .B(n735), .Y(n57) );
  AND2X2 U203 ( .A(n1745), .B(n737), .Y(n58) );
  INVX12 U204 ( .A(proc_addr[1]), .Y(n533) );
  AND2X1 U205 ( .A(n1746), .B(n738), .Y(n59) );
  AND2X1 U206 ( .A(n1747), .B(n734), .Y(n60) );
  AND2X6 U207 ( .A(n59), .B(n794), .Y(n61) );
  CLKBUFX3 U208 ( .A(n52), .Y(n666) );
  AND2X1 U209 ( .A(n1746), .B(n734), .Y(n63) );
  AND2X8 U210 ( .A(n63), .B(n794), .Y(n64) );
  AND2X2 U211 ( .A(n395), .B(n575), .Y(n65) );
  CLKINVX3 U212 ( .A(n555), .Y(n553) );
  CLKINVX3 U213 ( .A(n555), .Y(n554) );
  BUFX8 U214 ( .A(n739), .Y(n741) );
  BUFX16 U215 ( .A(n743), .Y(n738) );
  BUFX4 U216 ( .A(n743), .Y(n737) );
  BUFX16 U217 ( .A(n1749), .Y(n787) );
  MXI2X8 U218 ( .A(n920), .B(n919), .S0(n571), .Y(n68) );
  MXI2X8 U219 ( .A(n98), .B(n945), .S0(n572), .Y(n69) );
  AND2X6 U220 ( .A(n79), .B(n551), .Y(n70) );
  INVX16 U221 ( .A(n766), .Y(n747) );
  CLKBUFX3 U222 ( .A(n1711), .Y(n710) );
  CLKINVX1 U223 ( .A(n407), .Y(n408) );
  INVX1 U224 ( .A(proc_reset), .Y(n795) );
  BUFX6 U225 ( .A(n795), .Y(n794) );
  MXI2X4 U226 ( .A(n894), .B(n893), .S0(n560), .Y(n72) );
  MXI2X4 U227 ( .A(n925), .B(n924), .S0(n565), .Y(n73) );
  MXI2X4 U228 ( .A(n912), .B(n911), .S0(n572), .Y(n74) );
  INVX6 U229 ( .A(n504), .Y(n505) );
  CLKAND2X12 U230 ( .A(n533), .B(n1545), .Y(n78) );
  AND2X4 U231 ( .A(n65), .B(n557), .Y(n79) );
  INVXL U232 ( .A(proc_addr[16]), .Y(n908) );
  INVX3 U233 ( .A(n961), .Y(n1543) );
  CLKINVX1 U234 ( .A(mem_ready), .Y(n965) );
  CLKINVX3 U235 ( .A(proc_addr[14]), .Y(n104) );
  OR2X8 U236 ( .A(n101), .B(n102), .Y(n80) );
  CLKINVX4 U237 ( .A(proc_addr[21]), .Y(n397) );
  CLKINVX1 U238 ( .A(n1536), .Y(n98) );
  CLKBUFX3 U239 ( .A(n54), .Y(n650) );
  CLKBUFX3 U240 ( .A(n53), .Y(n681) );
  INVX1 U241 ( .A(n1355), .Y(n555) );
  NAND2X1 U242 ( .A(mem_rdata[63]), .B(n1511), .Y(n1220) );
  NAND2XL U243 ( .A(mem_rdata[66]), .B(n1511), .Y(n1233) );
  NAND2XL U244 ( .A(mem_rdata[84]), .B(n1511), .Y(n1305) );
  NAND2XL U245 ( .A(mem_rdata[7]), .B(n1511), .Y(n995) );
  NAND2XL U246 ( .A(mem_rdata[40]), .B(n1511), .Y(n1128) );
  MX2X1 U247 ( .A(n909), .B(n908), .S0(n1511), .Y(n910) );
  MX2X1 U248 ( .A(n424), .B(n397), .S0(n1511), .Y(n913) );
  NAND2X6 U249 ( .A(n79), .B(n553), .Y(n963) );
  CLKINVX12 U250 ( .A(n963), .Y(n1092) );
  OAI221X4 U251 ( .A0(n1389), .A1(n551), .B0(n1584), .B1(n545), .C0(n991), .Y(
        block_next[6]) );
  BUFX20 U252 ( .A(n1092), .Y(n545) );
  BUFX12 U253 ( .A(n1511), .Y(n558) );
  NAND2X2 U254 ( .A(mem_ready), .B(n1517), .Y(n808) );
  NAND2X8 U255 ( .A(n959), .B(n447), .Y(n960) );
  INVX6 U256 ( .A(n967), .Y(n959) );
  OAI221X4 U257 ( .A0(n1656), .A1(n550), .B0(n1464), .B1(n556), .C0(n1309), 
        .Y(block_next[85]) );
  INVX3 U258 ( .A(n808), .Y(n958) );
  OAI221X4 U259 ( .A0(n1359), .A1(n551), .B0(n1554), .B1(n545), .C0(n964), .Y(
        block_next[0]) );
  OAI221X4 U260 ( .A0(n1646), .A1(n550), .B0(n1454), .B1(n557), .C0(n1301), 
        .Y(block_next[83]) );
  OAI221X4 U261 ( .A0(n1464), .A1(n551), .B0(n1659), .B1(n1092), .C0(n1051), 
        .Y(block_next[21]) );
  OAI221X4 U262 ( .A0(n1661), .A1(n550), .B0(n1469), .B1(n556), .C0(n1313), 
        .Y(block_next[86]) );
  OAI221X4 U263 ( .A0(n1626), .A1(n550), .B0(n1434), .B1(n556), .C0(n1285), 
        .Y(block_next[79]) );
  OAI221X4 U264 ( .A0(n1449), .A1(n552), .B0(n1644), .B1(n1092), .C0(n1039), 
        .Y(block_next[18]) );
  OAI221X4 U265 ( .A0(n1364), .A1(n551), .B0(n1559), .B1(n545), .C0(n971), .Y(
        block_next[1]) );
  OAI221X4 U266 ( .A0(n1621), .A1(n550), .B0(n1429), .B1(n556), .C0(n1281), 
        .Y(block_next[78]) );
  OAI221X4 U267 ( .A0(n1676), .A1(n550), .B0(n1484), .B1(n557), .C0(n1325), 
        .Y(block_next[89]) );
  OAI221X4 U268 ( .A0(n1671), .A1(n550), .B0(n1479), .B1(n556), .C0(n1321), 
        .Y(block_next[88]) );
  OAI221X4 U269 ( .A0(n1439), .A1(n552), .B0(n1634), .B1(n1092), .C0(n1031), 
        .Y(block_next[16]) );
  OAI221X4 U270 ( .A0(n1384), .A1(n551), .B0(n1579), .B1(n545), .C0(n987), .Y(
        block_next[5]) );
  OAI221X4 U271 ( .A0(n1651), .A1(n550), .B0(n1459), .B1(n556), .C0(n1305), 
        .Y(block_next[84]) );
  OAI221X4 U272 ( .A0(n1636), .A1(n550), .B0(n1444), .B1(n556), .C0(n1293), 
        .Y(block_next[81]) );
  OAI221X4 U273 ( .A0(n1631), .A1(n550), .B0(n1439), .B1(n556), .C0(n1289), 
        .Y(block_next[80]) );
  OAI221X4 U274 ( .A0(n1429), .A1(n552), .B0(n1624), .B1(n1092), .C0(n1023), 
        .Y(block_next[14]) );
  OAI221X4 U275 ( .A0(n1404), .A1(n552), .B0(n1599), .B1(n545), .C0(n1003), 
        .Y(block_next[9]) );
  OAI221X4 U276 ( .A0(n1434), .A1(n552), .B0(n1629), .B1(n1092), .C0(n1027), 
        .Y(block_next[15]) );
  OAI221X4 U277 ( .A0(n1379), .A1(n551), .B0(n1574), .B1(n545), .C0(n983), .Y(
        block_next[4]) );
  OAI221X4 U278 ( .A0(n1444), .A1(n552), .B0(n1639), .B1(n1092), .C0(n1035), 
        .Y(block_next[17]) );
  OAI221X4 U279 ( .A0(n1369), .A1(n551), .B0(n1564), .B1(n545), .C0(n975), .Y(
        block_next[2]) );
  OAI221X4 U280 ( .A0(n1419), .A1(n552), .B0(n1614), .B1(n1092), .C0(n1015), 
        .Y(block_next[12]) );
  OAI221X4 U281 ( .A0(n1399), .A1(n552), .B0(n1594), .B1(n545), .C0(n999), .Y(
        block_next[8]) );
  OAI221X4 U282 ( .A0(n1691), .A1(n549), .B0(n1499), .B1(n557), .C0(n1337), 
        .Y(block_next[92]) );
  OAI221X4 U283 ( .A0(n1666), .A1(n550), .B0(n1474), .B1(n557), .C0(n1317), 
        .Y(block_next[87]) );
  BUFX12 U284 ( .A(n1350), .Y(n550) );
  OAI221X4 U285 ( .A0(n1681), .A1(n550), .B0(n1489), .B1(n556), .C0(n1329), 
        .Y(block_next[90]) );
  OAI221X4 U286 ( .A0(n1641), .A1(n550), .B0(n1449), .B1(n556), .C0(n1297), 
        .Y(block_next[82]) );
  OAI221X4 U287 ( .A0(n1424), .A1(n552), .B0(n1619), .B1(n1092), .C0(n1019), 
        .Y(block_next[13]) );
  OAI221X4 U288 ( .A0(n1374), .A1(n552), .B0(n1569), .B1(n545), .C0(n979), .Y(
        block_next[3]) );
  OAI221X4 U289 ( .A0(n1616), .A1(n550), .B0(n1424), .B1(n556), .C0(n1277), 
        .Y(block_next[77]) );
  OAI221X4 U290 ( .A0(n1454), .A1(n551), .B0(n1649), .B1(n1092), .C0(n1043), 
        .Y(block_next[19]) );
  OAI221X4 U291 ( .A0(n1409), .A1(n552), .B0(n1604), .B1(n545), .C0(n1007), 
        .Y(block_next[10]) );
  OAI221X4 U292 ( .A0(n1474), .A1(n551), .B0(n1669), .B1(n1092), .C0(n1059), 
        .Y(block_next[23]) );
  OAI221X4 U293 ( .A0(n1414), .A1(n552), .B0(n1609), .B1(n545), .C0(n1011), 
        .Y(block_next[11]) );
  OAI221X4 U294 ( .A0(n1469), .A1(n551), .B0(n1664), .B1(n1092), .C0(n1055), 
        .Y(block_next[22]) );
  OAI221X4 U295 ( .A0(n1394), .A1(n552), .B0(n1589), .B1(n545), .C0(n995), .Y(
        block_next[7]) );
  BUFX16 U296 ( .A(n768), .Y(n766) );
  CLKINVX8 U297 ( .A(n765), .Y(n542) );
  CLKINVX6 U298 ( .A(n765), .Y(n749) );
  INVX8 U299 ( .A(n765), .Y(n441) );
  INVX8 U300 ( .A(n532), .Y(n442) );
  MX4X4 U301 ( .A(n81), .B(n82), .C(n83), .D(n84), .S0(n415), .S1(n724), .Y(
        n829) );
  XNOR2X4 U302 ( .A(n85), .B(n888), .Y(n817) );
  MX4X4 U303 ( .A(\blocktag[0][16] ), .B(\blocktag[2][16] ), .C(
        \blocktag[1][16] ), .D(\blocktag[3][16] ), .S0(n751), .S1(n724), .Y(
        n830) );
  MXI4X4 U304 ( .A(n517), .B(n518), .C(n515), .D(n516), .S0(n761), .S1(n725), 
        .Y(n822) );
  MXI2X4 U305 ( .A(n829), .B(n830), .S0(n86), .Y(n419) );
  CLKMX2X2 U306 ( .A(n805), .B(n804), .S0(n780), .Y(n418) );
  MX4X4 U307 ( .A(\blocktag[3][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[0][18] ), .S0(n768), .S1(n744), .Y(
        n810) );
  CLKMX2X6 U308 ( .A(n824), .B(n823), .S0(n779), .Y(n1524) );
  NAND3X6 U309 ( .A(n93), .B(n1548), .C(n92), .Y(n1705) );
  CLKINVX1 U310 ( .A(n894), .Y(n436) );
  AO22X1 U311 ( .A0(proc_addr[10]), .A1(mem_read), .B0(mem_write), .B1(n436), 
        .Y(n1768) );
  XOR2X4 U312 ( .A(n1531), .B(n94), .Y(n880) );
  CLKMX2X6 U313 ( .A(n854), .B(n853), .S0(n779), .Y(n1535) );
  MXI2X4 U314 ( .A(n878), .B(n877), .S0(n779), .Y(n95) );
  INVX16 U315 ( .A(n766), .Y(n746) );
  INVX4 U316 ( .A(n883), .Y(n1511) );
  BUFX20 U317 ( .A(n558), .Y(n571) );
  BUFX20 U318 ( .A(n558), .Y(n568) );
  BUFX16 U319 ( .A(n559), .Y(n570) );
  BUFX20 U320 ( .A(n558), .Y(n566) );
  BUFX20 U321 ( .A(n570), .Y(n563) );
  BUFX20 U322 ( .A(n571), .Y(n562) );
  BUFX20 U323 ( .A(n572), .Y(n561) );
  BUFX20 U324 ( .A(n558), .Y(n567) );
  BUFX20 U325 ( .A(n569), .Y(n565) );
  BUFX20 U326 ( .A(n570), .Y(n564) );
  CLKINVX1 U327 ( .A(mem_write), .Y(n99) );
  INVX3 U328 ( .A(mem_read), .Y(n100) );
  NOR2X4 U329 ( .A(n98), .B(n99), .Y(n101) );
  CLKBUFX12 U330 ( .A(n767), .Y(n765) );
  XOR2X4 U331 ( .A(n402), .B(n104), .Y(n827) );
  CLKBUFX2 U332 ( .A(n10), .Y(n105) );
  CLKMX2X6 U333 ( .A(n832), .B(n831), .S0(n779), .Y(n1529) );
  BUFX20 U334 ( .A(n572), .Y(n560) );
  BUFX20 U335 ( .A(n559), .Y(n572) );
  MXI4X4 U336 ( .A(n114), .B(n115), .C(n116), .D(n117), .S0(n764), .S1(n744), 
        .Y(n811) );
  AND4X8 U337 ( .A(n869), .B(n867), .C(n868), .D(n870), .Y(n531) );
  INVX20 U338 ( .A(n502), .Y(n751) );
  MXI2X4 U339 ( .A(n819), .B(n820), .S0(n107), .Y(n402) );
  INVX1 U340 ( .A(n13), .Y(n504) );
  NAND2X2 U341 ( .A(mem_rdata[35]), .B(n570), .Y(n1108) );
  CLKINVX3 U342 ( .A(n1518), .Y(n1749) );
  OAI221X4 U343 ( .A0(n1679), .A1(n505), .B0(n1678), .B1(n520), .C0(n1677), 
        .Y(proc_rdata[25]) );
  OAI221X4 U344 ( .A0(n1674), .A1(n505), .B0(n1673), .B1(n520), .C0(n1672), 
        .Y(proc_rdata[24]) );
  MXI4X4 U345 ( .A(n108), .B(n109), .C(n110), .D(n111), .S0(n764), .S1(n723), 
        .Y(n814) );
  INVX16 U346 ( .A(n744), .Y(n723) );
  AO22XL U347 ( .A0(proc_addr[5]), .A1(mem_read), .B0(mem_write), .B1(n1521), 
        .Y(n1773) );
  INVX8 U348 ( .A(n1773), .Y(n122) );
  CLKMX2X6 U349 ( .A(n850), .B(n849), .S0(n779), .Y(n1537) );
  CLKBUFX2 U350 ( .A(n25), .Y(n112) );
  MX2X4 U351 ( .A(n878), .B(n877), .S0(n779), .Y(n113) );
  BUFX20 U352 ( .A(n769), .Y(n502) );
  INVX6 U353 ( .A(n768), .Y(n439) );
  INVX4 U354 ( .A(n766), .Y(n756) );
  INVX8 U355 ( .A(n532), .Y(n760) );
  CLKINVX20 U356 ( .A(n409), .Y(n759) );
  CLKMX2X6 U357 ( .A(n866), .B(n865), .S0(n779), .Y(n1522) );
  OAI221X4 U358 ( .A0(n1629), .A1(n505), .B0(n1628), .B1(n583), .C0(n1627), 
        .Y(proc_rdata[15]) );
  OAI221X4 U359 ( .A0(n1589), .A1(n505), .B0(n1588), .B1(n582), .C0(n1587), 
        .Y(proc_rdata[7]) );
  OAI221X4 U360 ( .A0(n1564), .A1(n505), .B0(n1563), .B1(n582), .C0(n1562), 
        .Y(proc_rdata[2]) );
  OAI221X4 U361 ( .A0(n1609), .A1(n505), .B0(n1608), .B1(n582), .C0(n1607), 
        .Y(proc_rdata[11]) );
  OAI221X4 U362 ( .A0(n1584), .A1(n505), .B0(n1583), .B1(n582), .C0(n1582), 
        .Y(proc_rdata[6]) );
  MX4X2 U363 ( .A(\blocktag[0][20] ), .B(\blocktag[2][20] ), .C(
        \blocktag[1][20] ), .D(\blocktag[3][20] ), .S0(n753), .S1(n726), .Y(
        n872) );
  MX4X2 U364 ( .A(\blocktag[4][20] ), .B(\blocktag[6][20] ), .C(
        \blocktag[5][20] ), .D(\blocktag[7][20] ), .S0(n753), .S1(n726), .Y(
        n871) );
  CLKINVX12 U365 ( .A(N32), .Y(n770) );
  MX4X4 U366 ( .A(\blocktag[3][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[0][13] ), .S0(n762), .S1(n736), .Y(
        n878) );
  MX4X1 U367 ( .A(\block[4][43] ), .B(\block[6][43] ), .C(\block[5][43] ), .D(
        \block[7][43] ), .S0(n759), .S1(n733), .Y(n1138) );
  INVX12 U368 ( .A(n760), .Y(n409) );
  INVXL U369 ( .A(n1535), .Y(n937) );
  CLKINVX12 U370 ( .A(n1775), .Y(n118) );
  CLKINVX20 U371 ( .A(n118), .Y(mem_wdata[126]) );
  CLKINVX12 U372 ( .A(n1812), .Y(n120) );
  CLKINVX20 U373 ( .A(n120), .Y(mem_wdata[80]) );
  BUFX6 U374 ( .A(n55), .Y(n600) );
  CLKINVX20 U375 ( .A(n122), .Y(mem_addr[3]) );
  CLKINVX12 U376 ( .A(n1772), .Y(n124) );
  CLKINVX20 U377 ( .A(n124), .Y(mem_addr[4]) );
  CLKINVX12 U378 ( .A(n1771), .Y(n126) );
  CLKINVX20 U379 ( .A(n126), .Y(mem_addr[5]) );
  CLKINVX12 U380 ( .A(n1770), .Y(n128) );
  CLKINVX20 U381 ( .A(n128), .Y(mem_addr[6]) );
  CLKINVX12 U382 ( .A(n1769), .Y(n130) );
  CLKINVX20 U383 ( .A(n130), .Y(mem_addr[7]) );
  CLKINVX12 U384 ( .A(n1768), .Y(n132) );
  CLKINVX20 U385 ( .A(n132), .Y(mem_addr[8]) );
  CLKINVX12 U386 ( .A(n1767), .Y(n134) );
  CLKINVX20 U387 ( .A(n134), .Y(mem_addr[9]) );
  CLKINVX12 U388 ( .A(n1766), .Y(n136) );
  CLKINVX20 U389 ( .A(n136), .Y(mem_addr[10]) );
  CLKINVX12 U390 ( .A(n1765), .Y(n138) );
  CLKINVX20 U391 ( .A(n138), .Y(mem_addr[11]) );
  CLKINVX12 U392 ( .A(n1764), .Y(n140) );
  CLKINVX20 U393 ( .A(n140), .Y(mem_addr[12]) );
  CLKINVX12 U394 ( .A(n1763), .Y(n142) );
  CLKINVX20 U395 ( .A(n142), .Y(mem_addr[13]) );
  CLKINVX12 U396 ( .A(n1762), .Y(n144) );
  CLKINVX20 U397 ( .A(n144), .Y(mem_addr[14]) );
  CLKINVX12 U398 ( .A(n1761), .Y(n146) );
  CLKINVX20 U399 ( .A(n146), .Y(mem_addr[15]) );
  CLKINVX12 U400 ( .A(n1760), .Y(n148) );
  CLKINVX20 U401 ( .A(n148), .Y(mem_addr[16]) );
  CLKINVX12 U402 ( .A(n1759), .Y(n150) );
  CLKINVX20 U403 ( .A(n150), .Y(mem_addr[17]) );
  CLKINVX12 U404 ( .A(n1758), .Y(n152) );
  CLKINVX20 U405 ( .A(n152), .Y(mem_addr[18]) );
  CLKINVX12 U406 ( .A(n1757), .Y(n154) );
  CLKINVX20 U407 ( .A(n154), .Y(mem_addr[19]) );
  CLKINVX12 U408 ( .A(n1756), .Y(n156) );
  CLKINVX20 U409 ( .A(n156), .Y(mem_addr[20]) );
  CLKINVX12 U410 ( .A(n1755), .Y(n158) );
  CLKINVX20 U411 ( .A(n158), .Y(mem_addr[21]) );
  CLKINVX12 U412 ( .A(n1754), .Y(n160) );
  CLKINVX20 U413 ( .A(n160), .Y(mem_addr[22]) );
  CLKINVX12 U414 ( .A(n1753), .Y(n162) );
  CLKINVX20 U415 ( .A(n162), .Y(mem_addr[23]) );
  CLKINVX20 U416 ( .A(n164), .Y(mem_addr[24]) );
  CLKINVX12 U417 ( .A(n80), .Y(n166) );
  CLKINVX20 U418 ( .A(n166), .Y(mem_addr[26]) );
  CLKINVX12 U419 ( .A(n1750), .Y(n168) );
  CLKINVX20 U420 ( .A(n168), .Y(mem_addr[27]) );
  CLKAND2X12 U421 ( .A(mem_write), .B(n968), .Y(mem_wdata[0]) );
  CLKBUFX20 U422 ( .A(n787), .Y(mem_write) );
  CLKINVX8 U423 ( .A(n1887), .Y(n170) );
  CLKINVX20 U424 ( .A(n170), .Y(mem_wdata[1]) );
  CLKINVX8 U425 ( .A(n1886), .Y(n172) );
  CLKINVX20 U426 ( .A(n172), .Y(mem_wdata[2]) );
  CLKINVX8 U427 ( .A(n1885), .Y(n174) );
  CLKINVX20 U428 ( .A(n174), .Y(mem_wdata[3]) );
  CLKINVX8 U429 ( .A(n1884), .Y(n176) );
  CLKINVX20 U430 ( .A(n176), .Y(mem_wdata[4]) );
  CLKINVX8 U431 ( .A(n1883), .Y(n178) );
  CLKINVX20 U432 ( .A(n178), .Y(mem_wdata[5]) );
  CLKINVX8 U433 ( .A(n1882), .Y(n180) );
  CLKINVX20 U434 ( .A(n180), .Y(mem_wdata[6]) );
  CLKINVX8 U435 ( .A(n1881), .Y(n182) );
  CLKINVX20 U436 ( .A(n182), .Y(mem_wdata[8]) );
  CLKINVX8 U437 ( .A(n1880), .Y(n184) );
  CLKINVX20 U438 ( .A(n184), .Y(mem_wdata[9]) );
  CLKINVX8 U439 ( .A(n1879), .Y(n186) );
  CLKINVX20 U440 ( .A(n186), .Y(mem_wdata[10]) );
  CLKINVX8 U441 ( .A(n1878), .Y(n188) );
  CLKINVX20 U442 ( .A(n188), .Y(mem_wdata[11]) );
  CLKINVX8 U443 ( .A(n1877), .Y(n190) );
  CLKINVX20 U444 ( .A(n190), .Y(mem_wdata[12]) );
  CLKINVX8 U445 ( .A(n1876), .Y(n192) );
  CLKINVX20 U446 ( .A(n192), .Y(mem_wdata[13]) );
  CLKINVX8 U447 ( .A(n1875), .Y(n194) );
  CLKINVX20 U448 ( .A(n194), .Y(mem_wdata[14]) );
  CLKINVX8 U449 ( .A(n1874), .Y(n196) );
  CLKINVX20 U450 ( .A(n196), .Y(mem_wdata[15]) );
  CLKINVX8 U451 ( .A(n1873), .Y(n198) );
  CLKINVX20 U452 ( .A(n198), .Y(mem_wdata[16]) );
  CLKINVX8 U453 ( .A(n1872), .Y(n200) );
  CLKINVX20 U454 ( .A(n200), .Y(mem_wdata[17]) );
  CLKINVX8 U455 ( .A(n1871), .Y(n202) );
  CLKINVX20 U456 ( .A(n202), .Y(mem_wdata[18]) );
  CLKINVX8 U457 ( .A(n1870), .Y(n204) );
  CLKINVX20 U458 ( .A(n204), .Y(mem_wdata[19]) );
  CLKINVX8 U459 ( .A(n1869), .Y(n206) );
  CLKINVX20 U460 ( .A(n206), .Y(mem_wdata[20]) );
  CLKINVX8 U461 ( .A(n1868), .Y(n208) );
  CLKINVX20 U462 ( .A(n208), .Y(mem_wdata[21]) );
  CLKINVX8 U463 ( .A(n1867), .Y(n210) );
  CLKINVX20 U464 ( .A(n210), .Y(mem_wdata[22]) );
  CLKINVX8 U465 ( .A(n1866), .Y(n212) );
  CLKINVX20 U466 ( .A(n212), .Y(mem_wdata[23]) );
  CLKINVX8 U467 ( .A(n1865), .Y(n214) );
  CLKINVX20 U468 ( .A(n214), .Y(mem_wdata[24]) );
  CLKINVX8 U469 ( .A(n1864), .Y(n216) );
  CLKINVX20 U470 ( .A(n216), .Y(mem_wdata[25]) );
  CLKINVX8 U471 ( .A(n1863), .Y(n218) );
  CLKINVX20 U472 ( .A(n218), .Y(mem_wdata[26]) );
  CLKINVX8 U473 ( .A(n1862), .Y(n220) );
  CLKINVX20 U474 ( .A(n220), .Y(mem_wdata[28]) );
  CLKINVX8 U475 ( .A(n1861), .Y(n222) );
  CLKINVX20 U476 ( .A(n222), .Y(mem_wdata[29]) );
  CLKINVX8 U477 ( .A(n1860), .Y(n224) );
  CLKINVX20 U478 ( .A(n224), .Y(mem_wdata[30]) );
  CLKINVX8 U479 ( .A(n1859), .Y(n226) );
  CLKINVX20 U480 ( .A(n226), .Y(mem_wdata[31]) );
  CLKINVX8 U481 ( .A(n1858), .Y(n228) );
  CLKINVX20 U482 ( .A(n228), .Y(mem_wdata[32]) );
  CLKINVX8 U483 ( .A(n1857), .Y(n230) );
  CLKINVX20 U484 ( .A(n230), .Y(mem_wdata[33]) );
  CLKINVX8 U485 ( .A(n1856), .Y(n232) );
  CLKINVX20 U486 ( .A(n232), .Y(mem_wdata[34]) );
  CLKINVX8 U487 ( .A(n1855), .Y(n234) );
  CLKINVX20 U488 ( .A(n234), .Y(mem_wdata[35]) );
  CLKINVX8 U489 ( .A(n1854), .Y(n236) );
  CLKINVX20 U490 ( .A(n236), .Y(mem_wdata[36]) );
  CLKINVX8 U491 ( .A(n1853), .Y(n238) );
  CLKINVX20 U492 ( .A(n238), .Y(mem_wdata[37]) );
  CLKINVX8 U493 ( .A(n1852), .Y(n240) );
  CLKINVX20 U494 ( .A(n240), .Y(mem_wdata[38]) );
  CLKINVX8 U495 ( .A(n1851), .Y(n242) );
  CLKINVX20 U496 ( .A(n242), .Y(mem_wdata[39]) );
  CLKINVX8 U497 ( .A(n1850), .Y(n244) );
  CLKINVX20 U498 ( .A(n244), .Y(mem_wdata[40]) );
  CLKINVX8 U499 ( .A(n1849), .Y(n246) );
  CLKINVX20 U500 ( .A(n246), .Y(mem_wdata[41]) );
  CLKINVX8 U501 ( .A(n1848), .Y(n248) );
  CLKINVX20 U502 ( .A(n248), .Y(mem_wdata[42]) );
  CLKINVX8 U503 ( .A(n1847), .Y(n250) );
  CLKINVX20 U504 ( .A(n250), .Y(mem_wdata[43]) );
  CLKINVX8 U505 ( .A(n1846), .Y(n252) );
  CLKINVX20 U506 ( .A(n252), .Y(mem_wdata[44]) );
  CLKINVX8 U507 ( .A(n1845), .Y(n254) );
  CLKINVX20 U508 ( .A(n254), .Y(mem_wdata[45]) );
  CLKINVX8 U509 ( .A(n1844), .Y(n256) );
  CLKINVX20 U510 ( .A(n256), .Y(mem_wdata[47]) );
  CLKINVX8 U511 ( .A(n1843), .Y(n258) );
  CLKINVX20 U512 ( .A(n258), .Y(mem_wdata[48]) );
  CLKINVX8 U513 ( .A(n1842), .Y(n260) );
  CLKINVX20 U514 ( .A(n260), .Y(mem_wdata[49]) );
  CLKINVX8 U515 ( .A(n1841), .Y(n262) );
  CLKINVX20 U516 ( .A(n262), .Y(mem_wdata[50]) );
  CLKINVX8 U517 ( .A(n1840), .Y(n264) );
  CLKINVX20 U518 ( .A(n264), .Y(mem_wdata[51]) );
  CLKINVX8 U519 ( .A(n1839), .Y(n266) );
  CLKINVX20 U520 ( .A(n266), .Y(mem_wdata[52]) );
  CLKINVX8 U521 ( .A(n1838), .Y(n268) );
  CLKINVX20 U522 ( .A(n268), .Y(mem_wdata[53]) );
  CLKINVX8 U523 ( .A(n1837), .Y(n270) );
  CLKINVX20 U524 ( .A(n270), .Y(mem_wdata[54]) );
  CLKINVX8 U525 ( .A(n1836), .Y(n272) );
  CLKINVX20 U526 ( .A(n272), .Y(mem_wdata[55]) );
  CLKINVX8 U527 ( .A(n1835), .Y(n274) );
  CLKINVX20 U528 ( .A(n274), .Y(mem_wdata[56]) );
  CLKINVX8 U529 ( .A(n1834), .Y(n276) );
  CLKINVX20 U530 ( .A(n276), .Y(mem_wdata[57]) );
  CLKINVX8 U531 ( .A(n1833), .Y(n278) );
  CLKINVX20 U532 ( .A(n278), .Y(mem_wdata[58]) );
  CLKINVX8 U533 ( .A(n1832), .Y(n280) );
  CLKINVX20 U534 ( .A(n280), .Y(mem_wdata[60]) );
  CLKINVX8 U535 ( .A(n1831), .Y(n282) );
  CLKINVX20 U536 ( .A(n282), .Y(mem_wdata[61]) );
  CLKINVX8 U537 ( .A(n1830), .Y(n284) );
  CLKINVX20 U538 ( .A(n284), .Y(mem_wdata[62]) );
  CLKINVX8 U539 ( .A(n1829), .Y(n286) );
  CLKINVX20 U540 ( .A(n286), .Y(mem_wdata[63]) );
  CLKINVX8 U541 ( .A(n1828), .Y(n288) );
  CLKINVX20 U542 ( .A(n288), .Y(mem_wdata[64]) );
  CLKINVX8 U543 ( .A(n1827), .Y(n290) );
  CLKINVX20 U544 ( .A(n290), .Y(mem_wdata[65]) );
  CLKINVX8 U545 ( .A(n1826), .Y(n292) );
  CLKINVX20 U546 ( .A(n292), .Y(mem_wdata[66]) );
  CLKINVX8 U547 ( .A(n1825), .Y(n294) );
  CLKINVX20 U548 ( .A(n294), .Y(mem_wdata[67]) );
  CLKINVX8 U549 ( .A(n1824), .Y(n296) );
  CLKINVX20 U550 ( .A(n296), .Y(mem_wdata[68]) );
  CLKINVX8 U551 ( .A(n1823), .Y(n298) );
  CLKINVX20 U552 ( .A(n298), .Y(mem_wdata[69]) );
  CLKINVX8 U553 ( .A(n1822), .Y(n300) );
  CLKINVX20 U554 ( .A(n300), .Y(mem_wdata[70]) );
  CLKINVX8 U555 ( .A(n1821), .Y(n302) );
  CLKINVX20 U556 ( .A(n302), .Y(mem_wdata[71]) );
  CLKINVX8 U557 ( .A(n1820), .Y(n304) );
  CLKINVX20 U558 ( .A(n304), .Y(mem_wdata[72]) );
  CLKINVX8 U559 ( .A(n1819), .Y(n306) );
  CLKINVX20 U560 ( .A(n306), .Y(mem_wdata[73]) );
  CLKINVX8 U561 ( .A(n1818), .Y(n308) );
  CLKINVX20 U562 ( .A(n308), .Y(mem_wdata[74]) );
  CLKINVX8 U563 ( .A(n1817), .Y(n310) );
  CLKINVX20 U564 ( .A(n310), .Y(mem_wdata[75]) );
  CLKINVX8 U565 ( .A(n1816), .Y(n312) );
  CLKINVX20 U566 ( .A(n312), .Y(mem_wdata[76]) );
  CLKINVX8 U567 ( .A(n1815), .Y(n314) );
  CLKINVX20 U568 ( .A(n314), .Y(mem_wdata[77]) );
  CLKINVX8 U569 ( .A(n1814), .Y(n316) );
  CLKINVX20 U570 ( .A(n316), .Y(mem_wdata[78]) );
  CLKINVX8 U571 ( .A(n1813), .Y(n318) );
  CLKINVX20 U572 ( .A(n318), .Y(mem_wdata[79]) );
  INVX12 U573 ( .A(n1811), .Y(n320) );
  CLKINVX20 U574 ( .A(n320), .Y(mem_wdata[84]) );
  INVX12 U575 ( .A(n1810), .Y(n322) );
  CLKINVX20 U576 ( .A(n322), .Y(mem_wdata[85]) );
  INVX12 U577 ( .A(n1809), .Y(n324) );
  CLKINVX20 U578 ( .A(n324), .Y(mem_wdata[86]) );
  INVX12 U579 ( .A(n1808), .Y(n326) );
  CLKINVX20 U580 ( .A(n326), .Y(mem_wdata[87]) );
  INVX12 U581 ( .A(n1807), .Y(n328) );
  CLKINVX20 U582 ( .A(n328), .Y(mem_wdata[88]) );
  INVX12 U583 ( .A(n1806), .Y(n330) );
  CLKINVX20 U584 ( .A(n330), .Y(mem_wdata[89]) );
  INVX12 U585 ( .A(n1805), .Y(n332) );
  CLKINVX20 U586 ( .A(n332), .Y(mem_wdata[90]) );
  INVX12 U587 ( .A(n1804), .Y(n334) );
  CLKINVX20 U588 ( .A(n334), .Y(mem_wdata[94]) );
  INVX12 U589 ( .A(n1803), .Y(n336) );
  CLKINVX20 U590 ( .A(n336), .Y(mem_wdata[96]) );
  INVX12 U591 ( .A(n1802), .Y(n338) );
  CLKINVX20 U592 ( .A(n338), .Y(mem_wdata[97]) );
  INVX12 U593 ( .A(n1801), .Y(n340) );
  CLKINVX20 U594 ( .A(n340), .Y(mem_wdata[98]) );
  INVX12 U595 ( .A(n1800), .Y(n342) );
  CLKINVX20 U596 ( .A(n342), .Y(mem_wdata[99]) );
  INVX12 U597 ( .A(n1799), .Y(n344) );
  CLKINVX20 U598 ( .A(n344), .Y(mem_wdata[100]) );
  INVX12 U599 ( .A(n1798), .Y(n346) );
  CLKINVX20 U600 ( .A(n346), .Y(mem_wdata[101]) );
  INVX12 U601 ( .A(n1797), .Y(n348) );
  CLKINVX20 U602 ( .A(n348), .Y(mem_wdata[102]) );
  INVX12 U603 ( .A(n1796), .Y(n350) );
  CLKINVX20 U604 ( .A(n350), .Y(mem_wdata[103]) );
  INVX12 U605 ( .A(n1795), .Y(n352) );
  CLKINVX20 U606 ( .A(n352), .Y(mem_wdata[104]) );
  INVX12 U607 ( .A(n1794), .Y(n354) );
  CLKINVX20 U608 ( .A(n354), .Y(mem_wdata[105]) );
  INVX12 U609 ( .A(n1793), .Y(n356) );
  CLKINVX20 U610 ( .A(n356), .Y(mem_wdata[106]) );
  INVX12 U611 ( .A(n1792), .Y(n358) );
  CLKINVX20 U612 ( .A(n358), .Y(mem_wdata[107]) );
  INVX12 U613 ( .A(n1791), .Y(n360) );
  CLKINVX20 U614 ( .A(n360), .Y(mem_wdata[108]) );
  INVX12 U615 ( .A(n1790), .Y(n362) );
  CLKINVX20 U616 ( .A(n362), .Y(mem_wdata[109]) );
  INVX12 U617 ( .A(n1789), .Y(n364) );
  CLKINVX20 U618 ( .A(n364), .Y(mem_wdata[110]) );
  INVX12 U619 ( .A(n1788), .Y(n366) );
  CLKINVX20 U620 ( .A(n366), .Y(mem_wdata[111]) );
  INVX12 U621 ( .A(n1787), .Y(n368) );
  CLKINVX20 U622 ( .A(n368), .Y(mem_wdata[112]) );
  INVX12 U623 ( .A(n1786), .Y(n370) );
  CLKINVX20 U624 ( .A(n370), .Y(mem_wdata[113]) );
  INVX12 U625 ( .A(n1785), .Y(n372) );
  CLKINVX20 U626 ( .A(n372), .Y(mem_wdata[114]) );
  INVX12 U627 ( .A(n1784), .Y(n374) );
  CLKINVX20 U628 ( .A(n374), .Y(mem_wdata[115]) );
  INVX12 U629 ( .A(n1783), .Y(n376) );
  CLKINVX20 U630 ( .A(n376), .Y(mem_wdata[116]) );
  INVX12 U631 ( .A(n1782), .Y(n378) );
  CLKINVX20 U632 ( .A(n378), .Y(mem_wdata[117]) );
  INVX12 U633 ( .A(n1781), .Y(n380) );
  CLKINVX20 U634 ( .A(n380), .Y(mem_wdata[118]) );
  INVX12 U635 ( .A(n1780), .Y(n382) );
  CLKINVX20 U636 ( .A(n382), .Y(mem_wdata[119]) );
  INVX12 U637 ( .A(n1779), .Y(n384) );
  CLKINVX20 U638 ( .A(n384), .Y(mem_wdata[120]) );
  INVX12 U639 ( .A(n1778), .Y(n386) );
  CLKINVX20 U640 ( .A(n386), .Y(mem_wdata[121]) );
  INVX12 U641 ( .A(n1777), .Y(n388) );
  CLKINVX20 U642 ( .A(n388), .Y(mem_wdata[122]) );
  CLKINVX20 U643 ( .A(n390), .Y(mem_wdata[125]) );
  INVX8 U644 ( .A(n1774), .Y(n392) );
  CLKINVX20 U645 ( .A(n392), .Y(mem_addr[1]) );
  CLKAND2X12 U646 ( .A(n1519), .B(n780), .Y(mem_addr[2]) );
  AOI221X2 U647 ( .A0(n796), .A1(n1538), .B0(n965), .B1(n1542), .C0(n67), .Y(
        n395) );
  INVX8 U648 ( .A(n1545), .Y(n1542) );
  BUFX20 U649 ( .A(n769), .Y(n764) );
  XOR2X4 U650 ( .A(n419), .B(n396), .Y(n525) );
  MXI4X4 U651 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n532), .S1(n724), 
        .Y(n823) );
  MXI2X4 U652 ( .A(n841), .B(n842), .S0(n398), .Y(n417) );
  XNOR2X4 U653 ( .A(n399), .B(n884), .Y(n818) );
  MXI2X4 U654 ( .A(n805), .B(n804), .S0(n780), .Y(n399) );
  MX2X6 U655 ( .A(n872), .B(n871), .S0(n779), .Y(n1534) );
  MXI2X4 U656 ( .A(n400), .B(n401), .S0(n779), .Y(n1531) );
  MX4X1 U657 ( .A(n431), .B(n432), .C(n433), .D(n434), .S0(n765), .S1(n741), 
        .Y(n401) );
  CLKMX2X6 U658 ( .A(n838), .B(n837), .S0(n779), .Y(n1528) );
  XOR2X4 U659 ( .A(n417), .B(n403), .Y(n843) );
  INVX2 U660 ( .A(n439), .Y(n404) );
  INVX16 U661 ( .A(n762), .Y(n444) );
  INVX16 U662 ( .A(n762), .Y(n754) );
  CLKMX2X6 U663 ( .A(n852), .B(n851), .S0(n779), .Y(n1521) );
  MXI4X2 U664 ( .A(\blocktag[7][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[4][22] ), .S0(n768), .S1(n738), .Y(
        n861) );
  INVX16 U665 ( .A(n744), .Y(n726) );
  CLKINVX4 U666 ( .A(n925), .Y(n405) );
  INVXL U667 ( .A(n1532), .Y(n925) );
  INVXL U668 ( .A(n1537), .Y(n943) );
  XOR2X4 U669 ( .A(n406), .B(n898), .Y(n826) );
  MXI2X4 U670 ( .A(n821), .B(n822), .S0(n435), .Y(n406) );
  CLKINVX2 U671 ( .A(proc_addr[11]), .Y(n898) );
  INVXL U672 ( .A(n1523), .Y(n407) );
  NAND2X8 U673 ( .A(n521), .B(n1543), .Y(n520) );
  CLKMX2X6 U674 ( .A(n864), .B(n863), .S0(n779), .Y(n1532) );
  BUFX8 U675 ( .A(n520), .Y(n582) );
  MXI2XL U676 ( .A(n820), .B(n819), .S0(n780), .Y(n416) );
  MX4X1 U677 ( .A(\block[2][95] ), .B(\block[0][95] ), .C(\block[3][95] ), .D(
        \block[1][95] ), .S0(n766), .S1(n734), .Y(n1348) );
  INVX4 U678 ( .A(n765), .Y(n748) );
  MXI4X2 U679 ( .A(n420), .B(n421), .C(n422), .D(n423), .S0(n763), .S1(n726), 
        .Y(n859) );
  MXI2XL U680 ( .A(n830), .B(n829), .S0(n779), .Y(n424) );
  MXI4X4 U681 ( .A(n425), .B(n426), .C(n427), .D(n428), .S0(n751), .S1(n725), 
        .Y(n842) );
  BUFX20 U682 ( .A(n767), .Y(n768) );
  CLKBUFX2 U683 ( .A(n1530), .Y(n429) );
  INVX4 U684 ( .A(n765), .Y(n755) );
  CLKAND2X12 U685 ( .A(mem_write), .B(n1495), .Y(mem_wdata[123]) );
  INVX4 U686 ( .A(n1495), .Y(n1688) );
  MX2X1 U687 ( .A(n1492), .B(n1491), .S0(n772), .Y(n1495) );
  INVX1 U688 ( .A(n743), .Y(n438) );
  BUFX20 U689 ( .A(n745), .Y(n743) );
  INVXL U690 ( .A(n25), .Y(n922) );
  BUFX20 U691 ( .A(n767), .Y(n532) );
  CLKINVX2 U692 ( .A(n912), .Y(n440) );
  MXI4X4 U693 ( .A(n461), .B(n462), .C(n459), .D(n460), .S0(n751), .S1(n738), 
        .Y(n819) );
  INVXL U694 ( .A(n418), .Y(n885) );
  MX4X4 U695 ( .A(\blocktag[4][8] ), .B(\blocktag[6][8] ), .C(\blocktag[5][8] ), .D(\blocktag[7][8] ), .S0(n752), .S1(n725), .Y(n841) );
  CLKBUFX12 U696 ( .A(n744), .Y(n736) );
  INVXL U697 ( .A(n1521), .Y(n940) );
  INVXL U698 ( .A(n1527), .Y(n927) );
  CLKMX2X6 U699 ( .A(n840), .B(n839), .S0(n779), .Y(n1526) );
  CLKINVX2 U700 ( .A(n424), .Y(n443) );
  XOR2X4 U701 ( .A(n1534), .B(n445), .Y(n876) );
  XOR2X4 U702 ( .A(n1526), .B(n446), .Y(n844) );
  CLKBUFX3 U703 ( .A(n520), .Y(n583) );
  INVXL U704 ( .A(n1529), .Y(n912) );
  CLKINVX6 U705 ( .A(n1542), .Y(n447) );
  CLKMX2X6 U706 ( .A(n798), .B(n797), .S0(n772), .Y(n1545) );
  CLKINVX2 U707 ( .A(n909), .Y(n448) );
  XOR2X4 U708 ( .A(n1522), .B(n921), .Y(n867) );
  CLKINVX3 U709 ( .A(proc_addr[6]), .Y(n921) );
  XOR2X4 U710 ( .A(n1528), .B(proc_addr[16]), .Y(n845) );
  INVXL U711 ( .A(n2), .Y(n453) );
  MXI4X4 U712 ( .A(n454), .B(n455), .C(n456), .D(n457), .S0(n441), .S1(n728), 
        .Y(n877) );
  MX4X2 U713 ( .A(\blocktag[0][12] ), .B(\blocktag[2][12] ), .C(
        \blocktag[1][12] ), .D(\blocktag[3][12] ), .S0(n415), .S1(n724), .Y(
        n832) );
  INVX20 U714 ( .A(n736), .Y(n734) );
  XOR2X4 U715 ( .A(n1527), .B(n926), .Y(n870) );
  CLKINVX2 U716 ( .A(proc_addr[15]), .Y(n926) );
  CLKBUFX2 U717 ( .A(n1531), .Y(n458) );
  XOR2X4 U718 ( .A(n1537), .B(n942), .Y(n858) );
  CLKINVX2 U719 ( .A(proc_addr[29]), .Y(n942) );
  MX4X4 U720 ( .A(\blocktag[2][3] ), .B(\blocktag[0][3] ), .C(\blocktag[3][3] ), .D(\blocktag[1][3] ), .S0(n532), .S1(n723), .Y(n805) );
  INVXL U721 ( .A(n437), .Y(n889) );
  XOR2X4 U722 ( .A(n1535), .B(n936), .Y(n855) );
  CLKINVX2 U723 ( .A(proc_addr[26]), .Y(n936) );
  CLKINVX2 U724 ( .A(proc_addr[24]), .Y(n930) );
  MXI4X4 U725 ( .A(n510), .B(n511), .C(n512), .D(n513), .S0(n761), .S1(n723), 
        .Y(n833) );
  XOR2X4 U726 ( .A(n1524), .B(n514), .Y(n825) );
  BUFX20 U727 ( .A(n770), .Y(n769) );
  XOR2X4 U728 ( .A(n1521), .B(n939), .Y(n856) );
  CLKINVX3 U729 ( .A(proc_addr[5]), .Y(n939) );
  INVX20 U730 ( .A(n761), .Y(n752) );
  CLKINVX2 U731 ( .A(proc_addr[25]), .Y(n933) );
  INVXL U732 ( .A(n18), .Y(n894) );
  MX4X4 U733 ( .A(\blocktag[6][3] ), .B(\blocktag[4][3] ), .C(\blocktag[7][3] ), .D(\blocktag[5][3] ), .S0(n532), .S1(n723), .Y(n804) );
  BUFX8 U734 ( .A(n91), .Y(n579) );
  BUFX8 U735 ( .A(n579), .Y(n581) );
  CLKINVX2 U736 ( .A(n416), .Y(n522) );
  INVX8 U737 ( .A(n539), .Y(n540) );
  NAND3X8 U738 ( .A(n835), .B(n525), .C(n836), .Y(n846) );
  OAI221X4 U739 ( .A0(n1704), .A1(n548), .B0(n1513), .B1(n553), .C0(n1220), 
        .Y(block_next[63]) );
  BUFX12 U740 ( .A(n70), .Y(n548) );
  OAI221X4 U741 ( .A0(n1695), .A1(n548), .B0(n1502), .B1(n553), .C0(n1212), 
        .Y(block_next[61]) );
  OAI221X4 U742 ( .A0(n1685), .A1(n548), .B0(n1494), .B1(n553), .C0(n1204), 
        .Y(block_next[59]) );
  OAI221X4 U743 ( .A0(n1690), .A1(n548), .B0(n1499), .B1(n553), .C0(n1208), 
        .Y(block_next[60]) );
  OAI221X4 U744 ( .A0(n1699), .A1(n548), .B0(n1507), .B1(n553), .C0(n1216), 
        .Y(block_next[62]) );
  OAI221X4 U745 ( .A0(n1660), .A1(n547), .B0(n1469), .B1(n553), .C0(n1184), 
        .Y(block_next[54]) );
  OAI221X4 U746 ( .A0(n1655), .A1(n547), .B0(n1464), .B1(n553), .C0(n1180), 
        .Y(block_next[53]) );
  OAI221X4 U747 ( .A0(n1680), .A1(n548), .B0(n1489), .B1(n553), .C0(n1200), 
        .Y(block_next[58]) );
  OAI221X4 U748 ( .A0(n1675), .A1(n547), .B0(n1484), .B1(n553), .C0(n1196), 
        .Y(block_next[57]) );
  OAI221X4 U749 ( .A0(n1670), .A1(n547), .B0(n1479), .B1(n554), .C0(n1192), 
        .Y(block_next[56]) );
  OAI221X4 U750 ( .A0(n1665), .A1(n547), .B0(n1474), .B1(n553), .C0(n1188), 
        .Y(block_next[55]) );
  OAI221X4 U751 ( .A0(n1551), .A1(n549), .B0(n1359), .B1(n557), .C0(n1225), 
        .Y(block_next[64]) );
  OAI221X4 U752 ( .A0(n1556), .A1(n549), .B0(n1364), .B1(n557), .C0(n1229), 
        .Y(block_next[65]) );
  BUFX16 U753 ( .A(n1350), .Y(n549) );
  XOR2X4 U754 ( .A(n1532), .B(n924), .Y(n868) );
  BUFX16 U755 ( .A(n785), .Y(n783) );
  NOR2BX4 U756 ( .AN(n1544), .B(n1542), .Y(n523) );
  CLKINVX2 U757 ( .A(proc_addr[22]), .Y(n924) );
  CLKINVX12 U758 ( .A(n1540), .Y(n1547) );
  CLKINVX2 U759 ( .A(proc_addr[20]), .Y(n919) );
  XOR2X4 U760 ( .A(n1523), .B(n524), .Y(n816) );
  CLKINVX2 U761 ( .A(proc_addr[13]), .Y(n902) );
  XOR2X4 U762 ( .A(n1529), .B(n911), .Y(n836) );
  CLKINVX2 U763 ( .A(proc_addr[17]), .Y(n911) );
  OAI221X4 U764 ( .A0(n1645), .A1(n547), .B0(n1454), .B1(n553), .C0(n1172), 
        .Y(block_next[51]) );
  OAI221X4 U765 ( .A0(n1499), .A1(n551), .B0(n1694), .B1(n546), .C0(n1079), 
        .Y(block_next[28]) );
  OAI221X4 U766 ( .A0(n1595), .A1(n548), .B0(n1404), .B1(n554), .C0(n1132), 
        .Y(block_next[41]) );
  OAI221X4 U767 ( .A0(n1625), .A1(n547), .B0(n1434), .B1(n554), .C0(n1156), 
        .Y(block_next[47]) );
  OAI221X4 U768 ( .A0(n1600), .A1(n548), .B0(n1409), .B1(n554), .C0(n1136), 
        .Y(block_next[42]) );
  OAI221X4 U769 ( .A0(n1590), .A1(n548), .B0(n1399), .B1(n554), .C0(n1128), 
        .Y(block_next[40]) );
  OAI221X4 U770 ( .A0(n1580), .A1(n548), .B0(n1389), .B1(n554), .C0(n1120), 
        .Y(block_next[38]) );
  OAI221X4 U771 ( .A0(n1555), .A1(n548), .B0(n1364), .B1(n1355), .C0(n1100), 
        .Y(block_next[33]) );
  OAI221X4 U772 ( .A0(n1507), .A1(n551), .B0(n1703), .B1(n546), .C0(n1087), 
        .Y(block_next[30]) );
  OAI221X4 U773 ( .A0(n1550), .A1(n548), .B0(n1359), .B1(n554), .C0(n1096), 
        .Y(block_next[32]) );
  OAI221X4 U774 ( .A0(n1615), .A1(n547), .B0(n1424), .B1(n554), .C0(n1148), 
        .Y(block_next[45]) );
  OAI221X4 U775 ( .A0(n1570), .A1(n548), .B0(n1379), .B1(n554), .C0(n1112), 
        .Y(block_next[36]) );
  OAI221X4 U776 ( .A0(n1575), .A1(n548), .B0(n1384), .B1(n554), .C0(n1116), 
        .Y(block_next[37]) );
  OAI221X4 U777 ( .A0(n1560), .A1(n548), .B0(n1369), .B1(n554), .C0(n1104), 
        .Y(block_next[34]) );
  OAI221X4 U778 ( .A0(n1605), .A1(n548), .B0(n1414), .B1(n554), .C0(n1140), 
        .Y(block_next[43]) );
  OAI221X4 U779 ( .A0(n1494), .A1(n551), .B0(n1689), .B1(n546), .C0(n1075), 
        .Y(block_next[27]) );
  OAI221X4 U780 ( .A0(n1585), .A1(n548), .B0(n1394), .B1(n554), .C0(n1124), 
        .Y(block_next[39]) );
  OAI221X4 U781 ( .A0(n1513), .A1(n551), .B0(n1710), .B1(n546), .C0(n1091), 
        .Y(block_next[31]) );
  OAI221X4 U782 ( .A0(n1650), .A1(n547), .B0(n1459), .B1(n553), .C0(n1176), 
        .Y(block_next[52]) );
  OAI221X4 U783 ( .A0(n1640), .A1(n547), .B0(n1449), .B1(n554), .C0(n1168), 
        .Y(block_next[50]) );
  OAI221X4 U784 ( .A0(n1635), .A1(n547), .B0(n1444), .B1(n554), .C0(n1164), 
        .Y(block_next[49]) );
  OAI221X4 U785 ( .A0(n1630), .A1(n547), .B0(n1439), .B1(n554), .C0(n1160), 
        .Y(block_next[48]) );
  OAI221X4 U786 ( .A0(n1610), .A1(n548), .B0(n1419), .B1(n554), .C0(n1144), 
        .Y(block_next[44]) );
  OAI221X4 U787 ( .A0(n1502), .A1(n551), .B0(n1698), .B1(n546), .C0(n1083), 
        .Y(block_next[29]) );
  BUFX12 U788 ( .A(n1092), .Y(n546) );
  OAI221X4 U789 ( .A0(n1620), .A1(n547), .B0(n1429), .B1(n554), .C0(n1152), 
        .Y(block_next[46]) );
  OAI221X4 U790 ( .A0(n1565), .A1(n548), .B0(n1374), .B1(n554), .C0(n1108), 
        .Y(block_next[35]) );
  CLKINVX2 U791 ( .A(proc_addr[19]), .Y(n914) );
  CLKINVX2 U792 ( .A(proc_addr[23]), .Y(n888) );
  CLKAND2X12 U793 ( .A(mem_write), .B(n1500), .Y(mem_wdata[124]) );
  INVX8 U794 ( .A(n1500), .Y(n1693) );
  CLKMX2X8 U795 ( .A(n1497), .B(n1496), .S0(n772), .Y(n1500) );
  CLKINVX2 U796 ( .A(proc_addr[10]), .Y(n893) );
  CLKINVX2 U797 ( .A(proc_addr[8]), .Y(n884) );
  NOR4X8 U798 ( .A(n846), .B(n844), .C(n843), .D(n845), .Y(n847) );
  MX2X4 U799 ( .A(n528), .B(n529), .S0(n772), .Y(n527) );
  MXI4XL U800 ( .A(\block[0][125] ), .B(\block[2][125] ), .C(\block[1][125] ), 
        .D(\block[3][125] ), .S0(n750), .S1(n722), .Y(n528) );
  MXI4XL U801 ( .A(\block[4][125] ), .B(\block[6][125] ), .C(\block[5][125] ), 
        .D(\block[7][125] ), .S0(n750), .S1(n722), .Y(n529) );
  NAND4X8 U802 ( .A(n530), .B(n531), .C(n881), .D(n882), .Y(n1541) );
  AND4X8 U803 ( .A(n857), .B(n858), .C(n855), .D(n856), .Y(n530) );
  CLKINVX2 U804 ( .A(proc_addr[12]), .Y(n905) );
  CLKINVX2 U805 ( .A(proc_addr[9]), .Y(n895) );
  AND2X4 U806 ( .A(mem_write), .B(n1516), .Y(mem_wdata[127]) );
  INVX8 U807 ( .A(n1516), .Y(n1708) );
  MX4X4 U808 ( .A(\blocktag[0][10] ), .B(\blocktag[2][10] ), .C(
        \blocktag[1][10] ), .D(\blocktag[3][10] ), .S0(n753), .S1(n726), .Y(
        n860) );
  MX4X2 U809 ( .A(\blocktag[4][19] ), .B(\blocktag[6][19] ), .C(
        \blocktag[5][19] ), .D(\blocktag[7][19] ), .S0(n442), .S1(n724), .Y(
        n873) );
  INVX20 U810 ( .A(n763), .Y(n753) );
  NOR2X8 U811 ( .A(n875), .B(n876), .Y(n882) );
  MX4X2 U812 ( .A(\blocktag[4][24] ), .B(\blocktag[6][24] ), .C(
        \blocktag[5][24] ), .D(\blocktag[7][24] ), .S0(n752), .S1(n725), .Y(
        n849) );
  CLKINVX16 U813 ( .A(n771), .Y(n785) );
  BUFX20 U814 ( .A(n785), .Y(n784) );
  BUFX8 U815 ( .A(n785), .Y(n782) );
  INVX4 U816 ( .A(n532), .Y(n750) );
  NOR2X8 U817 ( .A(n880), .B(n879), .Y(n881) );
  MX4X2 U818 ( .A(\blocktag[0][11] ), .B(\blocktag[2][11] ), .C(
        \blocktag[1][11] ), .D(\blocktag[3][11] ), .S0(n415), .S1(n725), .Y(
        n838) );
  BUFX20 U819 ( .A(N33), .Y(n771) );
  CLKINVX2 U820 ( .A(proc_addr[7]), .Y(n891) );
  NAND2X2 U821 ( .A(n22), .B(n1546), .Y(n967) );
  NOR4X8 U822 ( .A(n828), .B(n825), .C(n826), .D(n827), .Y(n848) );
  CLKMX2X6 U823 ( .A(n860), .B(n859), .S0(n779), .Y(n1527) );
  MX4X2 U824 ( .A(\blocktag[0][0] ), .B(\blocktag[2][0] ), .C(\blocktag[1][0] ), .D(\blocktag[3][0] ), .S0(n752), .S1(n725), .Y(n852) );
  OAI221X4 U825 ( .A0(n1561), .A1(n549), .B0(n1369), .B1(n557), .C0(n1233), 
        .Y(block_next[66]) );
  NAND2X8 U826 ( .A(n793), .B(n1538), .Y(n1539) );
  NAND3X8 U827 ( .A(n1546), .B(n1547), .C(n78), .Y(n1549) );
  CLKINVX8 U828 ( .A(proc_addr[0]), .Y(n1544) );
  NAND4BX2 U829 ( .AN(n1517), .B(n967), .C(n966), .D(n965), .Y(n1518) );
  CLKAND2X12 U830 ( .A(n789), .B(n996), .Y(mem_wdata[7]) );
  BUFX20 U831 ( .A(n767), .Y(n763) );
  BUFX20 U832 ( .A(n769), .Y(n761) );
  NAND3BX4 U833 ( .AN(mem_ready), .B(proc_stall), .C(n1517), .Y(n1520) );
  CLKINVX2 U834 ( .A(n1520), .Y(n1748) );
  AND2XL U835 ( .A(n735), .B(n1519), .Y(mem_addr[0]) );
  BUFX20 U836 ( .A(n787), .Y(n789) );
  NAND2X6 U837 ( .A(n946), .B(n447), .Y(n1517) );
  CLKMX2X4 U838 ( .A(n807), .B(n806), .S0(n780), .Y(n946) );
  OA22X1 U839 ( .A0(n1581), .A1(n579), .B0(n1580), .B1(n540), .Y(n1582) );
  INVX20 U840 ( .A(n738), .Y(n711) );
  BUFX20 U841 ( .A(n787), .Y(n791) );
  CLKAND2X12 U842 ( .A(n791), .B(n1153), .Y(mem_wdata[46]) );
  CLKMX2X4 U843 ( .A(n1505), .B(n1504), .S0(n772), .Y(n1508) );
  BUFX20 U844 ( .A(n768), .Y(n762) );
  INVX20 U845 ( .A(n738), .Y(n728) );
  AND2X8 U846 ( .A(mem_write), .B(n1508), .Y(n1775) );
  BUFX20 U847 ( .A(n1749), .Y(n790) );
  AND2X8 U848 ( .A(n790), .B(n1290), .Y(n1812) );
  AND2XL U849 ( .A(n790), .B(n1294), .Y(mem_wdata[81]) );
  AND2XL U850 ( .A(n790), .B(n1298), .Y(mem_wdata[82]) );
  AND2XL U851 ( .A(n790), .B(n1302), .Y(mem_wdata[83]) );
  NAND2X8 U852 ( .A(n847), .B(n848), .Y(n1540) );
  CLKMX2X2 U853 ( .A(n407), .B(n891), .S0(n568), .Y(n892) );
  BUFX20 U854 ( .A(n770), .Y(n767) );
  NAND2X2 U855 ( .A(proc_addr[1]), .B(proc_addr[0]), .Y(n961) );
  AO22XL U856 ( .A0(proc_addr[27]), .A1(mem_read), .B0(mem_write), .B1(n453), 
        .Y(n1751) );
  CLKAND2X12 U857 ( .A(n790), .B(n1205), .Y(mem_wdata[59]) );
  CLKAND2X12 U858 ( .A(n791), .B(n1076), .Y(mem_wdata[27]) );
  CLKAND2X12 U859 ( .A(n789), .B(n1351), .Y(mem_wdata[95]) );
  CLKAND2X12 U860 ( .A(n789), .B(n1342), .Y(mem_wdata[93]) );
  CLKAND2X12 U861 ( .A(n789), .B(n1338), .Y(mem_wdata[92]) );
  CLKAND2X12 U862 ( .A(n789), .B(n1334), .Y(mem_wdata[91]) );
  BUFX8 U863 ( .A(n628), .Y(n623) );
  CLKBUFX6 U864 ( .A(n628), .Y(n624) );
  CLKBUFX4 U865 ( .A(n61), .Y(n648) );
  BUFX3 U866 ( .A(n585), .Y(n599) );
  NAND2XL U867 ( .A(n1747), .B(n739), .Y(n802) );
  BUFX12 U868 ( .A(n579), .Y(n580) );
  INVXL U869 ( .A(n1052), .Y(n1659) );
  INVXL U870 ( .A(n1056), .Y(n1664) );
  NAND2XL U871 ( .A(mem_rdata[0]), .B(n570), .Y(n964) );
  INVX1 U872 ( .A(n736), .Y(n544) );
  INVX2 U873 ( .A(n1197), .Y(n1675) );
  INVX2 U874 ( .A(n1193), .Y(n1670) );
  INVX3 U875 ( .A(n1262), .Y(n1596) );
  INVX3 U876 ( .A(n1133), .Y(n1595) );
  INVX3 U877 ( .A(n1004), .Y(n1599) );
  INVX3 U878 ( .A(n1189), .Y(n1665) );
  CLKINVX8 U879 ( .A(n887), .Y(n1711) );
  INVX3 U880 ( .A(n1508), .Y(n1702) );
  CLKINVX1 U881 ( .A(n1326), .Y(n1676) );
  CLKINVX1 U882 ( .A(n1310), .Y(n1656) );
  INVX1 U883 ( .A(n1068), .Y(n1679) );
  INVX1 U884 ( .A(n1485), .Y(n1678) );
  INVXL U885 ( .A(n1470), .Y(n1663) );
  CLKINVX1 U886 ( .A(n1302), .Y(n1646) );
  CLKINVX1 U887 ( .A(n1173), .Y(n1645) );
  CLKINVX1 U888 ( .A(n1181), .Y(n1655) );
  CLKINVX1 U889 ( .A(n1161), .Y(n1630) );
  CLKINVX1 U890 ( .A(n1185), .Y(n1660) );
  CLKINVX3 U891 ( .A(n1165), .Y(n1635) );
  NAND2X1 U892 ( .A(mem_rdata[90]), .B(n565), .Y(n1329) );
  MX4X1 U893 ( .A(\block[4][47] ), .B(\block[6][47] ), .C(\block[5][47] ), .D(
        \block[7][47] ), .S0(n760), .S1(n734), .Y(n1154) );
  MX4X1 U894 ( .A(\block[4][111] ), .B(\block[6][111] ), .C(\block[5][111] ), 
        .D(\block[7][111] ), .S0(n749), .S1(n720), .Y(n1431) );
  MX4X1 U895 ( .A(\block[4][46] ), .B(\block[6][46] ), .C(\block[5][46] ), .D(
        \block[7][46] ), .S0(n760), .S1(n734), .Y(n1150) );
  MX4X1 U896 ( .A(\block[4][75] ), .B(\block[6][75] ), .C(\block[5][75] ), .D(
        \block[7][75] ), .S0(n754), .S1(n715), .Y(n1267) );
  CLKBUFX4 U897 ( .A(n645), .Y(n643) );
  CLKBUFX4 U898 ( .A(n627), .Y(n625) );
  CLKBUFX4 U899 ( .A(n679), .Y(n677) );
  CLKBUFX4 U900 ( .A(n709), .Y(n707) );
  CLKBUFX4 U901 ( .A(n650), .Y(n661) );
  CLKBUFX4 U902 ( .A(n694), .Y(n692) );
  CLKBUFX4 U903 ( .A(n600), .Y(n612) );
  CLKBUFX4 U904 ( .A(n584), .Y(n595) );
  BUFX4 U905 ( .A(n627), .Y(n631) );
  CLKBUFX2 U906 ( .A(n64), .Y(n632) );
  BUFX4 U907 ( .A(n681), .Y(n696) );
  INVX3 U908 ( .A(n801), .Y(n952) );
  NAND2XL U909 ( .A(n1745), .B(n734), .Y(n801) );
  NOR2XL U910 ( .A(n772), .B(n760), .Y(n1744) );
  INVX3 U911 ( .A(n800), .Y(n951) );
  NAND2XL U912 ( .A(n1744), .B(n736), .Y(n800) );
  NAND2X4 U913 ( .A(n951), .B(n794), .Y(n887) );
  CLKINVX4 U914 ( .A(n802), .Y(n953) );
  OA22XL U915 ( .A0(n1591), .A1(n579), .B0(n1590), .B1(n540), .Y(n1592) );
  OA22XL U916 ( .A0(n1606), .A1(n579), .B0(n1605), .B1(n540), .Y(n1607) );
  OA22XL U917 ( .A0(n1611), .A1(n579), .B0(n1610), .B1(n540), .Y(n1612) );
  OA22XL U918 ( .A0(n1586), .A1(n581), .B0(n1585), .B1(n540), .Y(n1587) );
  OA22XL U919 ( .A0(n1576), .A1(n579), .B0(n1575), .B1(n540), .Y(n1577) );
  OA22XL U920 ( .A0(n1561), .A1(n579), .B0(n1560), .B1(n540), .Y(n1562) );
  OA22XL U921 ( .A0(n1551), .A1(n579), .B0(n1550), .B1(n540), .Y(n1552) );
  OA22XL U922 ( .A0(n1566), .A1(n579), .B0(n1565), .B1(n540), .Y(n1567) );
  OA22XL U923 ( .A0(n1556), .A1(n579), .B0(n1555), .B1(n540), .Y(n1557) );
  OA22XL U924 ( .A0(n1626), .A1(n579), .B0(n1625), .B1(n540), .Y(n1627) );
  OA22XL U925 ( .A0(n1621), .A1(n579), .B0(n1620), .B1(n540), .Y(n1622) );
  OA22XL U926 ( .A0(n1571), .A1(n579), .B0(n1570), .B1(n540), .Y(n1572) );
  OA22XL U927 ( .A0(n1656), .A1(n580), .B0(n1655), .B1(n540), .Y(n1657) );
  OA22XL U928 ( .A0(n1646), .A1(n580), .B0(n1645), .B1(n540), .Y(n1647) );
  OA22XL U929 ( .A0(n1661), .A1(n580), .B0(n1660), .B1(n540), .Y(n1662) );
  OA22XL U930 ( .A0(n1641), .A1(n580), .B0(n1640), .B1(n540), .Y(n1642) );
  OA22XL U931 ( .A0(n1651), .A1(n580), .B0(n1650), .B1(n540), .Y(n1652) );
  OA22XL U932 ( .A0(n1631), .A1(n580), .B0(n1630), .B1(n540), .Y(n1632) );
  OA22XL U933 ( .A0(n1636), .A1(n580), .B0(n1635), .B1(n540), .Y(n1637) );
  OA22XL U934 ( .A0(n1666), .A1(n580), .B0(n1665), .B1(n540), .Y(n1667) );
  OA22XL U935 ( .A0(n1681), .A1(n580), .B0(n1680), .B1(n540), .Y(n1682) );
  INVX3 U936 ( .A(n1405), .Y(n1598) );
  INVXL U937 ( .A(n946), .Y(n947) );
  INVX3 U938 ( .A(n1360), .Y(n1553) );
  INVX3 U939 ( .A(n1395), .Y(n1588) );
  INVX3 U940 ( .A(n1375), .Y(n1568) );
  INVX3 U941 ( .A(n1385), .Y(n1578) );
  INVX3 U942 ( .A(n1365), .Y(n1558) );
  INVX3 U943 ( .A(n1370), .Y(n1563) );
  INVX3 U944 ( .A(n1435), .Y(n1628) );
  INVX3 U945 ( .A(n1430), .Y(n1623) );
  INVX3 U946 ( .A(n1400), .Y(n1593) );
  INVX3 U947 ( .A(n1380), .Y(n1573) );
  INVX3 U948 ( .A(n968), .Y(n1554) );
  INVX3 U949 ( .A(n1415), .Y(n1608) );
  INVX3 U950 ( .A(n1410), .Y(n1603) );
  INVX3 U951 ( .A(n1390), .Y(n1583) );
  INVX3 U952 ( .A(n1425), .Y(n1618) );
  INVX3 U953 ( .A(n1420), .Y(n1613) );
  INVX3 U954 ( .A(n1286), .Y(n1626) );
  INVX3 U955 ( .A(n1282), .Y(n1621) );
  INVX3 U956 ( .A(n1278), .Y(n1616) );
  INVX3 U957 ( .A(n1274), .Y(n1611) );
  INVX3 U958 ( .A(n1226), .Y(n1551) );
  INVX3 U959 ( .A(n1238), .Y(n1566) );
  INVX3 U960 ( .A(n1254), .Y(n1586) );
  INVX3 U961 ( .A(n1246), .Y(n1576) );
  INVX3 U962 ( .A(n1230), .Y(n1556) );
  INVX3 U963 ( .A(n1234), .Y(n1561) );
  INVX3 U964 ( .A(n1270), .Y(n1606) );
  INVX3 U965 ( .A(n1266), .Y(n1601) );
  INVX3 U966 ( .A(n1250), .Y(n1581) );
  INVX3 U967 ( .A(n1258), .Y(n1591) );
  INVX3 U968 ( .A(n1242), .Y(n1571) );
  INVX3 U969 ( .A(n1125), .Y(n1585) );
  INVX3 U970 ( .A(n1141), .Y(n1605) );
  INVX3 U971 ( .A(n1157), .Y(n1625) );
  INVX3 U972 ( .A(n1137), .Y(n1600) );
  INVX3 U973 ( .A(n1153), .Y(n1620) );
  INVX3 U974 ( .A(n1149), .Y(n1615) );
  INVX3 U975 ( .A(n1129), .Y(n1590) );
  INVX3 U976 ( .A(n1145), .Y(n1610) );
  INVX3 U977 ( .A(n1097), .Y(n1550) );
  INVX3 U978 ( .A(n1109), .Y(n1565) );
  INVX3 U979 ( .A(n1117), .Y(n1575) );
  INVX3 U980 ( .A(n1101), .Y(n1555) );
  INVX3 U981 ( .A(n1105), .Y(n1560) );
  INVX3 U982 ( .A(n1121), .Y(n1580) );
  INVX3 U983 ( .A(n1113), .Y(n1570) );
  INVX3 U984 ( .A(n1028), .Y(n1629) );
  INVX3 U985 ( .A(n1024), .Y(n1624) );
  INVX3 U986 ( .A(n980), .Y(n1569) );
  INVX3 U987 ( .A(n976), .Y(n1564) );
  INVX3 U988 ( .A(n1008), .Y(n1604) );
  INVX3 U989 ( .A(n1012), .Y(n1609) );
  INVX3 U990 ( .A(n1020), .Y(n1619) );
  INVX3 U991 ( .A(n1016), .Y(n1614) );
  INVX1 U992 ( .A(n1048), .Y(n1654) );
  INVX1 U993 ( .A(n1064), .Y(n1674) );
  INVX1 U994 ( .A(n1060), .Y(n1669) );
  INVXL U995 ( .A(n1072), .Y(n1684) );
  INVXL U996 ( .A(n1455), .Y(n1648) );
  INVXL U997 ( .A(n1440), .Y(n1633) );
  INVX1 U998 ( .A(n1445), .Y(n1638) );
  INVXL U999 ( .A(n1465), .Y(n1658) );
  INVX1 U1000 ( .A(n1450), .Y(n1643) );
  INVX1 U1001 ( .A(n1460), .Y(n1653) );
  INVX1 U1002 ( .A(n1475), .Y(n1668) );
  INVX1 U1003 ( .A(n1480), .Y(n1673) );
  INVXL U1004 ( .A(n1490), .Y(n1683) );
  INVX1 U1005 ( .A(n1298), .Y(n1641) );
  INVX1 U1006 ( .A(n1306), .Y(n1651) );
  INVXL U1007 ( .A(n1330), .Y(n1681) );
  INVX1 U1008 ( .A(n1169), .Y(n1640) );
  INVX1 U1009 ( .A(n1177), .Y(n1650) );
  INVXL U1010 ( .A(n1201), .Y(n1680) );
  NAND3BXL U1011 ( .AN(n533), .B(n962), .C(n1544), .Y(n1356) );
  NAND2XL U1012 ( .A(n962), .B(n1543), .Y(n1514) );
  CLKMX2X4 U1013 ( .A(n1332), .B(n1331), .S0(n774), .Y(n1334) );
  MX4XL U1014 ( .A(\block[4][124] ), .B(\block[6][124] ), .C(\block[5][124] ), 
        .D(\block[7][124] ), .S0(n750), .S1(n722), .Y(n1496) );
  NAND2XL U1015 ( .A(mem_rdata[1]), .B(n570), .Y(n971) );
  NAND2XL U1016 ( .A(mem_rdata[14]), .B(n568), .Y(n1023) );
  NAND2XL U1017 ( .A(mem_rdata[53]), .B(n568), .Y(n1180) );
  NAND2X1 U1018 ( .A(mem_rdata[91]), .B(n563), .Y(n1333) );
  NAND2X1 U1019 ( .A(mem_rdata[80]), .B(n567), .Y(n1289) );
  NAND2X1 U1020 ( .A(mem_rdata[81]), .B(n563), .Y(n1293) );
  NAND2X1 U1021 ( .A(mem_rdata[82]), .B(n568), .Y(n1297) );
  NAND2X1 U1022 ( .A(mem_rdata[83]), .B(n559), .Y(n1301) );
  NAND2X1 U1023 ( .A(mem_rdata[85]), .B(n571), .Y(n1309) );
  NAND2X1 U1024 ( .A(mem_rdata[86]), .B(n568), .Y(n1313) );
  NAND2X1 U1025 ( .A(mem_rdata[87]), .B(n564), .Y(n1317) );
  NAND2X1 U1026 ( .A(mem_rdata[88]), .B(n565), .Y(n1321) );
  NAND2X1 U1027 ( .A(mem_rdata[89]), .B(n558), .Y(n1325) );
  NAND2X2 U1028 ( .A(mem_rdata[79]), .B(n568), .Y(n1285) );
  NAND2XL U1029 ( .A(mem_rdata[27]), .B(n568), .Y(n1075) );
  MX4XL U1030 ( .A(\block[4][79] ), .B(\block[6][79] ), .C(\block[5][79] ), 
        .D(\block[7][79] ), .S0(n754), .S1(n716), .Y(n1283) );
  MX4XL U1031 ( .A(\block[4][78] ), .B(\block[6][78] ), .C(\block[5][78] ), 
        .D(\block[7][78] ), .S0(n103), .S1(n715), .Y(n1279) );
  MX4XL U1032 ( .A(\block[0][39] ), .B(\block[2][39] ), .C(\block[1][39] ), 
        .D(\block[3][39] ), .S0(n758), .S1(n732), .Y(n1123) );
  MX4XL U1033 ( .A(\block[0][103] ), .B(\block[2][103] ), .C(\block[1][103] ), 
        .D(\block[3][103] ), .S0(n758), .S1(n718), .Y(n1392) );
  MX4XL U1034 ( .A(\block[4][99] ), .B(\block[6][99] ), .C(\block[5][99] ), 
        .D(\block[7][99] ), .S0(n758), .S1(n718), .Y(n1371) );
  MX4XL U1035 ( .A(\block[0][101] ), .B(\block[2][101] ), .C(\block[1][101] ), 
        .D(\block[3][101] ), .S0(n758), .S1(n718), .Y(n1382) );
  MX4XL U1036 ( .A(\block[4][42] ), .B(\block[6][42] ), .C(\block[5][42] ), 
        .D(\block[7][42] ), .S0(n759), .S1(n733), .Y(n1134) );
  MX4XL U1037 ( .A(\block[4][35] ), .B(\block[6][35] ), .C(\block[5][35] ), 
        .D(\block[7][35] ), .S0(n442), .S1(n732), .Y(n1106) );
  MX4XL U1038 ( .A(\block[0][69] ), .B(\block[2][69] ), .C(\block[1][69] ), 
        .D(\block[3][69] ), .S0(n754), .S1(n714), .Y(n1244) );
  MX4XL U1039 ( .A(\block[4][68] ), .B(\block[6][68] ), .C(\block[5][68] ), 
        .D(\block[7][68] ), .S0(n754), .S1(n714), .Y(n1239) );
  MXI2X1 U1040 ( .A(n1743), .B(n954), .S0(n951), .Y(n1727) );
  MXI2X1 U1041 ( .A(n1742), .B(n954), .S0(n57), .Y(n1726) );
  MXI2X1 U1042 ( .A(n1741), .B(n954), .S0(n58), .Y(n1725) );
  MXI2X1 U1043 ( .A(n1740), .B(n954), .S0(n952), .Y(n1724) );
  MXI2X1 U1044 ( .A(n1739), .B(n954), .S0(n59), .Y(n1723) );
  MXI2X1 U1045 ( .A(n1738), .B(n954), .S0(n63), .Y(n1722) );
  MXI2X1 U1046 ( .A(n1737), .B(n954), .S0(n953), .Y(n1721) );
  MXI2X1 U1047 ( .A(n1736), .B(n954), .S0(n60), .Y(n1720) );
  NAND2XL U1048 ( .A(mem_rdata[105]), .B(n567), .Y(n1403) );
  NAND2XL U1049 ( .A(mem_rdata[92]), .B(n562), .Y(n1337) );
  NAND2XL U1050 ( .A(mem_rdata[118]), .B(n572), .Y(n1468) );
  MX2X1 U1051 ( .A(n998), .B(n997), .S0(n778), .Y(n1000) );
  MX4XL U1052 ( .A(\block[4][8] ), .B(\block[6][8] ), .C(\block[5][8] ), .D(
        \block[7][8] ), .S0(n542), .S1(n727), .Y(n997) );
  MX4XL U1053 ( .A(\block[0][8] ), .B(\block[2][8] ), .C(\block[1][8] ), .D(
        \block[3][8] ), .S0(n444), .S1(n727), .Y(n998) );
  MX2X1 U1054 ( .A(n990), .B(n989), .S0(n778), .Y(n992) );
  MX4XL U1055 ( .A(\block[0][6] ), .B(\block[2][6] ), .C(\block[1][6] ), .D(
        \block[3][6] ), .S0(n444), .S1(n727), .Y(n990) );
  MX4XL U1056 ( .A(\block[4][6] ), .B(\block[6][6] ), .C(\block[5][6] ), .D(
        \block[7][6] ), .S0(n444), .S1(n727), .Y(n989) );
  MX2XL U1057 ( .A(n982), .B(n981), .S0(n778), .Y(n984) );
  MX4XL U1058 ( .A(\block[4][4] ), .B(\block[6][4] ), .C(\block[5][4] ), .D(
        \block[7][4] ), .S0(n444), .S1(n727), .Y(n981) );
  MX4XL U1059 ( .A(\block[0][4] ), .B(\block[2][4] ), .C(\block[1][4] ), .D(
        \block[3][4] ), .S0(n754), .S1(n727), .Y(n982) );
  MX2XL U1060 ( .A(n994), .B(n993), .S0(n778), .Y(n996) );
  MX4XL U1061 ( .A(\block[4][7] ), .B(\block[6][7] ), .C(\block[5][7] ), .D(
        \block[7][7] ), .S0(n754), .S1(n727), .Y(n993) );
  MX4XL U1062 ( .A(\block[4][107] ), .B(\block[6][107] ), .C(\block[5][107] ), 
        .D(\block[7][107] ), .S0(n103), .S1(n719), .Y(n1411) );
  MX4XL U1063 ( .A(\block[0][37] ), .B(\block[2][37] ), .C(\block[1][37] ), 
        .D(\block[3][37] ), .S0(n758), .S1(n732), .Y(n1115) );
  MX4XL U1064 ( .A(\block[4][34] ), .B(\block[6][34] ), .C(\block[5][34] ), 
        .D(\block[7][34] ), .S0(n758), .S1(n732), .Y(n1102) );
  MX4XL U1065 ( .A(\block[4][74] ), .B(\block[6][74] ), .C(\block[5][74] ), 
        .D(\block[7][74] ), .S0(n754), .S1(n715), .Y(n1263) );
  MX4XL U1066 ( .A(\block[4][71] ), .B(\block[6][71] ), .C(\block[5][71] ), 
        .D(\block[7][71] ), .S0(n754), .S1(n714), .Y(n1251) );
  MX4XL U1067 ( .A(\block[0][49] ), .B(\block[2][49] ), .C(\block[1][49] ), 
        .D(\block[3][49] ), .S0(n760), .S1(n734), .Y(n1163) );
  MX2XL U1068 ( .A(n1042), .B(n1041), .S0(n778), .Y(n1044) );
  MX4XL U1069 ( .A(\block[0][19] ), .B(\block[2][19] ), .C(\block[1][19] ), 
        .D(\block[3][19] ), .S0(n755), .S1(n729), .Y(n1042) );
  MX4XL U1070 ( .A(\block[4][19] ), .B(\block[6][19] ), .C(\block[5][19] ), 
        .D(\block[7][19] ), .S0(n755), .S1(n729), .Y(n1041) );
  MX2XL U1071 ( .A(n1038), .B(n1037), .S0(n778), .Y(n1040) );
  MX4XL U1072 ( .A(\block[0][18] ), .B(\block[2][18] ), .C(\block[1][18] ), 
        .D(\block[3][18] ), .S0(n755), .S1(n729), .Y(n1038) );
  MX4XL U1073 ( .A(\block[4][18] ), .B(\block[6][18] ), .C(\block[5][18] ), 
        .D(\block[7][18] ), .S0(n755), .S1(n729), .Y(n1037) );
  MX2XL U1074 ( .A(n1030), .B(n1029), .S0(n778), .Y(n1032) );
  MX4XL U1075 ( .A(\block[0][16] ), .B(\block[2][16] ), .C(\block[1][16] ), 
        .D(\block[3][16] ), .S0(n755), .S1(n729), .Y(n1030) );
  MX4XL U1076 ( .A(\block[4][16] ), .B(\block[6][16] ), .C(\block[5][16] ), 
        .D(\block[7][16] ), .S0(n755), .S1(n729), .Y(n1029) );
  MX2XL U1077 ( .A(n1034), .B(n1033), .S0(n778), .Y(n1036) );
  MX4XL U1078 ( .A(\block[0][17] ), .B(\block[2][17] ), .C(\block[1][17] ), 
        .D(\block[3][17] ), .S0(n755), .S1(n729), .Y(n1034) );
  MX4XL U1079 ( .A(\block[4][17] ), .B(\block[6][17] ), .C(\block[5][17] ), 
        .D(\block[7][17] ), .S0(n755), .S1(n729), .Y(n1033) );
  MX4XL U1080 ( .A(\block[0][85] ), .B(\block[2][85] ), .C(\block[1][85] ), 
        .D(\block[3][85] ), .S0(n754), .S1(n716), .Y(n1308) );
  MX4XL U1081 ( .A(\block[0][121] ), .B(\block[2][121] ), .C(\block[1][121] ), 
        .D(\block[3][121] ), .S0(n542), .S1(n721), .Y(n1482) );
  NAND3BXL U1082 ( .AN(proc_addr[0]), .B(n962), .C(n533), .Y(n1354) );
  CLKBUFX3 U1083 ( .A(n680), .Y(n675) );
  CLKBUFX3 U1084 ( .A(n666), .Y(n674) );
  CLKBUFX3 U1085 ( .A(n666), .Y(n673) );
  CLKBUFX3 U1086 ( .A(n666), .Y(n672) );
  CLKBUFX3 U1087 ( .A(n679), .Y(n671) );
  CLKBUFX3 U1088 ( .A(n679), .Y(n670) );
  CLKBUFX3 U1089 ( .A(n679), .Y(n669) );
  CLKBUFX3 U1090 ( .A(n666), .Y(n668) );
  CLKBUFX3 U1091 ( .A(n666), .Y(n667) );
  CLKBUFX3 U1092 ( .A(n680), .Y(n676) );
  CLKBUFX3 U1093 ( .A(n663), .Y(n659) );
  CLKBUFX3 U1094 ( .A(n650), .Y(n658) );
  CLKBUFX3 U1095 ( .A(n664), .Y(n657) );
  CLKBUFX3 U1096 ( .A(n664), .Y(n656) );
  CLKBUFX3 U1097 ( .A(n664), .Y(n655) );
  CLKBUFX3 U1098 ( .A(n663), .Y(n654) );
  CLKBUFX3 U1099 ( .A(n650), .Y(n653) );
  CLKBUFX3 U1100 ( .A(n664), .Y(n652) );
  CLKBUFX3 U1101 ( .A(n650), .Y(n651) );
  CLKBUFX3 U1102 ( .A(n663), .Y(n660) );
  CLKBUFX3 U1103 ( .A(n710), .Y(n705) );
  CLKBUFX3 U1104 ( .A(n1711), .Y(n704) );
  CLKBUFX3 U1105 ( .A(n1711), .Y(n703) );
  CLKBUFX3 U1106 ( .A(n710), .Y(n702) );
  CLKBUFX3 U1107 ( .A(n710), .Y(n701) );
  CLKBUFX3 U1108 ( .A(n1711), .Y(n700) );
  CLKBUFX3 U1109 ( .A(n1711), .Y(n699) );
  CLKBUFX3 U1110 ( .A(n1711), .Y(n698) );
  CLKBUFX3 U1111 ( .A(n1711), .Y(n697) );
  CLKBUFX3 U1112 ( .A(n709), .Y(n706) );
  CLKBUFX3 U1113 ( .A(n53), .Y(n690) );
  CLKBUFX3 U1114 ( .A(n694), .Y(n689) );
  CLKBUFX3 U1115 ( .A(n694), .Y(n688) );
  CLKBUFX3 U1116 ( .A(n695), .Y(n687) );
  CLKBUFX3 U1117 ( .A(n695), .Y(n686) );
  CLKBUFX3 U1118 ( .A(n696), .Y(n685) );
  CLKBUFX3 U1119 ( .A(n696), .Y(n684) );
  CLKBUFX3 U1120 ( .A(n696), .Y(n683) );
  CLKBUFX3 U1121 ( .A(n696), .Y(n682) );
  CLKBUFX3 U1122 ( .A(n681), .Y(n691) );
  CLKBUFX3 U1123 ( .A(n646), .Y(n641) );
  CLKBUFX3 U1124 ( .A(n647), .Y(n640) );
  CLKBUFX3 U1125 ( .A(n647), .Y(n639) );
  CLKBUFX3 U1126 ( .A(n648), .Y(n638) );
  CLKBUFX3 U1127 ( .A(n648), .Y(n637) );
  CLKBUFX3 U1128 ( .A(n649), .Y(n636) );
  CLKBUFX3 U1129 ( .A(n649), .Y(n635) );
  CLKBUFX3 U1130 ( .A(n649), .Y(n634) );
  CLKBUFX3 U1131 ( .A(n645), .Y(n633) );
  CLKBUFX3 U1132 ( .A(n629), .Y(n622) );
  CLKBUFX3 U1133 ( .A(n629), .Y(n621) );
  CLKBUFX3 U1134 ( .A(n630), .Y(n620) );
  CLKBUFX3 U1135 ( .A(n630), .Y(n619) );
  CLKBUFX3 U1136 ( .A(n631), .Y(n618) );
  CLKBUFX3 U1137 ( .A(n631), .Y(n617) );
  CLKBUFX3 U1138 ( .A(n632), .Y(n616) );
  CLKBUFX3 U1139 ( .A(n632), .Y(n615) );
  CLKBUFX3 U1140 ( .A(n646), .Y(n642) );
  CLKBUFX3 U1141 ( .A(n600), .Y(n610) );
  CLKBUFX3 U1142 ( .A(n601), .Y(n609) );
  CLKBUFX3 U1143 ( .A(n601), .Y(n608) );
  CLKBUFX3 U1144 ( .A(n600), .Y(n607) );
  CLKBUFX3 U1145 ( .A(n600), .Y(n606) );
  CLKBUFX3 U1146 ( .A(n614), .Y(n605) );
  CLKBUFX3 U1147 ( .A(n614), .Y(n604) );
  CLKBUFX3 U1148 ( .A(n600), .Y(n603) );
  CLKBUFX3 U1149 ( .A(n600), .Y(n602) );
  CLKBUFX3 U1150 ( .A(n598), .Y(n594) );
  CLKBUFX3 U1151 ( .A(n598), .Y(n593) );
  CLKBUFX3 U1152 ( .A(n599), .Y(n592) );
  CLKBUFX3 U1153 ( .A(n599), .Y(n591) );
  CLKBUFX3 U1154 ( .A(n586), .Y(n590) );
  CLKBUFX3 U1155 ( .A(n586), .Y(n589) );
  CLKBUFX3 U1156 ( .A(n586), .Y(n588) );
  CLKBUFX3 U1157 ( .A(n586), .Y(n587) );
  CLKBUFX3 U1158 ( .A(n600), .Y(n611) );
  CLKBUFX3 U1159 ( .A(n679), .Y(n678) );
  CLKBUFX3 U1160 ( .A(n664), .Y(n662) );
  CLKBUFX3 U1161 ( .A(n709), .Y(n708) );
  CLKBUFX3 U1162 ( .A(n695), .Y(n693) );
  CLKBUFX3 U1163 ( .A(n645), .Y(n644) );
  CLKBUFX3 U1164 ( .A(n627), .Y(n626) );
  CLKBUFX3 U1165 ( .A(n600), .Y(n613) );
  CLKBUFX3 U1166 ( .A(n584), .Y(n596) );
  CLKBUFX3 U1167 ( .A(n665), .Y(n680) );
  CLKBUFX3 U1168 ( .A(n54), .Y(n664) );
  CLKBUFX3 U1169 ( .A(n54), .Y(n663) );
  CLKBUFX3 U1170 ( .A(n53), .Y(n694) );
  CLKBUFX3 U1171 ( .A(n53), .Y(n695) );
  CLKBUFX3 U1172 ( .A(n665), .Y(n679) );
  CLKBUFX3 U1173 ( .A(n1711), .Y(n709) );
  CLKBUFX3 U1174 ( .A(n61), .Y(n647) );
  CLKBUFX3 U1175 ( .A(n61), .Y(n649) );
  CLKBUFX3 U1176 ( .A(n64), .Y(n629) );
  CLKBUFX3 U1177 ( .A(n64), .Y(n630) );
  CLKBUFX3 U1178 ( .A(n61), .Y(n646) );
  CLKBUFX3 U1179 ( .A(n630), .Y(n628) );
  CLKBUFX3 U1180 ( .A(n601), .Y(n614) );
  CLKBUFX3 U1181 ( .A(n585), .Y(n598) );
  CLKBUFX3 U1182 ( .A(n584), .Y(n597) );
  CLKBUFX3 U1183 ( .A(n61), .Y(n645) );
  CLKBUFX3 U1184 ( .A(n64), .Y(n627) );
  CLKBUFX3 U1185 ( .A(n52), .Y(n665) );
  CLKBUFX3 U1186 ( .A(n56), .Y(n585) );
  CLKBUFX3 U1187 ( .A(n56), .Y(n586) );
  CLKBUFX3 U1188 ( .A(n56), .Y(n584) );
  INVX3 U1189 ( .A(n737), .Y(n731) );
  INVX3 U1190 ( .A(n737), .Y(n730) );
  INVX3 U1191 ( .A(n744), .Y(n722) );
  INVX3 U1192 ( .A(n742), .Y(n712) );
  INVX3 U1193 ( .A(n740), .Y(n717) );
  NOR2X1 U1194 ( .A(n766), .B(n772), .Y(n1745) );
  INVX3 U1195 ( .A(n737), .Y(n732) );
  INVX3 U1196 ( .A(n738), .Y(n727) );
  INVX3 U1197 ( .A(n738), .Y(n729) );
  INVX3 U1198 ( .A(n740), .Y(n718) );
  INVX3 U1199 ( .A(n741), .Y(n714) );
  INVX3 U1200 ( .A(n737), .Y(n719) );
  INVX3 U1201 ( .A(n741), .Y(n715) );
  INVX3 U1202 ( .A(n740), .Y(n720) );
  INVX3 U1203 ( .A(n741), .Y(n716) );
  INVX3 U1204 ( .A(n740), .Y(n721) );
  INVX3 U1205 ( .A(n736), .Y(n733) );
  CLKINVX1 U1206 ( .A(n736), .Y(n735) );
  INVX4 U1207 ( .A(n782), .Y(n775) );
  INVX4 U1208 ( .A(n781), .Y(n777) );
  INVX3 U1209 ( .A(n783), .Y(n773) );
  INVX3 U1210 ( .A(n783), .Y(n774) );
  INVX3 U1211 ( .A(n782), .Y(n776) );
  BUFX8 U1212 ( .A(n70), .Y(n547) );
  NOR2XL U1213 ( .A(n784), .B(n760), .Y(n1746) );
  NOR2XL U1214 ( .A(n784), .B(n766), .Y(n1747) );
  INVX4 U1215 ( .A(n781), .Y(n778) );
  CLKBUFX3 U1216 ( .A(n1356), .Y(n556) );
  CLKBUFX3 U1217 ( .A(n1514), .Y(n574) );
  CLKBUFX3 U1218 ( .A(n1514), .Y(n573) );
  OAI221XL U1219 ( .A0(n1664), .A1(n505), .B0(n1663), .B1(n583), .C0(n1662), 
        .Y(proc_rdata[22]) );
  NAND3BXL U1220 ( .AN(n555), .B(n65), .C(n552), .Y(n1224) );
  BUFX8 U1221 ( .A(n1515), .Y(n577) );
  BUFX8 U1222 ( .A(n1515), .Y(n576) );
  OAI221X1 U1223 ( .A0(n1604), .A1(n505), .B0(n1603), .B1(n582), .C0(n1602), 
        .Y(proc_rdata[10]) );
  OA22X1 U1224 ( .A0(n1601), .A1(n581), .B0(n1600), .B1(n540), .Y(n1602) );
  OA22X1 U1225 ( .A0(n1596), .A1(n581), .B0(n1595), .B1(n540), .Y(n1597) );
  OAI221X1 U1226 ( .A0(n1619), .A1(n505), .B0(n1618), .B1(n583), .C0(n1617), 
        .Y(proc_rdata[13]) );
  OA22X1 U1227 ( .A0(n1616), .A1(n579), .B0(n1615), .B1(n540), .Y(n1617) );
  OAI221X1 U1228 ( .A0(n1614), .A1(n505), .B0(n1613), .B1(n583), .C0(n1612), 
        .Y(proc_rdata[12]) );
  OAI221XL U1229 ( .A0(n1649), .A1(n505), .B0(n1648), .B1(n583), .C0(n1647), 
        .Y(proc_rdata[19]) );
  OAI221XL U1230 ( .A0(n1659), .A1(n505), .B0(n1658), .B1(n583), .C0(n1657), 
        .Y(proc_rdata[21]) );
  OAI221XL U1231 ( .A0(n1644), .A1(n505), .B0(n1643), .B1(n583), .C0(n1642), 
        .Y(proc_rdata[18]) );
  OAI221XL U1232 ( .A0(n1654), .A1(n505), .B0(n1653), .B1(n583), .C0(n1652), 
        .Y(proc_rdata[20]) );
  OAI221XL U1233 ( .A0(n1634), .A1(n505), .B0(n1633), .B1(n583), .C0(n1632), 
        .Y(proc_rdata[16]) );
  OA22X1 U1234 ( .A0(n1671), .A1(n580), .B0(n1670), .B1(n540), .Y(n1672) );
  OA22X1 U1235 ( .A0(n1676), .A1(n580), .B0(n1675), .B1(n540), .Y(n1677) );
  OAI221XL U1236 ( .A0(n1669), .A1(n505), .B0(n1668), .B1(n583), .C0(n1667), 
        .Y(proc_rdata[23]) );
  OAI221XL U1237 ( .A0(n1639), .A1(n505), .B0(n1638), .B1(n583), .C0(n1637), 
        .Y(proc_rdata[17]) );
  BUFX4 U1238 ( .A(n1515), .Y(n578) );
  OAI221XL U1239 ( .A0(n1684), .A1(n505), .B0(n1683), .B1(n583), .C0(n1682), 
        .Y(proc_rdata[26]) );
  CLKBUFX3 U1240 ( .A(n1354), .Y(n552) );
  CLKBUFX3 U1241 ( .A(n1354), .Y(n551) );
  CLKBUFX3 U1242 ( .A(n1356), .Y(n557) );
  CLKBUFX3 U1243 ( .A(n1514), .Y(n575) );
  NAND2BX1 U1244 ( .AN(n949), .B(n955), .Y(n950) );
  NAND4XL U1245 ( .A(n395), .B(n557), .C(n1355), .D(n1354), .Y(n1357) );
  CLKINVX1 U1246 ( .A(n1334), .Y(n1686) );
  CLKINVX1 U1247 ( .A(n996), .Y(n1589) );
  CLKINVX1 U1248 ( .A(n992), .Y(n1584) );
  CLKINVX1 U1249 ( .A(n1000), .Y(n1594) );
  CLKINVX1 U1250 ( .A(n984), .Y(n1574) );
  CLKINVX1 U1251 ( .A(n1044), .Y(n1649) );
  CLKINVX1 U1252 ( .A(n1040), .Y(n1644) );
  CLKINVX1 U1253 ( .A(n1032), .Y(n1634) );
  CLKINVX1 U1254 ( .A(n1036), .Y(n1639) );
  CLKINVX1 U1255 ( .A(n1314), .Y(n1661) );
  CLKINVX1 U1256 ( .A(n1290), .Y(n1631) );
  CLKINVX1 U1257 ( .A(n1322), .Y(n1671) );
  CLKINVX1 U1258 ( .A(n1318), .Y(n1666) );
  CLKINVX1 U1259 ( .A(n1294), .Y(n1636) );
  CLKINVX1 U1260 ( .A(n955), .Y(n962) );
  NAND3BXL U1261 ( .AN(n1544), .B(n962), .C(n533), .Y(n1355) );
  NAND2XL U1262 ( .A(mem_rdata[2]), .B(n568), .Y(n975) );
  NAND2XL U1263 ( .A(mem_rdata[3]), .B(n568), .Y(n979) );
  NAND2XL U1264 ( .A(mem_rdata[4]), .B(n567), .Y(n983) );
  NAND2XL U1265 ( .A(mem_rdata[5]), .B(n570), .Y(n987) );
  NAND2XL U1266 ( .A(mem_rdata[6]), .B(n558), .Y(n991) );
  NAND2XL U1267 ( .A(mem_rdata[8]), .B(n566), .Y(n999) );
  NAND2XL U1268 ( .A(mem_rdata[9]), .B(n565), .Y(n1003) );
  NAND2XL U1269 ( .A(mem_rdata[10]), .B(n562), .Y(n1007) );
  NAND2XL U1270 ( .A(mem_rdata[11]), .B(n568), .Y(n1011) );
  NAND2XL U1271 ( .A(mem_rdata[12]), .B(n561), .Y(n1015) );
  NAND2XL U1272 ( .A(mem_rdata[13]), .B(n563), .Y(n1019) );
  NAND2XL U1273 ( .A(mem_rdata[15]), .B(n571), .Y(n1027) );
  NAND2XL U1274 ( .A(mem_rdata[16]), .B(n571), .Y(n1031) );
  NAND2XL U1275 ( .A(mem_rdata[17]), .B(n568), .Y(n1035) );
  NAND2XL U1276 ( .A(mem_rdata[18]), .B(n558), .Y(n1039) );
  NAND2XL U1277 ( .A(mem_rdata[19]), .B(n564), .Y(n1043) );
  NAND2XL U1278 ( .A(mem_rdata[20]), .B(n569), .Y(n1047) );
  NAND2XL U1279 ( .A(mem_rdata[21]), .B(n559), .Y(n1051) );
  NAND2XL U1280 ( .A(mem_rdata[22]), .B(n563), .Y(n1055) );
  NAND2XL U1281 ( .A(mem_rdata[23]), .B(n566), .Y(n1059) );
  NAND2XL U1282 ( .A(mem_rdata[24]), .B(n566), .Y(n1063) );
  NAND2XL U1283 ( .A(mem_rdata[25]), .B(n571), .Y(n1067) );
  NAND2XL U1284 ( .A(mem_rdata[26]), .B(n569), .Y(n1071) );
  NAND2XL U1285 ( .A(mem_rdata[28]), .B(n565), .Y(n1079) );
  NAND2XL U1286 ( .A(mem_rdata[29]), .B(n569), .Y(n1083) );
  NAND2XL U1287 ( .A(mem_rdata[30]), .B(n562), .Y(n1087) );
  NAND2XL U1288 ( .A(mem_rdata[31]), .B(n558), .Y(n1091) );
  NAND2XL U1289 ( .A(mem_rdata[32]), .B(n560), .Y(n1096) );
  NAND2XL U1290 ( .A(mem_rdata[33]), .B(n568), .Y(n1100) );
  NAND2XL U1291 ( .A(mem_rdata[34]), .B(n559), .Y(n1104) );
  NAND2XL U1292 ( .A(mem_rdata[36]), .B(n566), .Y(n1112) );
  NAND2XL U1293 ( .A(mem_rdata[37]), .B(n568), .Y(n1116) );
  NAND2XL U1294 ( .A(mem_rdata[38]), .B(n568), .Y(n1120) );
  NAND2XL U1295 ( .A(mem_rdata[39]), .B(n565), .Y(n1124) );
  NAND2XL U1296 ( .A(mem_rdata[41]), .B(n564), .Y(n1132) );
  NAND2XL U1297 ( .A(mem_rdata[42]), .B(n558), .Y(n1136) );
  NAND2XL U1298 ( .A(mem_rdata[43]), .B(n568), .Y(n1140) );
  NAND2XL U1299 ( .A(mem_rdata[44]), .B(n564), .Y(n1144) );
  NAND2XL U1300 ( .A(mem_rdata[45]), .B(n568), .Y(n1148) );
  NAND2XL U1301 ( .A(mem_rdata[46]), .B(n572), .Y(n1152) );
  NAND2XL U1302 ( .A(mem_rdata[47]), .B(n564), .Y(n1156) );
  NAND2XL U1303 ( .A(mem_rdata[48]), .B(n569), .Y(n1160) );
  NAND2XL U1304 ( .A(mem_rdata[49]), .B(n560), .Y(n1164) );
  NAND2XL U1305 ( .A(mem_rdata[50]), .B(n565), .Y(n1168) );
  NAND2XL U1306 ( .A(mem_rdata[51]), .B(n566), .Y(n1172) );
  NAND2XL U1307 ( .A(mem_rdata[52]), .B(n568), .Y(n1176) );
  NAND2XL U1308 ( .A(mem_rdata[54]), .B(n568), .Y(n1184) );
  NAND2XL U1309 ( .A(mem_rdata[55]), .B(n561), .Y(n1188) );
  NAND2XL U1310 ( .A(mem_rdata[56]), .B(n572), .Y(n1192) );
  NAND2XL U1311 ( .A(mem_rdata[57]), .B(n558), .Y(n1196) );
  NAND2XL U1312 ( .A(mem_rdata[58]), .B(n564), .Y(n1200) );
  NAND2XL U1313 ( .A(mem_rdata[59]), .B(n568), .Y(n1204) );
  NAND2XL U1314 ( .A(mem_rdata[60]), .B(n560), .Y(n1208) );
  NAND2XL U1315 ( .A(mem_rdata[61]), .B(n568), .Y(n1212) );
  NAND2XL U1316 ( .A(mem_rdata[62]), .B(n570), .Y(n1216) );
  NAND2XL U1317 ( .A(mem_rdata[64]), .B(n561), .Y(n1225) );
  NAND2XL U1318 ( .A(mem_rdata[65]), .B(n569), .Y(n1229) );
  NAND2XL U1319 ( .A(mem_rdata[67]), .B(n562), .Y(n1237) );
  NAND2XL U1320 ( .A(mem_rdata[68]), .B(n568), .Y(n1241) );
  NAND2XL U1321 ( .A(mem_rdata[69]), .B(n569), .Y(n1245) );
  NAND2XL U1322 ( .A(mem_rdata[70]), .B(n568), .Y(n1249) );
  NAND2XL U1323 ( .A(mem_rdata[71]), .B(n570), .Y(n1253) );
  NAND2XL U1324 ( .A(mem_rdata[72]), .B(n568), .Y(n1257) );
  NAND2XL U1325 ( .A(mem_rdata[73]), .B(n559), .Y(n1261) );
  NAND2XL U1326 ( .A(mem_rdata[74]), .B(n564), .Y(n1265) );
  NAND2XL U1327 ( .A(mem_rdata[75]), .B(n568), .Y(n1269) );
  NAND2XL U1328 ( .A(mem_rdata[76]), .B(n564), .Y(n1273) );
  NAND2XL U1329 ( .A(mem_rdata[77]), .B(n565), .Y(n1277) );
  NAND2XL U1330 ( .A(mem_rdata[78]), .B(n560), .Y(n1281) );
  NAND2XL U1331 ( .A(mem_rdata[93]), .B(n561), .Y(n1341) );
  NAND2XL U1332 ( .A(mem_rdata[94]), .B(n571), .Y(n1345) );
  NAND2XL U1333 ( .A(mem_rdata[95]), .B(n569), .Y(n1349) );
  MX4XL U1334 ( .A(blockdirty[4]), .B(blockdirty[6]), .C(blockdirty[5]), .D(
        blockdirty[7]), .S0(n444), .S1(n724), .Y(n806) );
  NAND2XL U1335 ( .A(mem_rdata[96]), .B(n568), .Y(n1358) );
  NAND2XL U1336 ( .A(mem_rdata[97]), .B(n568), .Y(n1363) );
  NAND2XL U1337 ( .A(mem_rdata[98]), .B(n560), .Y(n1368) );
  NAND2XL U1338 ( .A(mem_rdata[99]), .B(n568), .Y(n1373) );
  NAND2XL U1339 ( .A(mem_rdata[100]), .B(n567), .Y(n1378) );
  NAND2XL U1340 ( .A(mem_rdata[101]), .B(n561), .Y(n1383) );
  NAND2XL U1341 ( .A(mem_rdata[102]), .B(n568), .Y(n1388) );
  NAND2XL U1342 ( .A(mem_rdata[103]), .B(n570), .Y(n1393) );
  NAND2XL U1343 ( .A(mem_rdata[104]), .B(n569), .Y(n1398) );
  NAND2XL U1344 ( .A(mem_rdata[106]), .B(n567), .Y(n1408) );
  NAND2XL U1345 ( .A(mem_rdata[107]), .B(n559), .Y(n1413) );
  NAND2XL U1346 ( .A(mem_rdata[108]), .B(n563), .Y(n1418) );
  NAND2XL U1347 ( .A(mem_rdata[109]), .B(n562), .Y(n1423) );
  NAND2XL U1348 ( .A(mem_rdata[110]), .B(n563), .Y(n1428) );
  NAND2XL U1349 ( .A(mem_rdata[111]), .B(n567), .Y(n1433) );
  NAND2XL U1350 ( .A(mem_rdata[112]), .B(n562), .Y(n1438) );
  NAND2XL U1351 ( .A(mem_rdata[113]), .B(n561), .Y(n1443) );
  NAND2XL U1352 ( .A(mem_rdata[114]), .B(n572), .Y(n1448) );
  NAND2XL U1353 ( .A(mem_rdata[115]), .B(n568), .Y(n1453) );
  NAND2XL U1354 ( .A(mem_rdata[116]), .B(n561), .Y(n1458) );
  NAND2XL U1355 ( .A(mem_rdata[117]), .B(n565), .Y(n1463) );
  NAND2XL U1356 ( .A(mem_rdata[119]), .B(n572), .Y(n1473) );
  NAND2XL U1357 ( .A(mem_rdata[120]), .B(n571), .Y(n1478) );
  NAND2XL U1358 ( .A(mem_rdata[121]), .B(n565), .Y(n1483) );
  NAND2XL U1359 ( .A(mem_rdata[122]), .B(n565), .Y(n1488) );
  NAND2XL U1360 ( .A(mem_rdata[123]), .B(n568), .Y(n1493) );
  NAND2XL U1361 ( .A(mem_rdata[124]), .B(n562), .Y(n1498) );
  NAND2XL U1362 ( .A(mem_rdata[125]), .B(n562), .Y(n1501) );
  NAND2XL U1363 ( .A(mem_rdata[126]), .B(n568), .Y(n1506) );
  NAND2XL U1364 ( .A(mem_rdata[127]), .B(n568), .Y(n1512) );
  MX4XL U1365 ( .A(\block[4][127] ), .B(\block[6][127] ), .C(\block[5][127] ), 
        .D(\block[7][127] ), .S0(n750), .S1(n734), .Y(n1509) );
  MX4XL U1366 ( .A(\block[0][127] ), .B(\block[2][127] ), .C(\block[1][127] ), 
        .D(\block[3][127] ), .S0(n441), .S1(n722), .Y(n1510) );
  MX4X1 U1367 ( .A(\block[4][95] ), .B(\block[6][95] ), .C(\block[5][95] ), 
        .D(\block[7][95] ), .S0(n749), .S1(n734), .Y(n1347) );
  CLKMX2X2 U1368 ( .A(n1344), .B(n1343), .S0(n774), .Y(n1346) );
  MX2XL U1369 ( .A(n937), .B(n936), .S0(n571), .Y(n938) );
  MX2XL U1370 ( .A(n922), .B(n921), .S0(n566), .Y(n923) );
  CLKMX2X2 U1371 ( .A(n416), .B(n104), .S0(n568), .Y(n901) );
  INVXL U1372 ( .A(n1528), .Y(n909) );
  MX2XL U1373 ( .A(n885), .B(n884), .S0(n563), .Y(n886) );
  MX2XL U1374 ( .A(n917), .B(n916), .S0(n571), .Y(n918) );
  INVXL U1375 ( .A(n113), .Y(n917) );
  MX2XL U1376 ( .A(n931), .B(n930), .S0(n566), .Y(n932) );
  INVXL U1377 ( .A(n1533), .Y(n931) );
  MX2XL U1378 ( .A(n2), .B(n928), .S0(n559), .Y(n929) );
  INVXL U1379 ( .A(proc_addr[27]), .Y(n928) );
  MX2XL U1380 ( .A(n934), .B(n933), .S0(n569), .Y(n935) );
  INVXL U1381 ( .A(n1534), .Y(n934) );
  MX2XL U1382 ( .A(n940), .B(n939), .S0(n559), .Y(n941) );
  MX2XL U1383 ( .A(n906), .B(n905), .S0(n571), .Y(n907) );
  MX2XL U1384 ( .A(n896), .B(n895), .S0(n571), .Y(n897) );
  INVXL U1385 ( .A(n1524), .Y(n896) );
  MX2XL U1386 ( .A(n899), .B(n898), .S0(n569), .Y(n900) );
  INVXL U1387 ( .A(n1525), .Y(n899) );
  MX2XL U1388 ( .A(n903), .B(n902), .S0(n569), .Y(n904) );
  INVXL U1389 ( .A(n430), .Y(n903) );
  MX2XL U1390 ( .A(n889), .B(n888), .S0(n560), .Y(n890) );
  MX2XL U1391 ( .A(n943), .B(n942), .S0(n567), .Y(n944) );
  AO21XL U1392 ( .A0(mem_ready), .A1(n966), .B0(n447), .Y(n799) );
  MXI2X1 U1393 ( .A(n1735), .B(n803), .S0(n951), .Y(n1719) );
  MXI2X1 U1394 ( .A(n1734), .B(n803), .S0(n57), .Y(n1718) );
  MXI2X1 U1395 ( .A(n1733), .B(n803), .S0(n58), .Y(n1717) );
  MXI2X1 U1396 ( .A(n1732), .B(n803), .S0(n952), .Y(n1716) );
  MXI2X1 U1397 ( .A(n1731), .B(n803), .S0(n59), .Y(n1715) );
  MXI2X1 U1398 ( .A(n1730), .B(n803), .S0(n63), .Y(n1714) );
  MXI2X1 U1399 ( .A(n1729), .B(n803), .S0(n953), .Y(n1713) );
  MXI2X1 U1400 ( .A(n1728), .B(n803), .S0(n60), .Y(n1712) );
  MX2XL U1401 ( .A(n1462), .B(n1461), .S0(n772), .Y(n1465) );
  MX4X1 U1402 ( .A(\block[4][117] ), .B(\block[6][117] ), .C(\block[5][117] ), 
        .D(\block[7][117] ), .S0(n759), .S1(n721), .Y(n1461) );
  MX2XL U1403 ( .A(n1467), .B(n1466), .S0(n772), .Y(n1470) );
  MX4X1 U1404 ( .A(\block[0][118] ), .B(\block[2][118] ), .C(\block[1][118] ), 
        .D(\block[3][118] ), .S0(n759), .S1(n721), .Y(n1467) );
  MX4X1 U1405 ( .A(\block[4][118] ), .B(\block[6][118] ), .C(\block[5][118] ), 
        .D(\block[7][118] ), .S0(n759), .S1(n721), .Y(n1466) );
  MX2XL U1406 ( .A(n1487), .B(n1486), .S0(n772), .Y(n1490) );
  MX4XL U1407 ( .A(\block[0][122] ), .B(\block[2][122] ), .C(\block[1][122] ), 
        .D(\block[3][122] ), .S0(n760), .S1(n722), .Y(n1487) );
  MX4XL U1408 ( .A(\block[4][122] ), .B(\block[6][122] ), .C(\block[5][122] ), 
        .D(\block[7][122] ), .S0(n750), .S1(n722), .Y(n1486) );
  MX2XL U1409 ( .A(n1457), .B(n1456), .S0(n772), .Y(n1460) );
  MX4X1 U1410 ( .A(\block[4][116] ), .B(\block[6][116] ), .C(\block[5][116] ), 
        .D(\block[7][116] ), .S0(n759), .S1(n721), .Y(n1456) );
  MX4X1 U1411 ( .A(\block[0][116] ), .B(\block[2][116] ), .C(\block[1][116] ), 
        .D(\block[3][116] ), .S0(n542), .S1(n721), .Y(n1457) );
  MX2XL U1412 ( .A(n1447), .B(n1446), .S0(n772), .Y(n1450) );
  MX4X1 U1413 ( .A(\block[4][114] ), .B(\block[6][114] ), .C(\block[5][114] ), 
        .D(\block[7][114] ), .S0(n758), .S1(n720), .Y(n1446) );
  MX2XL U1414 ( .A(n1477), .B(n1476), .S0(n772), .Y(n1480) );
  MX4X1 U1415 ( .A(\block[0][120] ), .B(\block[2][120] ), .C(\block[1][120] ), 
        .D(\block[3][120] ), .S0(n754), .S1(n721), .Y(n1477) );
  MX4X1 U1416 ( .A(\block[4][120] ), .B(\block[6][120] ), .C(\block[5][120] ), 
        .D(\block[7][120] ), .S0(n754), .S1(n721), .Y(n1476) );
  MX2XL U1417 ( .A(n1482), .B(n1481), .S0(n772), .Y(n1485) );
  MX4XL U1418 ( .A(\block[4][121] ), .B(\block[6][121] ), .C(\block[5][121] ), 
        .D(\block[7][121] ), .S0(n749), .S1(n722), .Y(n1481) );
  MX2XL U1419 ( .A(n1472), .B(n1471), .S0(n772), .Y(n1475) );
  MX4X1 U1420 ( .A(\block[0][119] ), .B(\block[2][119] ), .C(\block[1][119] ), 
        .D(\block[3][119] ), .S0(n754), .S1(n721), .Y(n1472) );
  MX2XL U1421 ( .A(n1095), .B(n1094), .S0(n777), .Y(n1097) );
  MX4XL U1422 ( .A(\block[4][32] ), .B(\block[6][32] ), .C(\block[5][32] ), 
        .D(\block[7][32] ), .S0(n757), .S1(n732), .Y(n1094) );
  MX4XL U1423 ( .A(\block[0][32] ), .B(\block[2][32] ), .C(\block[1][32] ), 
        .D(\block[3][32] ), .S0(n757), .S1(n732), .Y(n1095) );
  MX2XL U1424 ( .A(n1223), .B(n1222), .S0(n775), .Y(n1226) );
  MX4XL U1425 ( .A(\block[0][64] ), .B(\block[2][64] ), .C(\block[1][64] ), 
        .D(\block[3][64] ), .S0(n747), .S1(n713), .Y(n1223) );
  MX4XL U1426 ( .A(\block[4][64] ), .B(\block[6][64] ), .C(\block[5][64] ), 
        .D(\block[7][64] ), .S0(n747), .S1(n713), .Y(n1222) );
  MX2XL U1427 ( .A(n1353), .B(n1352), .S0(n774), .Y(n1360) );
  MX4XL U1428 ( .A(\block[4][96] ), .B(\block[6][96] ), .C(\block[5][96] ), 
        .D(\block[7][96] ), .S0(n748), .S1(n735), .Y(n1352) );
  MX4XL U1429 ( .A(\block[0][96] ), .B(\block[2][96] ), .C(\block[1][96] ), 
        .D(\block[3][96] ), .S0(n749), .S1(n735), .Y(n1353) );
  MX2XL U1430 ( .A(n957), .B(n956), .S0(n779), .Y(n968) );
  MX4XL U1431 ( .A(\block[4][0] ), .B(\block[6][0] ), .C(\block[5][0] ), .D(
        \block[7][0] ), .S0(n754), .S1(n544), .Y(n956) );
  MX4XL U1432 ( .A(\block[0][0] ), .B(\block[2][0] ), .C(\block[1][0] ), .D(
        \block[3][0] ), .S0(n444), .S1(n544), .Y(n957) );
  MX2XL U1433 ( .A(n1123), .B(n1122), .S0(n776), .Y(n1125) );
  MX2XL U1434 ( .A(n1107), .B(n1106), .S0(n777), .Y(n1109) );
  MX2XL U1435 ( .A(n1236), .B(n1235), .S0(n775), .Y(n1238) );
  MX4XL U1436 ( .A(\block[0][67] ), .B(\block[2][67] ), .C(\block[1][67] ), 
        .D(\block[3][67] ), .S0(n747), .S1(n713), .Y(n1236) );
  MX4XL U1437 ( .A(\block[4][67] ), .B(\block[6][67] ), .C(\block[5][67] ), 
        .D(\block[7][67] ), .S0(n747), .S1(n714), .Y(n1235) );
  MX2XL U1438 ( .A(n1252), .B(n1251), .S0(n775), .Y(n1254) );
  MX2XL U1439 ( .A(n1392), .B(n1391), .S0(n773), .Y(n1395) );
  MX2XL U1440 ( .A(n1115), .B(n1114), .S0(n777), .Y(n1117) );
  MX2XL U1441 ( .A(n1372), .B(n1371), .S0(n773), .Y(n1375) );
  MX2XL U1442 ( .A(n1244), .B(n1243), .S0(n775), .Y(n1246) );
  MX2XL U1443 ( .A(n1382), .B(n1381), .S0(n773), .Y(n1385) );
  CLKMX2X2 U1444 ( .A(n978), .B(n977), .S0(n778), .Y(n980) );
  MX4XL U1445 ( .A(\block[0][3] ), .B(\block[2][3] ), .C(\block[1][3] ), .D(
        \block[3][3] ), .S0(n755), .S1(n727), .Y(n978) );
  MX4XL U1446 ( .A(\block[4][3] ), .B(\block[6][3] ), .C(\block[5][3] ), .D(
        \block[7][3] ), .S0(n749), .S1(n727), .Y(n977) );
  MX2XL U1447 ( .A(n1099), .B(n1098), .S0(n777), .Y(n1101) );
  MX4XL U1448 ( .A(\block[0][33] ), .B(\block[2][33] ), .C(\block[1][33] ), 
        .D(\block[3][33] ), .S0(n757), .S1(n731), .Y(n1099) );
  MX2XL U1449 ( .A(n1228), .B(n1227), .S0(n775), .Y(n1230) );
  MX4XL U1450 ( .A(\block[0][65] ), .B(\block[2][65] ), .C(\block[1][65] ), 
        .D(\block[3][65] ), .S0(n747), .S1(n713), .Y(n1228) );
  MX4XL U1451 ( .A(\block[4][65] ), .B(\block[6][65] ), .C(\block[5][65] ), 
        .D(\block[7][65] ), .S0(n747), .S1(n713), .Y(n1227) );
  MX2XL U1452 ( .A(n1103), .B(n1102), .S0(n777), .Y(n1105) );
  MX2XL U1453 ( .A(n1232), .B(n1231), .S0(n775), .Y(n1234) );
  MX4XL U1454 ( .A(\block[0][66] ), .B(\block[2][66] ), .C(\block[1][66] ), 
        .D(\block[3][66] ), .S0(n747), .S1(n713), .Y(n1232) );
  MX4XL U1455 ( .A(\block[4][66] ), .B(\block[6][66] ), .C(\block[5][66] ), 
        .D(\block[7][66] ), .S0(n747), .S1(n713), .Y(n1231) );
  MX2XL U1456 ( .A(n1362), .B(n1361), .S0(n773), .Y(n1365) );
  MX4XL U1457 ( .A(\block[4][97] ), .B(\block[6][97] ), .C(\block[5][97] ), 
        .D(\block[7][97] ), .S0(n542), .S1(n718), .Y(n1361) );
  MX4XL U1458 ( .A(\block[0][97] ), .B(\block[2][97] ), .C(\block[1][97] ), 
        .D(\block[3][97] ), .S0(n758), .S1(n721), .Y(n1362) );
  MX2XL U1459 ( .A(n1139), .B(n1138), .S0(n776), .Y(n1141) );
  MX2XL U1460 ( .A(n1367), .B(n1366), .S0(n773), .Y(n1370) );
  MX4XL U1461 ( .A(\block[0][98] ), .B(\block[2][98] ), .C(\block[1][98] ), 
        .D(\block[3][98] ), .S0(n542), .S1(n718), .Y(n1367) );
  MX4XL U1462 ( .A(\block[4][1] ), .B(\block[6][1] ), .C(\block[5][1] ), .D(
        \block[7][1] ), .S0(n754), .S1(n544), .Y(n969) );
  MX4XL U1463 ( .A(\block[0][1] ), .B(\block[2][1] ), .C(\block[1][1] ), .D(
        \block[3][1] ), .S0(n746), .S1(n544), .Y(n970) );
  MX2XL U1464 ( .A(n1268), .B(n1267), .S0(n775), .Y(n1270) );
  MX2XL U1465 ( .A(n1155), .B(n1154), .S0(n776), .Y(n1157) );
  MX2XL U1466 ( .A(n1284), .B(n1283), .S0(n774), .Y(n1286) );
  MX2XL U1467 ( .A(n1412), .B(n1411), .S0(n773), .Y(n1415) );
  CLKMX2X2 U1468 ( .A(n974), .B(n973), .S0(n778), .Y(n976) );
  MX4XL U1469 ( .A(\block[0][2] ), .B(\block[2][2] ), .C(\block[1][2] ), .D(
        \block[3][2] ), .S0(n444), .S1(n544), .Y(n974) );
  MX4XL U1470 ( .A(\block[4][2] ), .B(\block[6][2] ), .C(\block[5][2] ), .D(
        \block[7][2] ), .S0(n444), .S1(n544), .Y(n973) );
  CLKMX2X2 U1471 ( .A(n1010), .B(n1009), .S0(n778), .Y(n1012) );
  MX4XL U1472 ( .A(\block[0][11] ), .B(\block[2][11] ), .C(\block[1][11] ), 
        .D(\block[3][11] ), .S0(n754), .S1(n728), .Y(n1010) );
  MX4XL U1473 ( .A(\block[4][11] ), .B(\block[6][11] ), .C(\block[5][11] ), 
        .D(\block[7][11] ), .S0(n444), .S1(n728), .Y(n1009) );
  MX2XL U1474 ( .A(n1432), .B(n1431), .S0(n773), .Y(n1435) );
  MX2X1 U1475 ( .A(n1026), .B(n1025), .S0(n778), .Y(n1028) );
  MX4XL U1476 ( .A(\block[0][15] ), .B(\block[2][15] ), .C(\block[1][15] ), 
        .D(\block[3][15] ), .S0(n754), .S1(n728), .Y(n1026) );
  MX4X1 U1477 ( .A(\block[4][15] ), .B(\block[6][15] ), .C(\block[5][15] ), 
        .D(\block[7][15] ), .S0(n755), .S1(n729), .Y(n1025) );
  MX2XL U1478 ( .A(n1151), .B(n1150), .S0(n776), .Y(n1153) );
  MX2XL U1479 ( .A(n1135), .B(n1134), .S0(n776), .Y(n1137) );
  MX2XL U1480 ( .A(n1280), .B(n1279), .S0(n774), .Y(n1282) );
  MX2XL U1481 ( .A(n1264), .B(n1263), .S0(n775), .Y(n1266) );
  MX2XL U1482 ( .A(n1407), .B(n1406), .S0(n773), .Y(n1410) );
  MX2XL U1483 ( .A(n1427), .B(n1426), .S0(n773), .Y(n1430) );
  MX2XL U1484 ( .A(n1119), .B(n1118), .S0(n777), .Y(n1121) );
  MX4X1 U1485 ( .A(\block[4][38] ), .B(\block[6][38] ), .C(\block[5][38] ), 
        .D(\block[7][38] ), .S0(n758), .S1(n733), .Y(n1118) );
  MX4X1 U1486 ( .A(\block[0][38] ), .B(\block[2][38] ), .C(\block[1][38] ), 
        .D(\block[3][38] ), .S0(n758), .S1(n733), .Y(n1119) );
  MX2X1 U1487 ( .A(n1006), .B(n1005), .S0(n778), .Y(n1008) );
  MX4XL U1488 ( .A(\block[0][10] ), .B(\block[2][10] ), .C(\block[1][10] ), 
        .D(\block[3][10] ), .S0(n754), .S1(n728), .Y(n1006) );
  MX4XL U1489 ( .A(\block[4][10] ), .B(\block[6][10] ), .C(\block[5][10] ), 
        .D(\block[7][10] ), .S0(n444), .S1(n728), .Y(n1005) );
  MX2X1 U1490 ( .A(n1022), .B(n1021), .S0(n778), .Y(n1024) );
  MX4XL U1491 ( .A(\block[0][14] ), .B(\block[2][14] ), .C(\block[1][14] ), 
        .D(\block[3][14] ), .S0(n444), .S1(n729), .Y(n1022) );
  MX4XL U1492 ( .A(\block[4][14] ), .B(\block[6][14] ), .C(\block[5][14] ), 
        .D(\block[7][14] ), .S0(n748), .S1(n729), .Y(n1021) );
  MX2XL U1493 ( .A(n1248), .B(n1247), .S0(n775), .Y(n1250) );
  MX4X1 U1494 ( .A(\block[4][70] ), .B(\block[6][70] ), .C(\block[5][70] ), 
        .D(\block[7][70] ), .S0(n754), .S1(n714), .Y(n1247) );
  MX4X1 U1495 ( .A(\block[0][70] ), .B(\block[2][70] ), .C(\block[1][70] ), 
        .D(\block[3][70] ), .S0(n754), .S1(n714), .Y(n1248) );
  MX2XL U1496 ( .A(n1387), .B(n1386), .S0(n773), .Y(n1390) );
  MX4X1 U1497 ( .A(\block[4][102] ), .B(\block[6][102] ), .C(\block[5][102] ), 
        .D(\block[7][102] ), .S0(n747), .S1(n718), .Y(n1386) );
  MX4X1 U1498 ( .A(\block[0][102] ), .B(\block[2][102] ), .C(\block[1][102] ), 
        .D(\block[3][102] ), .S0(n758), .S1(n718), .Y(n1387) );
  MX2XL U1499 ( .A(n1131), .B(n1130), .S0(n776), .Y(n1133) );
  MX4X1 U1500 ( .A(\block[4][41] ), .B(\block[6][41] ), .C(\block[5][41] ), 
        .D(\block[7][41] ), .S0(n759), .S1(n733), .Y(n1130) );
  MX4X1 U1501 ( .A(\block[0][41] ), .B(\block[2][41] ), .C(\block[1][41] ), 
        .D(\block[3][41] ), .S0(n759), .S1(n733), .Y(n1131) );
  MX2XL U1502 ( .A(n1260), .B(n1259), .S0(n775), .Y(n1262) );
  MX4X1 U1503 ( .A(\block[0][73] ), .B(\block[2][73] ), .C(\block[1][73] ), 
        .D(\block[3][73] ), .S0(n754), .S1(n714), .Y(n1260) );
  MX4X1 U1504 ( .A(\block[4][73] ), .B(\block[6][73] ), .C(\block[5][73] ), 
        .D(\block[7][73] ), .S0(n754), .S1(n715), .Y(n1259) );
  MX2XL U1505 ( .A(n1147), .B(n1146), .S0(n776), .Y(n1149) );
  MX4X1 U1506 ( .A(\block[0][45] ), .B(\block[2][45] ), .C(\block[1][45] ), 
        .D(\block[3][45] ), .S0(n759), .S1(n733), .Y(n1147) );
  MX4X1 U1507 ( .A(\block[4][45] ), .B(\block[6][45] ), .C(\block[5][45] ), 
        .D(\block[7][45] ), .S0(n760), .S1(n734), .Y(n1146) );
  MX2XL U1508 ( .A(n1402), .B(n1401), .S0(n773), .Y(n1405) );
  MX2XL U1509 ( .A(n1276), .B(n1275), .S0(n774), .Y(n1278) );
  MX4X1 U1510 ( .A(\block[0][77] ), .B(\block[2][77] ), .C(\block[1][77] ), 
        .D(\block[3][77] ), .S0(n754), .S1(n715), .Y(n1276) );
  MX4X1 U1511 ( .A(\block[4][77] ), .B(\block[6][77] ), .C(\block[5][77] ), 
        .D(\block[7][77] ), .S0(n754), .S1(n715), .Y(n1275) );
  CLKMX2X2 U1512 ( .A(n1002), .B(n1001), .S0(n778), .Y(n1004) );
  MX4XL U1513 ( .A(\block[4][9] ), .B(\block[6][9] ), .C(\block[5][9] ), .D(
        \block[7][9] ), .S0(n754), .S1(n728), .Y(n1001) );
  MX4XL U1514 ( .A(\block[0][9] ), .B(\block[2][9] ), .C(\block[1][9] ), .D(
        \block[3][9] ), .S0(n444), .S1(n728), .Y(n1002) );
  MX2XL U1515 ( .A(n1422), .B(n1421), .S0(n773), .Y(n1425) );
  MX4X1 U1516 ( .A(\block[0][109] ), .B(\block[2][109] ), .C(\block[1][109] ), 
        .D(\block[3][109] ), .S0(n759), .S1(n719), .Y(n1422) );
  CLKMX2X2 U1517 ( .A(n1018), .B(n1017), .S0(n778), .Y(n1020) );
  MX4XL U1518 ( .A(\block[0][13] ), .B(\block[2][13] ), .C(\block[1][13] ), 
        .D(\block[3][13] ), .S0(n755), .S1(n728), .Y(n1018) );
  MX4XL U1519 ( .A(\block[4][13] ), .B(\block[6][13] ), .C(\block[5][13] ), 
        .D(\block[7][13] ), .S0(n444), .S1(n728), .Y(n1017) );
  MX2XL U1520 ( .A(n1127), .B(n1126), .S0(n776), .Y(n1129) );
  MX4X1 U1521 ( .A(\block[4][40] ), .B(\block[6][40] ), .C(\block[5][40] ), 
        .D(\block[7][40] ), .S0(n759), .S1(n733), .Y(n1126) );
  MX4X1 U1522 ( .A(\block[0][40] ), .B(\block[2][40] ), .C(\block[1][40] ), 
        .D(\block[3][40] ), .S0(n759), .S1(n733), .Y(n1127) );
  MX2XL U1523 ( .A(n1256), .B(n1255), .S0(n775), .Y(n1258) );
  MX4X1 U1524 ( .A(\block[4][72] ), .B(\block[6][72] ), .C(\block[5][72] ), 
        .D(\block[7][72] ), .S0(n754), .S1(n714), .Y(n1255) );
  MX4X1 U1525 ( .A(\block[0][72] ), .B(\block[2][72] ), .C(\block[1][72] ), 
        .D(\block[3][72] ), .S0(n754), .S1(n714), .Y(n1256) );
  MX2XL U1526 ( .A(n1397), .B(n1396), .S0(n773), .Y(n1400) );
  MX4X1 U1527 ( .A(\block[0][104] ), .B(\block[2][104] ), .C(\block[1][104] ), 
        .D(\block[3][104] ), .S0(n758), .S1(n719), .Y(n1397) );
  MX2XL U1528 ( .A(n1111), .B(n1110), .S0(n777), .Y(n1113) );
  MX4X1 U1529 ( .A(\block[4][36] ), .B(\block[6][36] ), .C(\block[5][36] ), 
        .D(\block[7][36] ), .S0(n758), .S1(n732), .Y(n1110) );
  MX4X1 U1530 ( .A(\block[0][36] ), .B(\block[2][36] ), .C(\block[1][36] ), 
        .D(\block[3][36] ), .S0(n758), .S1(n732), .Y(n1111) );
  MX2XL U1531 ( .A(n1143), .B(n1142), .S0(n776), .Y(n1145) );
  MX4X1 U1532 ( .A(\block[4][44] ), .B(\block[6][44] ), .C(\block[5][44] ), 
        .D(\block[7][44] ), .S0(n759), .S1(n734), .Y(n1142) );
  MX4X1 U1533 ( .A(\block[0][44] ), .B(\block[2][44] ), .C(\block[1][44] ), 
        .D(\block[3][44] ), .S0(n759), .S1(n734), .Y(n1143) );
  MX2XL U1534 ( .A(n1240), .B(n1239), .S0(n775), .Y(n1242) );
  MX4XL U1535 ( .A(\block[0][68] ), .B(\block[2][68] ), .C(\block[1][68] ), 
        .D(\block[3][68] ), .S0(n747), .S1(n714), .Y(n1240) );
  MX2XL U1536 ( .A(n1377), .B(n1376), .S0(n773), .Y(n1380) );
  MX4X1 U1537 ( .A(\block[4][100] ), .B(\block[6][100] ), .C(\block[5][100] ), 
        .D(\block[7][100] ), .S0(n758), .S1(n718), .Y(n1376) );
  MX4X1 U1538 ( .A(\block[0][100] ), .B(\block[2][100] ), .C(\block[1][100] ), 
        .D(\block[3][100] ), .S0(n747), .S1(n718), .Y(n1377) );
  MX2XL U1539 ( .A(n1272), .B(n1271), .S0(n774), .Y(n1274) );
  MX4X1 U1540 ( .A(\block[4][76] ), .B(\block[6][76] ), .C(\block[5][76] ), 
        .D(\block[7][76] ), .S0(n749), .S1(n715), .Y(n1271) );
  MX4X1 U1541 ( .A(\block[0][76] ), .B(\block[2][76] ), .C(\block[1][76] ), 
        .D(\block[3][76] ), .S0(n754), .S1(n715), .Y(n1272) );
  MX2XL U1542 ( .A(n1417), .B(n1416), .S0(n773), .Y(n1420) );
  CLKMX2X2 U1543 ( .A(n1014), .B(n1013), .S0(n778), .Y(n1016) );
  MX4XL U1544 ( .A(\block[0][12] ), .B(\block[2][12] ), .C(\block[1][12] ), 
        .D(\block[3][12] ), .S0(n754), .S1(n728), .Y(n1014) );
  MX4XL U1545 ( .A(\block[4][12] ), .B(\block[6][12] ), .C(\block[5][12] ), 
        .D(\block[7][12] ), .S0(n444), .S1(n728), .Y(n1013) );
  MX2XL U1546 ( .A(n1179), .B(n1178), .S0(n776), .Y(n1181) );
  MX4XL U1547 ( .A(\block[0][53] ), .B(\block[2][53] ), .C(\block[1][53] ), 
        .D(\block[3][53] ), .S0(n758), .S1(n711), .Y(n1179) );
  MX4XL U1548 ( .A(\block[4][53] ), .B(\block[6][53] ), .C(\block[5][53] ), 
        .D(\block[7][53] ), .S0(n747), .S1(n711), .Y(n1178) );
  MX2XL U1549 ( .A(n1171), .B(n1170), .S0(n776), .Y(n1173) );
  MX4XL U1550 ( .A(\block[0][51] ), .B(\block[2][51] ), .C(\block[1][51] ), 
        .D(\block[3][51] ), .S0(n747), .S1(n711), .Y(n1171) );
  MX4XL U1551 ( .A(\block[4][51] ), .B(\block[6][51] ), .C(\block[5][51] ), 
        .D(\block[7][51] ), .S0(n747), .S1(n711), .Y(n1170) );
  MX2XL U1552 ( .A(n1308), .B(n1307), .S0(n774), .Y(n1310) );
  MX4XL U1553 ( .A(\block[4][85] ), .B(\block[6][85] ), .C(\block[5][85] ), 
        .D(\block[7][85] ), .S0(n754), .S1(n717), .Y(n1307) );
  MX2XL U1554 ( .A(n1300), .B(n1299), .S0(n5), .Y(n1302) );
  MX4X1 U1555 ( .A(\block[0][83] ), .B(\block[2][83] ), .C(\block[1][83] ), 
        .D(\block[3][83] ), .S0(n754), .S1(n716), .Y(n1300) );
  MX4X1 U1556 ( .A(\block[4][83] ), .B(\block[6][83] ), .C(\block[5][83] ), 
        .D(\block[7][83] ), .S0(n754), .S1(n716), .Y(n1299) );
  MX2XL U1557 ( .A(n1183), .B(n1182), .S0(n776), .Y(n1185) );
  MX4XL U1558 ( .A(\block[0][54] ), .B(\block[2][54] ), .C(\block[1][54] ), 
        .D(\block[3][54] ), .S0(n747), .S1(n711), .Y(n1183) );
  MX4XL U1559 ( .A(\block[4][54] ), .B(\block[6][54] ), .C(\block[5][54] ), 
        .D(\block[7][54] ), .S0(n747), .S1(n711), .Y(n1182) );
  MX2XL U1560 ( .A(n1312), .B(n1311), .S0(n774), .Y(n1314) );
  MX4XL U1561 ( .A(\block[0][86] ), .B(\block[2][86] ), .C(\block[1][86] ), 
        .D(\block[3][86] ), .S0(n754), .S1(n717), .Y(n1312) );
  MX4XL U1562 ( .A(\block[4][86] ), .B(\block[6][86] ), .C(\block[5][86] ), 
        .D(\block[7][86] ), .S0(n746), .S1(n717), .Y(n1311) );
  MX2XL U1563 ( .A(n1452), .B(n1451), .S0(n773), .Y(n1455) );
  MX2XL U1564 ( .A(n1050), .B(n1049), .S0(n777), .Y(n1052) );
  MX4X1 U1565 ( .A(\block[0][21] ), .B(\block[2][21] ), .C(\block[1][21] ), 
        .D(\block[3][21] ), .S0(n755), .S1(n729), .Y(n1050) );
  MX4XL U1566 ( .A(\block[4][21] ), .B(\block[6][21] ), .C(\block[5][21] ), 
        .D(\block[7][21] ), .S0(n756), .S1(n730), .Y(n1049) );
  MX2XL U1567 ( .A(n1054), .B(n1053), .S0(n777), .Y(n1056) );
  MX4XL U1568 ( .A(\block[0][22] ), .B(\block[2][22] ), .C(\block[1][22] ), 
        .D(\block[3][22] ), .S0(n756), .S1(n730), .Y(n1054) );
  MX4XL U1569 ( .A(\block[4][22] ), .B(\block[6][22] ), .C(\block[5][22] ), 
        .D(\block[7][22] ), .S0(n756), .S1(n730), .Y(n1053) );
  MX2XL U1570 ( .A(n1167), .B(n1166), .S0(n776), .Y(n1169) );
  MX4XL U1571 ( .A(\block[0][50] ), .B(\block[2][50] ), .C(\block[1][50] ), 
        .D(\block[3][50] ), .S0(n760), .S1(n711), .Y(n1167) );
  MX4XL U1572 ( .A(\block[4][50] ), .B(\block[6][50] ), .C(\block[5][50] ), 
        .D(\block[7][50] ), .S0(n746), .S1(n711), .Y(n1166) );
  MX2XL U1573 ( .A(n1175), .B(n1174), .S0(n776), .Y(n1177) );
  MX4XL U1574 ( .A(\block[0][52] ), .B(\block[2][52] ), .C(\block[1][52] ), 
        .D(\block[3][52] ), .S0(n758), .S1(n711), .Y(n1175) );
  MX4XL U1575 ( .A(\block[4][52] ), .B(\block[6][52] ), .C(\block[5][52] ), 
        .D(\block[7][52] ), .S0(n747), .S1(n711), .Y(n1174) );
  MX2XL U1576 ( .A(n1296), .B(n1295), .S0(n774), .Y(n1298) );
  MX4X1 U1577 ( .A(\block[0][82] ), .B(\block[2][82] ), .C(\block[1][82] ), 
        .D(\block[3][82] ), .S0(n754), .S1(n716), .Y(n1296) );
  MX4X1 U1578 ( .A(\block[4][82] ), .B(\block[6][82] ), .C(\block[5][82] ), 
        .D(\block[7][82] ), .S0(n754), .S1(n716), .Y(n1295) );
  MX2XL U1579 ( .A(n1304), .B(n1303), .S0(n774), .Y(n1306) );
  MX4X1 U1580 ( .A(\block[0][84] ), .B(\block[2][84] ), .C(\block[1][84] ), 
        .D(\block[3][84] ), .S0(n754), .S1(n716), .Y(n1304) );
  MX4X1 U1581 ( .A(\block[4][84] ), .B(\block[6][84] ), .C(\block[5][84] ), 
        .D(\block[7][84] ), .S0(n754), .S1(n716), .Y(n1303) );
  MX2XL U1582 ( .A(n1199), .B(n1198), .S0(n775), .Y(n1201) );
  MX4XL U1583 ( .A(\block[0][58] ), .B(\block[2][58] ), .C(\block[1][58] ), 
        .D(\block[3][58] ), .S0(n746), .S1(n712), .Y(n1199) );
  MX4XL U1584 ( .A(\block[4][58] ), .B(\block[6][58] ), .C(\block[5][58] ), 
        .D(\block[7][58] ), .S0(n746), .S1(n712), .Y(n1198) );
  MX2XL U1585 ( .A(n1159), .B(n1158), .S0(n776), .Y(n1161) );
  MX4X1 U1586 ( .A(\block[0][48] ), .B(\block[2][48] ), .C(\block[1][48] ), 
        .D(\block[3][48] ), .S0(n760), .S1(n734), .Y(n1159) );
  MX4X1 U1587 ( .A(\block[4][48] ), .B(\block[6][48] ), .C(\block[5][48] ), 
        .D(\block[7][48] ), .S0(n760), .S1(n734), .Y(n1158) );
  MX2XL U1588 ( .A(n1191), .B(n1190), .S0(n776), .Y(n1193) );
  MX4XL U1589 ( .A(\block[0][56] ), .B(\block[2][56] ), .C(\block[1][56] ), 
        .D(\block[3][56] ), .S0(n747), .S1(n712), .Y(n1191) );
  MX4XL U1590 ( .A(\block[4][56] ), .B(\block[6][56] ), .C(\block[5][56] ), 
        .D(\block[7][56] ), .S0(n746), .S1(n712), .Y(n1190) );
  MX2XL U1591 ( .A(n1195), .B(n1194), .S0(n775), .Y(n1197) );
  MX4XL U1592 ( .A(\block[0][57] ), .B(\block[2][57] ), .C(\block[1][57] ), 
        .D(\block[3][57] ), .S0(n746), .S1(n712), .Y(n1195) );
  MX4XL U1593 ( .A(\block[4][57] ), .B(\block[6][57] ), .C(\block[5][57] ), 
        .D(\block[7][57] ), .S0(n746), .S1(n712), .Y(n1194) );
  MX2XL U1594 ( .A(n1187), .B(n1186), .S0(n776), .Y(n1189) );
  MX4XL U1595 ( .A(\block[0][55] ), .B(\block[2][55] ), .C(\block[1][55] ), 
        .D(\block[3][55] ), .S0(n758), .S1(n711), .Y(n1187) );
  MX4XL U1596 ( .A(\block[4][55] ), .B(\block[6][55] ), .C(\block[5][55] ), 
        .D(\block[7][55] ), .S0(n747), .S1(n712), .Y(n1186) );
  MX2XL U1597 ( .A(n1163), .B(n1162), .S0(n776), .Y(n1165) );
  MX4XL U1598 ( .A(\block[4][49] ), .B(\block[6][49] ), .C(\block[5][49] ), 
        .D(\block[7][49] ), .S0(n760), .S1(n717), .Y(n1162) );
  MX2XL U1599 ( .A(n1328), .B(n1327), .S0(n5), .Y(n1330) );
  MX4XL U1600 ( .A(\block[0][90] ), .B(\block[2][90] ), .C(\block[1][90] ), 
        .D(\block[3][90] ), .S0(n750), .S1(n717), .Y(n1328) );
  MX4XL U1601 ( .A(\block[4][90] ), .B(\block[6][90] ), .C(\block[5][90] ), 
        .D(\block[7][90] ), .S0(n758), .S1(n717), .Y(n1327) );
  MX2XL U1602 ( .A(n1288), .B(n1287), .S0(n774), .Y(n1290) );
  MX4X1 U1603 ( .A(\block[0][80] ), .B(\block[2][80] ), .C(\block[1][80] ), 
        .D(\block[3][80] ), .S0(n754), .S1(n716), .Y(n1288) );
  MX4X1 U1604 ( .A(\block[4][80] ), .B(\block[6][80] ), .C(\block[5][80] ), 
        .D(\block[7][80] ), .S0(n754), .S1(n716), .Y(n1287) );
  MX2XL U1605 ( .A(n1320), .B(n1319), .S0(n5), .Y(n1322) );
  MX4XL U1606 ( .A(\block[0][88] ), .B(\block[2][88] ), .C(\block[1][88] ), 
        .D(\block[3][88] ), .S0(n746), .S1(n717), .Y(n1320) );
  MX4XL U1607 ( .A(\block[4][88] ), .B(\block[6][88] ), .C(\block[5][88] ), 
        .D(\block[7][88] ), .S0(n746), .S1(n717), .Y(n1319) );
  MX2XL U1608 ( .A(n1324), .B(n1323), .S0(n5), .Y(n1326) );
  MX4XL U1609 ( .A(\block[0][89] ), .B(\block[2][89] ), .C(\block[1][89] ), 
        .D(\block[3][89] ), .S0(n746), .S1(n735), .Y(n1324) );
  MX4XL U1610 ( .A(\block[4][89] ), .B(\block[6][89] ), .C(\block[5][89] ), 
        .D(\block[7][89] ), .S0(n746), .S1(n717), .Y(n1323) );
  MX2XL U1611 ( .A(n1316), .B(n1315), .S0(n774), .Y(n1318) );
  MX4XL U1612 ( .A(\block[0][87] ), .B(\block[2][87] ), .C(\block[1][87] ), 
        .D(\block[3][87] ), .S0(n746), .S1(n717), .Y(n1316) );
  MX4XL U1613 ( .A(\block[4][87] ), .B(\block[6][87] ), .C(\block[5][87] ), 
        .D(\block[7][87] ), .S0(n746), .S1(n717), .Y(n1315) );
  MX2XL U1614 ( .A(n1292), .B(n1291), .S0(n774), .Y(n1294) );
  MX4X1 U1615 ( .A(\block[0][81] ), .B(\block[2][81] ), .C(\block[1][81] ), 
        .D(\block[3][81] ), .S0(n754), .S1(n716), .Y(n1292) );
  MX4X1 U1616 ( .A(\block[4][81] ), .B(\block[6][81] ), .C(\block[5][81] ), 
        .D(\block[7][81] ), .S0(n754), .S1(n716), .Y(n1291) );
  MX2XL U1617 ( .A(n1046), .B(n1045), .S0(n777), .Y(n1048) );
  MX4XL U1618 ( .A(\block[0][20] ), .B(\block[2][20] ), .C(\block[1][20] ), 
        .D(\block[3][20] ), .S0(n755), .S1(n730), .Y(n1046) );
  MX4XL U1619 ( .A(\block[4][20] ), .B(\block[6][20] ), .C(\block[5][20] ), 
        .D(\block[7][20] ), .S0(n755), .S1(n730), .Y(n1045) );
  MX2XL U1620 ( .A(n1437), .B(n1436), .S0(n773), .Y(n1440) );
  MX4X1 U1621 ( .A(\block[0][112] ), .B(\block[2][112] ), .C(\block[1][112] ), 
        .D(\block[3][112] ), .S0(n749), .S1(n720), .Y(n1437) );
  MX2XL U1622 ( .A(n1442), .B(n1441), .S0(n773), .Y(n1445) );
  MX4X1 U1623 ( .A(\block[0][113] ), .B(\block[2][113] ), .C(\block[1][113] ), 
        .D(\block[3][113] ), .S0(n759), .S1(n720), .Y(n1442) );
  MX2XL U1624 ( .A(n1058), .B(n1057), .S0(n777), .Y(n1060) );
  MX4XL U1625 ( .A(\block[0][23] ), .B(\block[2][23] ), .C(\block[1][23] ), 
        .D(\block[3][23] ), .S0(n756), .S1(n730), .Y(n1058) );
  MX4XL U1626 ( .A(\block[4][23] ), .B(\block[6][23] ), .C(\block[5][23] ), 
        .D(\block[7][23] ), .S0(n756), .S1(n730), .Y(n1057) );
  MX2XL U1627 ( .A(n1062), .B(n1061), .S0(n777), .Y(n1064) );
  MX4XL U1628 ( .A(\block[0][24] ), .B(\block[2][24] ), .C(\block[1][24] ), 
        .D(\block[3][24] ), .S0(n756), .S1(n730), .Y(n1062) );
  MX4XL U1629 ( .A(\block[4][24] ), .B(\block[6][24] ), .C(\block[5][24] ), 
        .D(\block[7][24] ), .S0(n756), .S1(n730), .Y(n1061) );
  MX2XL U1630 ( .A(n1066), .B(n1065), .S0(n777), .Y(n1068) );
  MX4XL U1631 ( .A(\block[0][25] ), .B(\block[2][25] ), .C(\block[1][25] ), 
        .D(\block[3][25] ), .S0(n756), .S1(n730), .Y(n1066) );
  MX4XL U1632 ( .A(\block[4][25] ), .B(\block[6][25] ), .C(\block[5][25] ), 
        .D(\block[7][25] ), .S0(n756), .S1(n730), .Y(n1065) );
  MX2XL U1633 ( .A(n1070), .B(n1069), .S0(n777), .Y(n1072) );
  MX4XL U1634 ( .A(\block[0][26] ), .B(\block[2][26] ), .C(\block[1][26] ), 
        .D(\block[3][26] ), .S0(n756), .S1(n731), .Y(n1070) );
  MX4XL U1635 ( .A(\block[4][26] ), .B(\block[6][26] ), .C(\block[5][26] ), 
        .D(\block[7][26] ), .S0(n756), .S1(n731), .Y(n1069) );
  NAND3BXL U1636 ( .AN(n960), .B(proc_write), .C(n796), .Y(n955) );
  CLKINVX1 U1637 ( .A(proc_wdata[0]), .Y(n1359) );
  CLKINVX1 U1638 ( .A(proc_wdata[1]), .Y(n1364) );
  CLKINVX1 U1639 ( .A(proc_wdata[2]), .Y(n1369) );
  CLKINVX1 U1640 ( .A(proc_wdata[3]), .Y(n1374) );
  CLKINVX1 U1641 ( .A(proc_wdata[4]), .Y(n1379) );
  CLKINVX1 U1642 ( .A(proc_wdata[5]), .Y(n1384) );
  CLKINVX1 U1643 ( .A(proc_wdata[6]), .Y(n1389) );
  CLKINVX1 U1644 ( .A(proc_wdata[7]), .Y(n1394) );
  CLKINVX1 U1645 ( .A(proc_wdata[8]), .Y(n1399) );
  CLKINVX1 U1646 ( .A(proc_wdata[9]), .Y(n1404) );
  CLKINVX1 U1647 ( .A(proc_wdata[10]), .Y(n1409) );
  CLKINVX1 U1648 ( .A(proc_wdata[11]), .Y(n1414) );
  CLKINVX1 U1649 ( .A(proc_wdata[12]), .Y(n1419) );
  CLKINVX1 U1650 ( .A(proc_wdata[13]), .Y(n1424) );
  CLKINVX1 U1651 ( .A(proc_wdata[14]), .Y(n1429) );
  CLKINVX1 U1652 ( .A(proc_wdata[15]), .Y(n1434) );
  CLKINVX1 U1653 ( .A(proc_wdata[16]), .Y(n1439) );
  CLKINVX1 U1654 ( .A(proc_wdata[17]), .Y(n1444) );
  CLKINVX1 U1655 ( .A(proc_wdata[18]), .Y(n1449) );
  CLKINVX1 U1656 ( .A(proc_wdata[19]), .Y(n1454) );
  CLKINVX1 U1657 ( .A(proc_wdata[20]), .Y(n1459) );
  CLKINVX1 U1658 ( .A(proc_wdata[21]), .Y(n1464) );
  CLKINVX1 U1659 ( .A(proc_wdata[22]), .Y(n1469) );
  CLKINVX1 U1660 ( .A(proc_wdata[23]), .Y(n1474) );
  CLKINVX1 U1661 ( .A(proc_wdata[24]), .Y(n1479) );
  CLKINVX1 U1662 ( .A(proc_wdata[25]), .Y(n1484) );
  CLKINVX1 U1663 ( .A(proc_wdata[26]), .Y(n1489) );
  CLKINVX1 U1664 ( .A(proc_wdata[27]), .Y(n1494) );
  CLKINVX1 U1665 ( .A(proc_wdata[28]), .Y(n1499) );
  CLKINVX1 U1666 ( .A(proc_wdata[29]), .Y(n1502) );
  CLKINVX1 U1667 ( .A(proc_wdata[30]), .Y(n1507) );
  CLKINVX1 U1668 ( .A(proc_wdata[31]), .Y(n1513) );
  CLKINVX1 U1669 ( .A(proc_write), .Y(n1538) );
  NAND3BX4 U1670 ( .AN(n1549), .B(n1544), .C(n1548), .Y(n1709) );
  NAND2X2 U1671 ( .A(n1538), .B(n796), .Y(n966) );
  MX4X2 U1672 ( .A(blockvalid[0]), .B(blockvalid[2]), .C(blockvalid[1]), .D(
        blockvalid[3]), .S0(n103), .S1(n711), .Y(n798) );
  MX4X2 U1673 ( .A(blockvalid[4]), .B(blockvalid[6]), .C(blockvalid[5]), .D(
        blockvalid[7]), .S0(n444), .S1(n728), .Y(n797) );
  CLKINVX3 U1674 ( .A(n799), .Y(n803) );
  CLKINVX3 U1675 ( .A(n886), .Y(blocktag_next[3]) );
  CLKINVX3 U1676 ( .A(n890), .Y(blocktag_next[18]) );
  CLKINVX3 U1677 ( .A(n892), .Y(blocktag_next[2]) );
  CLKINVX3 U1678 ( .A(n897), .Y(blocktag_next[4]) );
  CLKINVX3 U1679 ( .A(n900), .Y(blocktag_next[6]) );
  CLKINVX3 U1680 ( .A(n901), .Y(blocktag_next[9]) );
  CLKINVX3 U1681 ( .A(n904), .Y(blocktag_next[8]) );
  CLKINVX3 U1682 ( .A(n907), .Y(blocktag_next[7]) );
  CLKINVX3 U1683 ( .A(n910), .Y(blocktag_next[11]) );
  CLKINVX3 U1684 ( .A(n913), .Y(blocktag_next[16]) );
  CLKINVX3 U1685 ( .A(n918), .Y(blocktag_next[13]) );
  CLKINVX3 U1686 ( .A(n923), .Y(blocktag_next[1]) );
  CLKINVX3 U1687 ( .A(n929), .Y(blocktag_next[22]) );
  CLKINVX3 U1688 ( .A(n932), .Y(blocktag_next[19]) );
  CLKINVX3 U1689 ( .A(n935), .Y(blocktag_next[20]) );
  CLKINVX3 U1690 ( .A(n938), .Y(blocktag_next[21]) );
  CLKINVX3 U1691 ( .A(n941), .Y(blocktag_next[0]) );
  CLKINVX3 U1692 ( .A(n944), .Y(blocktag_next[24]) );
  CLKINVX3 U1693 ( .A(n950), .Y(n954) );
  CLKMX2X4 U1694 ( .A(n970), .B(n969), .S0(n778), .Y(n972) );
  CLKINVX3 U1695 ( .A(n972), .Y(n1559) );
  CLKAND2X4 U1696 ( .A(n789), .B(n972), .Y(n1887) );
  CLKAND2X4 U1697 ( .A(n789), .B(n976), .Y(n1886) );
  CLKAND2X4 U1698 ( .A(n789), .B(n980), .Y(n1885) );
  CLKAND2X4 U1699 ( .A(n789), .B(n984), .Y(n1884) );
  CLKMX2X4 U1700 ( .A(n986), .B(n985), .S0(n778), .Y(n988) );
  CLKINVX3 U1701 ( .A(n988), .Y(n1579) );
  CLKAND2X4 U1702 ( .A(n789), .B(n988), .Y(n1883) );
  CLKAND2X4 U1703 ( .A(n789), .B(n992), .Y(n1882) );
  CLKAND2X4 U1704 ( .A(n791), .B(n1000), .Y(n1881) );
  CLKAND2X4 U1705 ( .A(n791), .B(n1004), .Y(n1880) );
  CLKAND2X4 U1706 ( .A(n791), .B(n1008), .Y(n1879) );
  CLKAND2X4 U1707 ( .A(n791), .B(n1012), .Y(n1878) );
  CLKAND2X4 U1708 ( .A(n791), .B(n1016), .Y(n1877) );
  CLKAND2X4 U1709 ( .A(n791), .B(n1020), .Y(n1876) );
  CLKAND2X4 U1710 ( .A(n791), .B(n1024), .Y(n1875) );
  CLKAND2X4 U1711 ( .A(n791), .B(n1028), .Y(n1874) );
  CLKAND2X4 U1712 ( .A(n791), .B(n1032), .Y(n1873) );
  CLKAND2X4 U1713 ( .A(n791), .B(n1036), .Y(n1872) );
  CLKAND2X4 U1714 ( .A(n791), .B(n1040), .Y(n1871) );
  CLKAND2X4 U1715 ( .A(n791), .B(n1044), .Y(n1870) );
  OAI221X2 U1716 ( .A0(n1459), .A1(n551), .B0(n1654), .B1(n545), .C0(n1047), 
        .Y(block_next[20]) );
  CLKAND2X4 U1717 ( .A(n791), .B(n1048), .Y(n1869) );
  CLKAND2X4 U1718 ( .A(n791), .B(n1052), .Y(n1868) );
  CLKAND2X4 U1719 ( .A(n791), .B(n1056), .Y(n1867) );
  CLKAND2X4 U1720 ( .A(n791), .B(n1060), .Y(n1866) );
  OAI221X2 U1721 ( .A0(n1479), .A1(n551), .B0(n1674), .B1(n546), .C0(n1063), 
        .Y(block_next[24]) );
  CLKAND2X4 U1722 ( .A(n791), .B(n1064), .Y(n1865) );
  OAI221X2 U1723 ( .A0(n1484), .A1(n551), .B0(n1679), .B1(n546), .C0(n1067), 
        .Y(block_next[25]) );
  CLKAND2X4 U1724 ( .A(n791), .B(n1068), .Y(n1864) );
  OAI221X2 U1725 ( .A0(n1489), .A1(n552), .B0(n1684), .B1(n546), .C0(n1071), 
        .Y(block_next[26]) );
  CLKAND2X4 U1726 ( .A(n791), .B(n1072), .Y(n1863) );
  MX4X2 U1727 ( .A(\block[0][27] ), .B(\block[2][27] ), .C(\block[1][27] ), 
        .D(\block[3][27] ), .S0(n756), .S1(n730), .Y(n1074) );
  CLKMX2X4 U1728 ( .A(n1074), .B(n1073), .S0(n777), .Y(n1076) );
  CLKINVX3 U1729 ( .A(n1076), .Y(n1689) );
  CLKMX2X4 U1730 ( .A(n1078), .B(n1077), .S0(n777), .Y(n1080) );
  CLKINVX3 U1731 ( .A(n1080), .Y(n1694) );
  CLKAND2X4 U1732 ( .A(n791), .B(n1080), .Y(n1862) );
  CLKMX2X4 U1733 ( .A(n1082), .B(n1081), .S0(n777), .Y(n1084) );
  CLKINVX3 U1734 ( .A(n1084), .Y(n1698) );
  CLKAND2X4 U1735 ( .A(n791), .B(n1084), .Y(n1861) );
  CLKMX2X4 U1736 ( .A(n1086), .B(n1085), .S0(n777), .Y(n1088) );
  CLKINVX3 U1737 ( .A(n1088), .Y(n1703) );
  CLKAND2X4 U1738 ( .A(n791), .B(n1088), .Y(n1860) );
  MX4X2 U1739 ( .A(\block[0][31] ), .B(\block[2][31] ), .C(\block[1][31] ), 
        .D(\block[3][31] ), .S0(n757), .S1(n731), .Y(n1090) );
  CLKMX2X4 U1740 ( .A(n1090), .B(n1089), .S0(n777), .Y(n1093) );
  CLKINVX3 U1741 ( .A(n1093), .Y(n1710) );
  CLKAND2X4 U1742 ( .A(n791), .B(n1093), .Y(n1859) );
  CLKAND2X4 U1743 ( .A(n791), .B(n1097), .Y(n1858) );
  CLKAND2X4 U1744 ( .A(n791), .B(n1101), .Y(n1857) );
  CLKAND2X4 U1745 ( .A(n791), .B(n1105), .Y(n1856) );
  CLKAND2X4 U1746 ( .A(n791), .B(n1109), .Y(n1855) );
  CLKAND2X4 U1747 ( .A(n791), .B(n1113), .Y(n1854) );
  CLKAND2X4 U1748 ( .A(n790), .B(n1117), .Y(n1853) );
  CLKAND2X4 U1749 ( .A(n791), .B(n1121), .Y(n1852) );
  CLKAND2X4 U1750 ( .A(n791), .B(n1125), .Y(n1851) );
  CLKAND2X4 U1751 ( .A(n791), .B(n1129), .Y(n1850) );
  CLKAND2X4 U1752 ( .A(n791), .B(n1133), .Y(n1849) );
  CLKAND2X4 U1753 ( .A(n791), .B(n1137), .Y(n1848) );
  CLKAND2X4 U1754 ( .A(n791), .B(n1141), .Y(n1847) );
  CLKAND2X4 U1755 ( .A(n791), .B(n1145), .Y(n1846) );
  CLKAND2X4 U1756 ( .A(n791), .B(n1149), .Y(n1845) );
  CLKAND2X4 U1757 ( .A(n790), .B(n1157), .Y(n1844) );
  CLKAND2X4 U1758 ( .A(n790), .B(n1161), .Y(n1843) );
  CLKAND2X4 U1759 ( .A(n790), .B(n1165), .Y(n1842) );
  CLKAND2X4 U1760 ( .A(n790), .B(n1169), .Y(n1841) );
  CLKAND2X4 U1761 ( .A(n790), .B(n1173), .Y(n1840) );
  CLKAND2X4 U1762 ( .A(n790), .B(n1177), .Y(n1839) );
  CLKAND2X4 U1763 ( .A(n790), .B(n1181), .Y(n1838) );
  CLKAND2X4 U1764 ( .A(n790), .B(n1185), .Y(n1837) );
  CLKAND2X4 U1765 ( .A(n790), .B(n1189), .Y(n1836) );
  CLKAND2X4 U1766 ( .A(n790), .B(n1193), .Y(n1835) );
  CLKAND2X4 U1767 ( .A(n790), .B(n1197), .Y(n1834) );
  CLKAND2X4 U1768 ( .A(n790), .B(n1201), .Y(n1833) );
  MX4X2 U1769 ( .A(\block[0][59] ), .B(\block[2][59] ), .C(\block[1][59] ), 
        .D(\block[3][59] ), .S0(n746), .S1(n712), .Y(n1203) );
  MX4X2 U1770 ( .A(\block[4][59] ), .B(\block[6][59] ), .C(\block[5][59] ), 
        .D(\block[7][59] ), .S0(n746), .S1(n712), .Y(n1202) );
  CLKMX2X4 U1771 ( .A(n1203), .B(n1202), .S0(n775), .Y(n1205) );
  CLKINVX3 U1772 ( .A(n1205), .Y(n1685) );
  MX4X2 U1773 ( .A(\block[0][60] ), .B(\block[2][60] ), .C(\block[1][60] ), 
        .D(\block[3][60] ), .S0(n746), .S1(n712), .Y(n1207) );
  MX4X2 U1774 ( .A(\block[4][60] ), .B(\block[6][60] ), .C(\block[5][60] ), 
        .D(\block[7][60] ), .S0(n746), .S1(n712), .Y(n1206) );
  CLKMX2X4 U1775 ( .A(n1207), .B(n1206), .S0(n775), .Y(n1209) );
  CLKINVX3 U1776 ( .A(n1209), .Y(n1690) );
  CLKAND2X4 U1777 ( .A(n790), .B(n1209), .Y(n1832) );
  MX4X2 U1778 ( .A(\block[0][61] ), .B(\block[2][61] ), .C(\block[1][61] ), 
        .D(\block[3][61] ), .S0(n746), .S1(n712), .Y(n1211) );
  CLKMX2X4 U1779 ( .A(n1211), .B(n1210), .S0(n775), .Y(n1213) );
  CLKINVX3 U1780 ( .A(n1213), .Y(n1695) );
  CLKAND2X4 U1781 ( .A(n790), .B(n1213), .Y(n1831) );
  MX4X2 U1782 ( .A(\block[0][62] ), .B(\block[2][62] ), .C(\block[1][62] ), 
        .D(\block[3][62] ), .S0(n746), .S1(n713), .Y(n1215) );
  MX4X2 U1783 ( .A(\block[4][62] ), .B(\block[6][62] ), .C(\block[5][62] ), 
        .D(\block[7][62] ), .S0(n747), .S1(n713), .Y(n1214) );
  CLKMX2X4 U1784 ( .A(n1215), .B(n1214), .S0(n775), .Y(n1217) );
  CLKINVX3 U1785 ( .A(n1217), .Y(n1699) );
  CLKAND2X4 U1786 ( .A(n790), .B(n1217), .Y(n1830) );
  MX4X2 U1787 ( .A(\block[0][63] ), .B(\block[2][63] ), .C(\block[1][63] ), 
        .D(\block[3][63] ), .S0(n747), .S1(n713), .Y(n1219) );
  MX4X2 U1788 ( .A(\block[4][63] ), .B(\block[6][63] ), .C(\block[5][63] ), 
        .D(\block[7][63] ), .S0(n747), .S1(n713), .Y(n1218) );
  CLKMX2X4 U1789 ( .A(n1219), .B(n1218), .S0(n775), .Y(n1221) );
  CLKINVX3 U1790 ( .A(n1221), .Y(n1704) );
  CLKAND2X4 U1791 ( .A(n790), .B(n1221), .Y(n1829) );
  CLKINVX3 U1792 ( .A(n1224), .Y(n1350) );
  CLKAND2X4 U1793 ( .A(n790), .B(n1226), .Y(n1828) );
  CLKAND2X4 U1794 ( .A(n790), .B(n1230), .Y(n1827) );
  CLKAND2X4 U1795 ( .A(n790), .B(n1234), .Y(n1826) );
  OAI221X2 U1796 ( .A0(n1566), .A1(n549), .B0(n1374), .B1(n557), .C0(n1237), 
        .Y(block_next[67]) );
  CLKAND2X4 U1797 ( .A(n790), .B(n1238), .Y(n1825) );
  OAI221X2 U1798 ( .A0(n1571), .A1(n549), .B0(n1379), .B1(n557), .C0(n1241), 
        .Y(block_next[68]) );
  CLKAND2X4 U1799 ( .A(n790), .B(n1242), .Y(n1824) );
  OAI221X2 U1800 ( .A0(n1576), .A1(n549), .B0(n1384), .B1(n557), .C0(n1245), 
        .Y(block_next[69]) );
  CLKAND2X4 U1801 ( .A(n790), .B(n1246), .Y(n1823) );
  OAI221X2 U1802 ( .A0(n1581), .A1(n549), .B0(n1389), .B1(n557), .C0(n1249), 
        .Y(block_next[70]) );
  CLKAND2X4 U1803 ( .A(n790), .B(n1250), .Y(n1822) );
  OAI221X2 U1804 ( .A0(n1586), .A1(n549), .B0(n1394), .B1(n557), .C0(n1253), 
        .Y(block_next[71]) );
  CLKAND2X4 U1805 ( .A(n790), .B(n1254), .Y(n1821) );
  OAI221X2 U1806 ( .A0(n1591), .A1(n549), .B0(n1399), .B1(n556), .C0(n1257), 
        .Y(block_next[72]) );
  CLKAND2X4 U1807 ( .A(n790), .B(n1258), .Y(n1820) );
  OAI221X2 U1808 ( .A0(n1596), .A1(n549), .B0(n1404), .B1(n556), .C0(n1261), 
        .Y(block_next[73]) );
  CLKAND2X4 U1809 ( .A(n790), .B(n1262), .Y(n1819) );
  OAI221X2 U1810 ( .A0(n1601), .A1(n549), .B0(n1409), .B1(n556), .C0(n1265), 
        .Y(block_next[74]) );
  CLKAND2X4 U1811 ( .A(n790), .B(n1266), .Y(n1818) );
  OAI221X2 U1812 ( .A0(n1606), .A1(n549), .B0(n1414), .B1(n556), .C0(n1269), 
        .Y(block_next[75]) );
  CLKAND2X4 U1813 ( .A(n790), .B(n1270), .Y(n1817) );
  OAI221X2 U1814 ( .A0(n1611), .A1(n549), .B0(n1419), .B1(n556), .C0(n1273), 
        .Y(block_next[76]) );
  CLKAND2X4 U1815 ( .A(n790), .B(n1274), .Y(n1816) );
  CLKAND2X4 U1816 ( .A(n790), .B(n1278), .Y(n1815) );
  CLKAND2X4 U1817 ( .A(n790), .B(n1282), .Y(n1814) );
  CLKAND2X4 U1818 ( .A(n790), .B(n1286), .Y(n1813) );
  CLKAND2X4 U1819 ( .A(n789), .B(n1306), .Y(n1811) );
  CLKAND2X4 U1820 ( .A(n789), .B(n1310), .Y(n1810) );
  CLKAND2X4 U1821 ( .A(n789), .B(n1314), .Y(n1809) );
  CLKAND2X4 U1822 ( .A(n789), .B(n1318), .Y(n1808) );
  CLKAND2X4 U1823 ( .A(n789), .B(n1322), .Y(n1807) );
  CLKAND2X4 U1824 ( .A(n789), .B(n1326), .Y(n1806) );
  CLKAND2X4 U1825 ( .A(n789), .B(n1330), .Y(n1805) );
  MX4X2 U1826 ( .A(\block[0][91] ), .B(\block[2][91] ), .C(\block[1][91] ), 
        .D(\block[3][91] ), .S0(n746), .S1(n717), .Y(n1332) );
  MX4X2 U1827 ( .A(\block[4][91] ), .B(\block[6][91] ), .C(\block[5][91] ), 
        .D(\block[7][91] ), .S0(n755), .S1(n734), .Y(n1331) );
  OAI221X2 U1828 ( .A0(n1686), .A1(n550), .B0(n1494), .B1(n1356), .C0(n1333), 
        .Y(block_next[91]) );
  MX4X2 U1829 ( .A(\block[0][92] ), .B(\block[2][92] ), .C(\block[1][92] ), 
        .D(\block[3][92] ), .S0(n746), .S1(n734), .Y(n1336) );
  MX4X2 U1830 ( .A(\block[4][92] ), .B(\block[6][92] ), .C(\block[5][92] ), 
        .D(\block[7][92] ), .S0(n748), .S1(n734), .Y(n1335) );
  CLKMX2X4 U1831 ( .A(n1336), .B(n1335), .S0(n776), .Y(n1338) );
  CLKINVX3 U1832 ( .A(n1338), .Y(n1691) );
  CLKMX2X4 U1833 ( .A(n1340), .B(n1339), .S0(n774), .Y(n1342) );
  CLKINVX3 U1834 ( .A(n1342), .Y(n1696) );
  OAI221X2 U1835 ( .A0(n1696), .A1(n550), .B0(n1502), .B1(n557), .C0(n1341), 
        .Y(block_next[93]) );
  OAI221X2 U1836 ( .A0(n1700), .A1(n550), .B0(n1507), .B1(n557), .C0(n1345), 
        .Y(block_next[94]) );
  CLKAND2X4 U1837 ( .A(n789), .B(n1346), .Y(n1804) );
  CLKMX2X4 U1838 ( .A(n1348), .B(n1347), .S0(n773), .Y(n1351) );
  CLKINVX3 U1839 ( .A(n1351), .Y(n1706) );
  OAI221X2 U1840 ( .A0(n1706), .A1(n550), .B0(n1513), .B1(n556), .C0(n1349), 
        .Y(block_next[95]) );
  CLKINVX3 U1841 ( .A(n1357), .Y(n1515) );
  OAI221X2 U1842 ( .A0(n1553), .A1(n576), .B0(n575), .B1(n1359), .C0(n1358), 
        .Y(block_next[96]) );
  CLKAND2X4 U1843 ( .A(n789), .B(n1360), .Y(n1803) );
  OAI221X2 U1844 ( .A0(n1558), .A1(n576), .B0(n575), .B1(n1364), .C0(n1363), 
        .Y(block_next[97]) );
  CLKAND2X4 U1845 ( .A(n789), .B(n1365), .Y(n1802) );
  OAI221X2 U1846 ( .A0(n1563), .A1(n576), .B0(n575), .B1(n1369), .C0(n1368), 
        .Y(block_next[98]) );
  CLKAND2X4 U1847 ( .A(n789), .B(n1370), .Y(n1801) );
  OAI221X2 U1848 ( .A0(n1568), .A1(n576), .B0(n575), .B1(n1374), .C0(n1373), 
        .Y(block_next[99]) );
  CLKAND2X4 U1849 ( .A(n789), .B(n1375), .Y(n1800) );
  OAI221X2 U1850 ( .A0(n1573), .A1(n576), .B0(n575), .B1(n1379), .C0(n1378), 
        .Y(block_next[100]) );
  CLKAND2X4 U1851 ( .A(n789), .B(n1380), .Y(n1799) );
  OAI221X2 U1852 ( .A0(n1578), .A1(n576), .B0(n575), .B1(n1384), .C0(n1383), 
        .Y(block_next[101]) );
  CLKAND2X4 U1853 ( .A(n789), .B(n1385), .Y(n1798) );
  OAI221X2 U1854 ( .A0(n1583), .A1(n576), .B0(n575), .B1(n1389), .C0(n1388), 
        .Y(block_next[102]) );
  CLKAND2X4 U1855 ( .A(n789), .B(n1390), .Y(n1797) );
  OAI221X2 U1856 ( .A0(n1588), .A1(n576), .B0(n575), .B1(n1394), .C0(n1393), 
        .Y(block_next[103]) );
  CLKAND2X4 U1857 ( .A(n789), .B(n1395), .Y(n1796) );
  OAI221X2 U1858 ( .A0(n1593), .A1(n576), .B0(n574), .B1(n1399), .C0(n1398), 
        .Y(block_next[104]) );
  CLKAND2X4 U1859 ( .A(n789), .B(n1400), .Y(n1795) );
  OAI221X2 U1860 ( .A0(n1598), .A1(n576), .B0(n574), .B1(n1404), .C0(n1403), 
        .Y(block_next[105]) );
  CLKAND2X4 U1861 ( .A(n789), .B(n1405), .Y(n1794) );
  OAI221X2 U1862 ( .A0(n1603), .A1(n576), .B0(n574), .B1(n1409), .C0(n1408), 
        .Y(block_next[106]) );
  CLKAND2X4 U1863 ( .A(n789), .B(n1410), .Y(n1793) );
  OAI221X2 U1864 ( .A0(n1608), .A1(n576), .B0(n574), .B1(n1414), .C0(n1413), 
        .Y(block_next[107]) );
  CLKAND2X4 U1865 ( .A(n789), .B(n1415), .Y(n1792) );
  OAI221X2 U1866 ( .A0(n1613), .A1(n576), .B0(n574), .B1(n1419), .C0(n1418), 
        .Y(block_next[108]) );
  CLKAND2X4 U1867 ( .A(n789), .B(n1420), .Y(n1791) );
  OAI221X2 U1868 ( .A0(n1618), .A1(n577), .B0(n574), .B1(n1424), .C0(n1423), 
        .Y(block_next[109]) );
  CLKAND2X4 U1869 ( .A(n789), .B(n1425), .Y(n1790) );
  OAI221X2 U1870 ( .A0(n1623), .A1(n577), .B0(n574), .B1(n1429), .C0(n1428), 
        .Y(block_next[110]) );
  CLKAND2X4 U1871 ( .A(n789), .B(n1430), .Y(n1789) );
  OAI221X2 U1872 ( .A0(n1628), .A1(n577), .B0(n574), .B1(n1434), .C0(n1433), 
        .Y(block_next[111]) );
  CLKAND2X4 U1873 ( .A(n789), .B(n1435), .Y(n1788) );
  OAI221X2 U1874 ( .A0(n1633), .A1(n577), .B0(n574), .B1(n1439), .C0(n1438), 
        .Y(block_next[112]) );
  CLKAND2X4 U1875 ( .A(n789), .B(n1440), .Y(n1787) );
  OAI221X2 U1876 ( .A0(n1638), .A1(n577), .B0(n574), .B1(n1444), .C0(n1443), 
        .Y(block_next[113]) );
  CLKAND2X4 U1877 ( .A(n789), .B(n1445), .Y(n1786) );
  OAI221X2 U1878 ( .A0(n1643), .A1(n577), .B0(n574), .B1(n1449), .C0(n1448), 
        .Y(block_next[114]) );
  CLKAND2X4 U1879 ( .A(n789), .B(n1450), .Y(n1785) );
  OAI221X2 U1880 ( .A0(n1648), .A1(n577), .B0(n574), .B1(n1454), .C0(n1453), 
        .Y(block_next[115]) );
  CLKAND2X4 U1881 ( .A(n789), .B(n1455), .Y(n1784) );
  OAI221X2 U1882 ( .A0(n1653), .A1(n577), .B0(n573), .B1(n1459), .C0(n1458), 
        .Y(block_next[116]) );
  CLKAND2X4 U1883 ( .A(n789), .B(n1460), .Y(n1783) );
  OAI221X2 U1884 ( .A0(n1658), .A1(n577), .B0(n573), .B1(n1464), .C0(n1463), 
        .Y(block_next[117]) );
  CLKAND2X4 U1885 ( .A(n789), .B(n1465), .Y(n1782) );
  OAI221X2 U1886 ( .A0(n1663), .A1(n577), .B0(n573), .B1(n1469), .C0(n1468), 
        .Y(block_next[118]) );
  CLKAND2X4 U1887 ( .A(n789), .B(n1470), .Y(n1781) );
  OAI221X2 U1888 ( .A0(n1668), .A1(n577), .B0(n573), .B1(n1474), .C0(n1473), 
        .Y(block_next[119]) );
  CLKAND2X4 U1889 ( .A(n789), .B(n1475), .Y(n1780) );
  OAI221X2 U1890 ( .A0(n1673), .A1(n577), .B0(n573), .B1(n1479), .C0(n1478), 
        .Y(block_next[120]) );
  CLKAND2X4 U1891 ( .A(n789), .B(n1480), .Y(n1779) );
  OAI221X2 U1892 ( .A0(n1678), .A1(n577), .B0(n573), .B1(n1484), .C0(n1483), 
        .Y(block_next[121]) );
  CLKAND2X4 U1893 ( .A(n789), .B(n1485), .Y(n1778) );
  OAI221X2 U1894 ( .A0(n1683), .A1(n578), .B0(n573), .B1(n1489), .C0(n1488), 
        .Y(block_next[122]) );
  CLKAND2X4 U1895 ( .A(mem_write), .B(n1490), .Y(n1777) );
  OAI221X2 U1896 ( .A0(n1688), .A1(n578), .B0(n573), .B1(n1494), .C0(n1493), 
        .Y(block_next[123]) );
  OAI221X2 U1897 ( .A0(n1693), .A1(n578), .B0(n573), .B1(n1499), .C0(n1498), 
        .Y(block_next[124]) );
  OAI221X2 U1898 ( .A0(n527), .A1(n578), .B0(n573), .B1(n1502), .C0(n1501), 
        .Y(block_next[125]) );
  CLKAND2X4 U1899 ( .A(mem_write), .B(n1503), .Y(n1776) );
  OAI221X2 U1900 ( .A0(n1702), .A1(n578), .B0(n573), .B1(n1507), .C0(n1506), 
        .Y(block_next[126]) );
  OAI221X2 U1901 ( .A0(n1708), .A1(n578), .B0(n573), .B1(n1513), .C0(n1512), 
        .Y(block_next[127]) );
  AO22X4 U1902 ( .A0(proc_addr[6]), .A1(mem_read), .B0(mem_write), .B1(n112), 
        .Y(n1772) );
  AO22X4 U1903 ( .A0(proc_addr[7]), .A1(mem_read), .B0(mem_write), .B1(n408), 
        .Y(n1771) );
  AO22X4 U1904 ( .A0(proc_addr[8]), .A1(mem_read), .B0(mem_write), .B1(n418), 
        .Y(n1770) );
  AO22X4 U1905 ( .A0(proc_addr[9]), .A1(mem_read), .B0(mem_write), .B1(n24), 
        .Y(n1769) );
  AO22X4 U1906 ( .A0(proc_addr[11]), .A1(mem_read), .B0(mem_write), .B1(n1525), 
        .Y(n1767) );
  AO22X4 U1907 ( .A0(proc_addr[12]), .A1(mem_read), .B0(mem_write), .B1(n105), 
        .Y(n1766) );
  AO22X4 U1908 ( .A0(proc_addr[13]), .A1(mem_read), .B0(mem_write), .B1(n430), 
        .Y(n1765) );
  AO22X4 U1909 ( .A0(proc_addr[14]), .A1(mem_read), .B0(mem_write), .B1(n522), 
        .Y(n1764) );
  AO22X4 U1910 ( .A0(proc_addr[16]), .A1(mem_read), .B0(mem_write), .B1(n448), 
        .Y(n1762) );
  AO22X4 U1911 ( .A0(proc_addr[17]), .A1(mem_read), .B0(mem_write), .B1(n440), 
        .Y(n1761) );
  AO22X4 U1912 ( .A0(proc_addr[18]), .A1(mem_read), .B0(mem_write), .B1(n113), 
        .Y(n1760) );
  AO22X4 U1913 ( .A0(proc_addr[19]), .A1(mem_read), .B0(mem_write), .B1(n429), 
        .Y(n1759) );
  AO22X4 U1914 ( .A0(proc_addr[20]), .A1(mem_read), .B0(mem_write), .B1(n458), 
        .Y(n1758) );
  AO22X4 U1915 ( .A0(proc_addr[21]), .A1(mem_read), .B0(mem_write), .B1(n443), 
        .Y(n1757) );
  AO22X4 U1916 ( .A0(proc_addr[22]), .A1(mem_read), .B0(mem_write), .B1(n405), 
        .Y(n1756) );
  AO22X4 U1917 ( .A0(proc_addr[23]), .A1(mem_read), .B0(mem_write), .B1(n437), 
        .Y(n1755) );
  AO22X4 U1918 ( .A0(proc_addr[24]), .A1(mem_read), .B0(mem_write), .B1(n1533), 
        .Y(n1754) );
  AO22X4 U1919 ( .A0(proc_addr[25]), .A1(mem_read), .B0(mem_write), .B1(n1534), 
        .Y(n1753) );
  AO22X4 U1920 ( .A0(proc_addr[29]), .A1(mem_read), .B0(mem_write), .B1(n3), 
        .Y(n1750) );
  OAI221X2 U1921 ( .A0(n1554), .A1(n505), .B0(n1553), .B1(n582), .C0(n1552), 
        .Y(proc_rdata[0]) );
  OAI221X2 U1922 ( .A0(n1559), .A1(n505), .B0(n1558), .B1(n582), .C0(n1557), 
        .Y(proc_rdata[1]) );
  OAI221X2 U1923 ( .A0(n1569), .A1(n505), .B0(n1568), .B1(n582), .C0(n1567), 
        .Y(proc_rdata[3]) );
  OAI221X2 U1924 ( .A0(n1574), .A1(n505), .B0(n1573), .B1(n582), .C0(n1572), 
        .Y(proc_rdata[4]) );
  OAI221X2 U1925 ( .A0(n1579), .A1(n505), .B0(n1578), .B1(n582), .C0(n1577), 
        .Y(proc_rdata[5]) );
  OAI221X2 U1926 ( .A0(n1594), .A1(n505), .B0(n1593), .B1(n582), .C0(n1592), 
        .Y(proc_rdata[8]) );
  OAI221X2 U1927 ( .A0(n1624), .A1(n505), .B0(n1623), .B1(n583), .C0(n1622), 
        .Y(proc_rdata[14]) );
  OA22X4 U1928 ( .A0(n1686), .A1(n91), .B0(n97), .B1(n1685), .Y(n1687) );
  OAI221X2 U1929 ( .A0(n96), .A1(n1689), .B0(n1688), .B1(n520), .C0(n1687), 
        .Y(proc_rdata[27]) );
  OA22X4 U1930 ( .A0(n1691), .A1(n1705), .B0(n541), .B1(n1690), .Y(n1692) );
  OAI221X2 U1931 ( .A0(n1694), .A1(n96), .B0(n1693), .B1(n520), .C0(n1692), 
        .Y(proc_rdata[28]) );
  OA22X4 U1932 ( .A0(n1705), .A1(n1696), .B0(n541), .B1(n1695), .Y(n1697) );
  OAI221X2 U1933 ( .A0(n96), .A1(n1698), .B0(n527), .B1(n520), .C0(n1697), .Y(
        proc_rdata[29]) );
  OA22X4 U1934 ( .A0(n1700), .A1(n91), .B0(n1699), .B1(n541), .Y(n1701) );
  OAI221X2 U1935 ( .A0(n1703), .A1(n96), .B0(n1702), .B1(n520), .C0(n1701), 
        .Y(proc_rdata[30]) );
  OA22X4 U1936 ( .A0(n91), .A1(n1706), .B0(n97), .B1(n1704), .Y(n1707) );
  OAI221X2 U1937 ( .A0(n1710), .A1(n96), .B0(n1708), .B1(n520), .C0(n1707), 
        .Y(proc_rdata[31]) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, ICACHE_ren, ICACHE_stall,
         DCACHE_ren, DCACHE_stall, n2, n3, n4, n6, n8, n10, n12, n14, n16, n18,
         n20, n22, n24, n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46,
         n48, n50, n52, n54, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74,
         n76, n78, n80, n82, n84, n86, n88, n90, n92, n94, n96, n98, n100,
         n102, n104, n106, n108, n110, n112, n114, n116, n118, n120, n122,
         n124, n126, n128, n130, n132, n134, n136, n138, n140, n142, n144,
         n146, n148, n150, n152, n154, n156, n158, n160, n162, n164, n166,
         n168, n170, n172, n174, n176, n178, n180, n182, n184, n186, n188,
         n190, n192, n194, n196, n198, n200, n202, n204, n206, n208, n210,
         n212, n214, n216, n218, n220, n222, n224, n226, n228, n230, n232,
         n234, n236, n238, n240, n242, n244, n246, n248, n250, n252, n254,
         n256, n258, n260, n262, n264, n266, n268, n270, n277, n278;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n277), .ICACHE_ren(ICACHE_ren), 
        .ICACHE_addr(ICACHE_addr), .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(
        ICACHE_rdata), .DCACHE_ren(DCACHE_ren), .DCACHE_wen(DCACHE_wen), 
        .DCACHE_addr({DCACHE_addr[29:5], n415, n416, n417, DCACHE_addr[1:0]}), 
        .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(DCACHE_stall), 
        .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n278), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:5], n415, n416, 
        n417, DCACHE_addr[1:0]}), .proc_wdata(DCACHE_wdata), .proc_stall(
        DCACHE_stall), .proc_rdata(DCACHE_rdata), .mem_read(n279), .mem_write(
        n280), .mem_addr({mem_addr_D[31:29], n281, mem_addr_D[27:25], n282, 
        n283, mem_addr_D[22:21], n284, n285, mem_addr_D[18:13], n286, 
        mem_addr_D[11:7], n287, mem_addr_D[5:4]}), .mem_rdata(mem_rdata_D), 
        .mem_wdata({n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
        n298, n299, n300, n301, n302, n303, n304, n305, n306, mem_wdata_D[108], 
        n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
        n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
        n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
        n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
        n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
        n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
        n379, n380, n381, mem_wdata_D[32], n382, n383, n384, n385, n386, n387, 
        n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
        n400, n401, n402, n403, n404, n405, n406, mem_wdata_D[6:1], n407}), 
        .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n278), .proc_read(ICACHE_ren), 
        .proc_write(1'b0), .proc_addr(ICACHE_addr), .proc_wdata({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .proc_stall(ICACHE_stall), 
        .proc_rdata(ICACHE_rdata), .mem_read(n408), .mem_write(n409), 
        .mem_addr({mem_addr_I[31:5], n410}), .mem_rdata(mem_rdata_I), 
        .mem_wdata({n411, mem_wdata_I[126:84], n412, n413, n414, 
        mem_wdata_I[80:0]}), .mem_ready(mem_ready_I) );
  INVX1 U2 ( .A(n381), .Y(n184) );
  INVX1 U3 ( .A(n380), .Y(n190) );
  INVX1 U4 ( .A(n379), .Y(n196) );
  INVX1 U5 ( .A(n378), .Y(n202) );
  INVX1 U6 ( .A(n376), .Y(n210) );
  INVX1 U7 ( .A(n375), .Y(n218) );
  INVX1 U8 ( .A(n374), .Y(n226) );
  INVX1 U9 ( .A(n373), .Y(n234) );
  INVX1 U10 ( .A(n372), .Y(n242) );
  INVX1 U11 ( .A(n371), .Y(n250) );
  INVX1 U12 ( .A(n370), .Y(n258) );
  INVX1 U13 ( .A(n369), .Y(n266) );
  INVX1 U14 ( .A(n343), .Y(n186) );
  INVX1 U15 ( .A(n342), .Y(n192) );
  INVX1 U16 ( .A(n341), .Y(n198) );
  INVX1 U17 ( .A(n340), .Y(n204) );
  INVX1 U18 ( .A(n339), .Y(n212) );
  INVX1 U19 ( .A(n338), .Y(n220) );
  INVX1 U20 ( .A(n337), .Y(n228) );
  INVX1 U21 ( .A(n336), .Y(n236) );
  INVX1 U22 ( .A(n335), .Y(n244) );
  INVX1 U23 ( .A(n334), .Y(n252) );
  INVX1 U24 ( .A(n333), .Y(n260) );
  INVX1 U25 ( .A(n332), .Y(n268) );
  INVX1 U26 ( .A(n294), .Y(n216) );
  INVX1 U27 ( .A(n293), .Y(n224) );
  INVX1 U28 ( .A(n292), .Y(n232) );
  INVX1 U29 ( .A(n291), .Y(n240) );
  INVX1 U30 ( .A(n290), .Y(n248) );
  INVX1 U31 ( .A(n289), .Y(n256) );
  INVX1 U32 ( .A(n288), .Y(n264) );
  INVX3 U33 ( .A(n282), .Y(n174) );
  INVX3 U34 ( .A(n281), .Y(n176) );
  INVXL U35 ( .A(n416), .Y(n2) );
  CLKINVX1 U36 ( .A(n2), .Y(n3) );
  INVXL U37 ( .A(n415), .Y(n4) );
  INVX12 U38 ( .A(n4), .Y(DCACHE_addr[4]) );
  INVXL U39 ( .A(n417), .Y(n6) );
  INVX12 U40 ( .A(n6), .Y(DCACHE_addr[2]) );
  CLKINVX6 U41 ( .A(n286), .Y(n8) );
  INVX20 U42 ( .A(n8), .Y(mem_addr_D[12]) );
  CLKINVX6 U43 ( .A(n285), .Y(n10) );
  INVX20 U44 ( .A(n10), .Y(mem_addr_D[19]) );
  CLKINVX6 U45 ( .A(n284), .Y(n12) );
  INVX20 U46 ( .A(n12), .Y(mem_addr_D[20]) );
  CLKINVX6 U47 ( .A(n283), .Y(n14) );
  INVX20 U48 ( .A(n14), .Y(mem_addr_D[23]) );
  INVX4 U49 ( .A(n377), .Y(n16) );
  CLKINVX20 U50 ( .A(n16), .Y(mem_wdata_D[37]) );
  INVX4 U51 ( .A(n368), .Y(n18) );
  CLKINVX20 U52 ( .A(n18), .Y(mem_wdata_D[46]) );
  INVX4 U53 ( .A(n367), .Y(n20) );
  CLKINVX20 U54 ( .A(n20), .Y(mem_wdata_D[47]) );
  INVX4 U55 ( .A(n366), .Y(n22) );
  CLKINVX20 U56 ( .A(n22), .Y(mem_wdata_D[48]) );
  INVX4 U57 ( .A(n365), .Y(n24) );
  CLKINVX20 U58 ( .A(n24), .Y(mem_wdata_D[49]) );
  INVX4 U59 ( .A(n406), .Y(n26) );
  CLKINVX20 U60 ( .A(n26), .Y(mem_wdata_D[7]) );
  INVX4 U61 ( .A(n364), .Y(n28) );
  CLKINVX20 U62 ( .A(n28), .Y(mem_wdata_D[50]) );
  INVX4 U63 ( .A(n405), .Y(n30) );
  CLKINVX20 U64 ( .A(n30), .Y(mem_wdata_D[8]) );
  INVX4 U65 ( .A(n363), .Y(n32) );
  CLKINVX20 U66 ( .A(n32), .Y(mem_wdata_D[51]) );
  INVX4 U67 ( .A(n404), .Y(n34) );
  CLKINVX20 U68 ( .A(n34), .Y(mem_wdata_D[9]) );
  INVX4 U69 ( .A(n362), .Y(n36) );
  CLKINVX20 U70 ( .A(n36), .Y(mem_wdata_D[52]) );
  INVX4 U71 ( .A(n331), .Y(n38) );
  CLKINVX20 U72 ( .A(n38), .Y(mem_wdata_D[83]) );
  INVX4 U73 ( .A(n403), .Y(n40) );
  CLKINVX20 U74 ( .A(n40), .Y(mem_wdata_D[10]) );
  INVX4 U75 ( .A(n361), .Y(n42) );
  CLKINVX20 U76 ( .A(n42), .Y(mem_wdata_D[53]) );
  INVX4 U77 ( .A(n330), .Y(n44) );
  CLKINVX20 U78 ( .A(n44), .Y(mem_wdata_D[84]) );
  INVX4 U79 ( .A(n402), .Y(n46) );
  CLKINVX20 U80 ( .A(n46), .Y(mem_wdata_D[11]) );
  INVX4 U81 ( .A(n360), .Y(n48) );
  CLKINVX20 U82 ( .A(n48), .Y(mem_wdata_D[54]) );
  INVX4 U83 ( .A(n329), .Y(n50) );
  CLKINVX20 U84 ( .A(n50), .Y(mem_wdata_D[85]) );
  INVX4 U85 ( .A(n401), .Y(n52) );
  CLKINVX20 U86 ( .A(n52), .Y(mem_wdata_D[12]) );
  INVX4 U87 ( .A(n359), .Y(n54) );
  CLKINVX20 U88 ( .A(n54), .Y(mem_wdata_D[55]) );
  INVX4 U89 ( .A(n328), .Y(n56) );
  CLKINVX20 U90 ( .A(n56), .Y(mem_wdata_D[86]) );
  INVX4 U91 ( .A(n400), .Y(n58) );
  CLKINVX20 U92 ( .A(n58), .Y(mem_wdata_D[13]) );
  INVX4 U93 ( .A(n358), .Y(n60) );
  CLKINVX20 U94 ( .A(n60), .Y(mem_wdata_D[56]) );
  INVX4 U95 ( .A(n327), .Y(n62) );
  CLKINVX20 U96 ( .A(n62), .Y(mem_wdata_D[87]) );
  INVX4 U97 ( .A(n399), .Y(n64) );
  CLKINVX20 U98 ( .A(n64), .Y(mem_wdata_D[14]) );
  INVX4 U99 ( .A(n357), .Y(n66) );
  CLKINVX20 U100 ( .A(n66), .Y(mem_wdata_D[57]) );
  INVX4 U101 ( .A(n326), .Y(n68) );
  CLKINVX20 U102 ( .A(n68), .Y(mem_wdata_D[88]) );
  INVX4 U103 ( .A(n398), .Y(n70) );
  CLKINVX20 U104 ( .A(n70), .Y(mem_wdata_D[15]) );
  INVX4 U105 ( .A(n356), .Y(n72) );
  CLKINVX20 U106 ( .A(n72), .Y(mem_wdata_D[58]) );
  INVX4 U107 ( .A(n325), .Y(n74) );
  CLKINVX20 U108 ( .A(n74), .Y(mem_wdata_D[89]) );
  INVX4 U109 ( .A(n397), .Y(n76) );
  CLKINVX20 U110 ( .A(n76), .Y(mem_wdata_D[16]) );
  INVX4 U111 ( .A(n355), .Y(n78) );
  CLKINVX20 U112 ( .A(n78), .Y(mem_wdata_D[59]) );
  INVX4 U113 ( .A(n324), .Y(n80) );
  CLKINVX20 U114 ( .A(n80), .Y(mem_wdata_D[90]) );
  INVX4 U115 ( .A(n396), .Y(n82) );
  CLKINVX20 U116 ( .A(n82), .Y(mem_wdata_D[17]) );
  INVX4 U117 ( .A(n354), .Y(n84) );
  CLKINVX20 U118 ( .A(n84), .Y(mem_wdata_D[60]) );
  INVX4 U119 ( .A(n323), .Y(n86) );
  CLKINVX20 U120 ( .A(n86), .Y(mem_wdata_D[91]) );
  INVX4 U121 ( .A(n395), .Y(n88) );
  CLKINVX20 U122 ( .A(n88), .Y(mem_wdata_D[18]) );
  INVX4 U123 ( .A(n353), .Y(n90) );
  CLKINVX20 U124 ( .A(n90), .Y(mem_wdata_D[61]) );
  INVX4 U125 ( .A(n322), .Y(n92) );
  CLKINVX20 U126 ( .A(n92), .Y(mem_wdata_D[92]) );
  INVX4 U127 ( .A(n394), .Y(n94) );
  CLKINVX20 U128 ( .A(n94), .Y(mem_wdata_D[19]) );
  INVX4 U129 ( .A(n352), .Y(n96) );
  CLKINVX20 U130 ( .A(n96), .Y(mem_wdata_D[62]) );
  INVX4 U131 ( .A(n321), .Y(n98) );
  CLKINVX20 U132 ( .A(n98), .Y(mem_wdata_D[93]) );
  INVX4 U133 ( .A(n393), .Y(n100) );
  CLKINVX20 U134 ( .A(n100), .Y(mem_wdata_D[20]) );
  INVX4 U135 ( .A(n351), .Y(n102) );
  CLKINVX20 U136 ( .A(n102), .Y(mem_wdata_D[63]) );
  INVX4 U137 ( .A(n320), .Y(n104) );
  CLKINVX20 U138 ( .A(n104), .Y(mem_wdata_D[94]) );
  INVX4 U139 ( .A(n392), .Y(n106) );
  CLKINVX20 U140 ( .A(n106), .Y(mem_wdata_D[21]) );
  INVX4 U141 ( .A(n350), .Y(n108) );
  CLKINVX20 U142 ( .A(n108), .Y(mem_wdata_D[64]) );
  INVX4 U143 ( .A(n319), .Y(n110) );
  CLKINVX20 U144 ( .A(n110), .Y(mem_wdata_D[95]) );
  INVX4 U145 ( .A(n391), .Y(n112) );
  CLKINVX20 U146 ( .A(n112), .Y(mem_wdata_D[22]) );
  INVX4 U147 ( .A(n349), .Y(n114) );
  CLKINVX20 U148 ( .A(n114), .Y(mem_wdata_D[65]) );
  INVX4 U149 ( .A(n318), .Y(n116) );
  CLKINVX20 U150 ( .A(n116), .Y(mem_wdata_D[96]) );
  INVX4 U151 ( .A(n390), .Y(n118) );
  CLKINVX20 U152 ( .A(n118), .Y(mem_wdata_D[23]) );
  INVX4 U153 ( .A(n348), .Y(n120) );
  CLKINVX20 U154 ( .A(n120), .Y(mem_wdata_D[66]) );
  INVX4 U155 ( .A(n317), .Y(n122) );
  CLKINVX20 U156 ( .A(n122), .Y(mem_wdata_D[97]) );
  INVX4 U157 ( .A(n389), .Y(n124) );
  CLKINVX20 U158 ( .A(n124), .Y(mem_wdata_D[24]) );
  INVX4 U159 ( .A(n347), .Y(n126) );
  CLKINVX20 U160 ( .A(n126), .Y(mem_wdata_D[67]) );
  INVX4 U161 ( .A(n316), .Y(n128) );
  CLKINVX20 U162 ( .A(n128), .Y(mem_wdata_D[98]) );
  INVX4 U163 ( .A(n388), .Y(n130) );
  CLKINVX20 U164 ( .A(n130), .Y(mem_wdata_D[25]) );
  INVX4 U165 ( .A(n346), .Y(n132) );
  CLKINVX20 U166 ( .A(n132), .Y(mem_wdata_D[68]) );
  INVX4 U167 ( .A(n315), .Y(n134) );
  CLKINVX20 U168 ( .A(n134), .Y(mem_wdata_D[99]) );
  INVX4 U169 ( .A(n387), .Y(n136) );
  CLKINVX20 U170 ( .A(n136), .Y(mem_wdata_D[26]) );
  INVX4 U171 ( .A(n345), .Y(n138) );
  CLKINVX20 U172 ( .A(n138), .Y(mem_wdata_D[69]) );
  INVX4 U173 ( .A(n314), .Y(n140) );
  CLKINVX20 U174 ( .A(n140), .Y(mem_wdata_D[100]) );
  INVX4 U175 ( .A(n386), .Y(n142) );
  CLKINVX20 U176 ( .A(n142), .Y(mem_wdata_D[27]) );
  INVX4 U177 ( .A(n344), .Y(n144) );
  CLKINVX20 U178 ( .A(n144), .Y(mem_wdata_D[70]) );
  INVX4 U179 ( .A(n313), .Y(n146) );
  CLKINVX20 U180 ( .A(n146), .Y(mem_wdata_D[101]) );
  INVX4 U181 ( .A(n385), .Y(n148) );
  CLKINVX20 U182 ( .A(n148), .Y(mem_wdata_D[28]) );
  INVX4 U183 ( .A(n312), .Y(n150) );
  CLKINVX20 U184 ( .A(n150), .Y(mem_wdata_D[102]) );
  INVX4 U185 ( .A(n384), .Y(n152) );
  CLKINVX20 U186 ( .A(n152), .Y(mem_wdata_D[29]) );
  INVX4 U187 ( .A(n311), .Y(n154) );
  CLKINVX20 U188 ( .A(n154), .Y(mem_wdata_D[103]) );
  INVX4 U189 ( .A(n383), .Y(n156) );
  CLKINVX20 U190 ( .A(n156), .Y(mem_wdata_D[30]) );
  INVX4 U191 ( .A(n310), .Y(n158) );
  CLKINVX20 U192 ( .A(n158), .Y(mem_wdata_D[104]) );
  INVX4 U193 ( .A(n382), .Y(n160) );
  CLKINVX20 U194 ( .A(n160), .Y(mem_wdata_D[31]) );
  INVX4 U195 ( .A(n309), .Y(n162) );
  CLKINVX20 U196 ( .A(n162), .Y(mem_wdata_D[105]) );
  INVX4 U197 ( .A(n308), .Y(n164) );
  CLKINVX20 U198 ( .A(n164), .Y(mem_wdata_D[106]) );
  INVX4 U199 ( .A(n307), .Y(n166) );
  CLKINVX20 U200 ( .A(n166), .Y(mem_wdata_D[107]) );
  INVX4 U201 ( .A(n410), .Y(n168) );
  CLKINVX20 U202 ( .A(n168), .Y(mem_addr_I[4]) );
  INVX4 U203 ( .A(n287), .Y(n170) );
  CLKINVX20 U204 ( .A(n170), .Y(mem_addr_D[6]) );
  CLKINVX6 U205 ( .A(n411), .Y(n172) );
  INVX20 U206 ( .A(n172), .Y(mem_wdata_I[127]) );
  INVX20 U207 ( .A(n174), .Y(mem_addr_D[24]) );
  INVX20 U208 ( .A(n176), .Y(mem_addr_D[28]) );
  CLKINVX6 U209 ( .A(n414), .Y(n178) );
  INVX20 U210 ( .A(n178), .Y(mem_wdata_I[81]) );
  CLKINVX6 U211 ( .A(n413), .Y(n180) );
  INVX20 U212 ( .A(n180), .Y(mem_wdata_I[82]) );
  CLKINVX6 U213 ( .A(n412), .Y(n182) );
  INVX20 U214 ( .A(n182), .Y(mem_wdata_I[83]) );
  INVX3 U215 ( .A(n306), .Y(n188) );
  INVX16 U216 ( .A(n188), .Y(mem_wdata_D[109]) );
  INVX3 U217 ( .A(n305), .Y(n194) );
  INVX16 U218 ( .A(n194), .Y(mem_wdata_D[110]) );
  INVX3 U219 ( .A(n304), .Y(n200) );
  INVX16 U220 ( .A(n200), .Y(mem_wdata_D[111]) );
  INVX3 U221 ( .A(n303), .Y(n206) );
  INVX16 U222 ( .A(n206), .Y(mem_wdata_D[112]) );
  INVX3 U223 ( .A(n302), .Y(n214) );
  INVX16 U224 ( .A(n214), .Y(mem_wdata_D[113]) );
  INVX3 U225 ( .A(n301), .Y(n222) );
  INVX16 U226 ( .A(n222), .Y(mem_wdata_D[114]) );
  INVX3 U227 ( .A(n300), .Y(n230) );
  INVX16 U228 ( .A(n230), .Y(mem_wdata_D[115]) );
  INVX3 U229 ( .A(n299), .Y(n238) );
  INVX16 U230 ( .A(n238), .Y(mem_wdata_D[116]) );
  INVX3 U231 ( .A(n298), .Y(n246) );
  INVX16 U232 ( .A(n246), .Y(mem_wdata_D[117]) );
  INVX3 U233 ( .A(n297), .Y(n254) );
  INVX16 U234 ( .A(n254), .Y(mem_wdata_D[118]) );
  INVX3 U235 ( .A(n296), .Y(n262) );
  INVX16 U236 ( .A(n262), .Y(mem_wdata_D[119]) );
  INVX3 U237 ( .A(n295), .Y(n270) );
  INVX16 U238 ( .A(n270), .Y(mem_wdata_D[120]) );
  INVXL U239 ( .A(n277), .Y(n278) );
  BUFX12 U240 ( .A(n3), .Y(DCACHE_addr[3]) );
  BUFX16 U241 ( .A(rst_n), .Y(n277) );
  BUFX12 U242 ( .A(n280), .Y(mem_write_D) );
  BUFX12 U243 ( .A(n409), .Y(mem_write_I) );
  BUFX12 U244 ( .A(n279), .Y(mem_read_D) );
  BUFX12 U245 ( .A(n408), .Y(mem_read_I) );
  INVX12 U246 ( .A(n208), .Y(mem_wdata_D[0]) );
  INVX1 U247 ( .A(n407), .Y(n208) );
  INVX12 U248 ( .A(n216), .Y(mem_wdata_D[121]) );
  INVX12 U249 ( .A(n224), .Y(mem_wdata_D[122]) );
  INVX12 U250 ( .A(n232), .Y(mem_wdata_D[123]) );
  INVX12 U251 ( .A(n240), .Y(mem_wdata_D[124]) );
  INVX12 U252 ( .A(n248), .Y(mem_wdata_D[125]) );
  INVX12 U253 ( .A(n256), .Y(mem_wdata_D[126]) );
  INVX12 U254 ( .A(n264), .Y(mem_wdata_D[127]) );
  INVX12 U255 ( .A(n184), .Y(mem_wdata_D[33]) );
  INVX12 U256 ( .A(n190), .Y(mem_wdata_D[34]) );
  INVX12 U257 ( .A(n196), .Y(mem_wdata_D[35]) );
  INVX12 U258 ( .A(n202), .Y(mem_wdata_D[36]) );
  INVX12 U259 ( .A(n210), .Y(mem_wdata_D[38]) );
  INVX12 U260 ( .A(n218), .Y(mem_wdata_D[39]) );
  INVX12 U261 ( .A(n226), .Y(mem_wdata_D[40]) );
  INVX12 U262 ( .A(n234), .Y(mem_wdata_D[41]) );
  INVX12 U263 ( .A(n242), .Y(mem_wdata_D[42]) );
  INVX12 U264 ( .A(n250), .Y(mem_wdata_D[43]) );
  INVX12 U265 ( .A(n258), .Y(mem_wdata_D[44]) );
  INVX12 U266 ( .A(n266), .Y(mem_wdata_D[45]) );
  INVX12 U267 ( .A(n186), .Y(mem_wdata_D[71]) );
  INVX12 U268 ( .A(n192), .Y(mem_wdata_D[72]) );
  INVX12 U269 ( .A(n198), .Y(mem_wdata_D[73]) );
  INVX12 U270 ( .A(n204), .Y(mem_wdata_D[74]) );
  INVX12 U271 ( .A(n212), .Y(mem_wdata_D[75]) );
  INVX12 U272 ( .A(n220), .Y(mem_wdata_D[76]) );
  INVX12 U273 ( .A(n228), .Y(mem_wdata_D[77]) );
  INVX12 U274 ( .A(n236), .Y(mem_wdata_D[78]) );
  INVX12 U275 ( .A(n244), .Y(mem_wdata_D[79]) );
  INVX12 U276 ( .A(n252), .Y(mem_wdata_D[80]) );
  INVX12 U277 ( .A(n260), .Y(mem_wdata_D[81]) );
  INVX12 U278 ( .A(n268), .Y(mem_wdata_D[82]) );
endmodule

