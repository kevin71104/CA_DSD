
module IF_DEC_regFile ( clk, rst_n, flush, stallcache, stall_lw_use, 
        instruction_next, PCplus4, branchOffset, opcode, Rs, Rt, Rd, shamt, 
        funct, immediate, instruction_regI, PCplus4_regI );
  input [31:0] instruction_next;
  input [31:0] PCplus4;
  output [15:0] branchOffset;
  output [5:0] opcode;
  output [4:0] Rs;
  output [4:0] Rt;
  output [4:0] Rd;
  output [4:0] shamt;
  output [5:0] funct;
  output [15:0] immediate;
  output [31:0] instruction_regI;
  output [31:0] PCplus4_regI;
  input clk, rst_n, flush, stallcache, stall_lw_use;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n1, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154;

  DFFRX4 \instruction_regI_reg[31]  ( .D(n34), .CK(clk), .RN(n132), .Q(
        opcode[5]) );
  DFFRX4 \instruction_regI_reg[29]  ( .D(n32), .CK(clk), .RN(n132), .Q(
        opcode[3]) );
  DFFRX4 \instruction_regI_reg[28]  ( .D(n31), .CK(clk), .RN(n132), .Q(
        opcode[2]) );
  DFFRX4 \instruction_regI_reg[27]  ( .D(n30), .CK(clk), .RN(n132), .Q(
        opcode[1]) );
  DFFRX4 \instruction_regI_reg[25]  ( .D(n28), .CK(clk), .RN(n132), .Q(Rs[4])
         );
  DFFRX4 \instruction_regI_reg[22]  ( .D(n25), .CK(clk), .RN(n131), .Q(Rs[1])
         );
  DFFRX1 \PCplus4_regI_reg[31]  ( .D(n66), .CK(clk), .RN(n135), .Q(
        PCplus4_regI[31]) );
  DFFRX1 \PCplus4_regI_reg[30]  ( .D(n65), .CK(clk), .RN(n135), .Q(
        PCplus4_regI[30]) );
  DFFRX1 \PCplus4_regI_reg[29]  ( .D(n64), .CK(clk), .RN(n135), .Q(
        PCplus4_regI[29]) );
  DFFRX1 \PCplus4_regI_reg[28]  ( .D(n63), .CK(clk), .RN(n135), .Q(
        PCplus4_regI[28]) );
  DFFRX1 \PCplus4_regI_reg[27]  ( .D(n62), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[27]) );
  DFFRX1 \PCplus4_regI_reg[26]  ( .D(n61), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[26]) );
  DFFRX1 \PCplus4_regI_reg[25]  ( .D(n60), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[25]) );
  DFFRX1 \PCplus4_regI_reg[24]  ( .D(n59), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[24]) );
  DFFRX1 \instruction_regI_reg[30]  ( .D(n33), .CK(clk), .RN(n132), .Q(
        opcode[4]) );
  DFFRX2 \instruction_regI_reg[5]  ( .D(n8), .CK(clk), .RN(n130), .Q(funct[5])
         );
  DFFRX2 \instruction_regI_reg[2]  ( .D(n5), .CK(clk), .RN(n130), .Q(funct[2])
         );
  DFFRX2 \instruction_regI_reg[4]  ( .D(n7), .CK(clk), .RN(n130), .Q(funct[4])
         );
  DFFRX2 \instruction_regI_reg[0]  ( .D(n3), .CK(clk), .RN(n130), .Q(funct[0])
         );
  DFFRX2 \instruction_regI_reg[3]  ( .D(n6), .CK(clk), .RN(n130), .Q(funct[3])
         );
  DFFRX2 \instruction_regI_reg[26]  ( .D(n29), .CK(clk), .RN(n132), .Q(
        opcode[0]) );
  DFFRX2 \instruction_regI_reg[1]  ( .D(n4), .CK(clk), .RN(n130), .Q(funct[1])
         );
  DFFRX1 \instruction_regI_reg[9]  ( .D(n12), .CK(clk), .RN(n130), .Q(shamt[3]) );
  DFFRX1 \instruction_regI_reg[8]  ( .D(n11), .CK(clk), .RN(n130), .Q(shamt[2]) );
  DFFRX1 \instruction_regI_reg[7]  ( .D(n10), .CK(clk), .RN(n130), .Q(shamt[1]) );
  DFFRX1 \instruction_regI_reg[6]  ( .D(n9), .CK(clk), .RN(n130), .Q(shamt[0])
         );
  DFFRX1 \instruction_regI_reg[14]  ( .D(n17), .CK(clk), .RN(n131), .Q(Rd[3])
         );
  DFFRX1 \instruction_regI_reg[13]  ( .D(n16), .CK(clk), .RN(n131), .Q(Rd[2])
         );
  DFFRX1 \instruction_regI_reg[12]  ( .D(n15), .CK(clk), .RN(n131), .Q(Rd[1])
         );
  DFFRX1 \instruction_regI_reg[15]  ( .D(n18), .CK(clk), .RN(n131), .Q(Rd[4])
         );
  DFFRX1 \instruction_regI_reg[10]  ( .D(n13), .CK(clk), .RN(n130), .Q(
        shamt[4]) );
  DFFRX1 \instruction_regI_reg[16]  ( .D(n19), .CK(clk), .RN(n131), .Q(Rt[0])
         );
  DFFRX2 \PCplus4_regI_reg[16]  ( .D(n51), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[16]) );
  DFFRX2 \PCplus4_regI_reg[1]  ( .D(n36), .CK(clk), .RN(n132), .Q(
        PCplus4_regI[1]) );
  DFFRX2 \PCplus4_regI_reg[2]  ( .D(n37), .CK(clk), .RN(n132), .Q(
        PCplus4_regI[2]) );
  DFFRX2 \PCplus4_regI_reg[4]  ( .D(n39), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[4]) );
  DFFRX4 \instruction_regI_reg[17]  ( .D(n20), .CK(clk), .RN(n131), .Q(Rt[1])
         );
  DFFRX4 \instruction_regI_reg[21]  ( .D(n24), .CK(clk), .RN(n131), .Q(Rs[0])
         );
  DFFRX4 \instruction_regI_reg[23]  ( .D(n26), .CK(clk), .RN(n131), .Q(Rs[2])
         );
  DFFRX4 \instruction_regI_reg[19]  ( .D(n22), .CK(clk), .RN(n131), .Q(Rt[3])
         );
  DFFRX4 \instruction_regI_reg[24]  ( .D(n27), .CK(clk), .RN(n132), .Q(Rs[3])
         );
  DFFRX4 \instruction_regI_reg[18]  ( .D(n21), .CK(clk), .RN(n131), .Q(Rt[2])
         );
  DFFRX4 \instruction_regI_reg[20]  ( .D(n23), .CK(clk), .RN(n131), .Q(Rt[4])
         );
  DFFRX2 \PCplus4_regI_reg[6]  ( .D(n41), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[6]) );
  DFFRX2 \PCplus4_regI_reg[7]  ( .D(n42), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[7]) );
  DFFRX2 \PCplus4_regI_reg[9]  ( .D(n44), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[9]) );
  DFFRX2 \PCplus4_regI_reg[23]  ( .D(n58), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[23]) );
  DFFRX2 \PCplus4_regI_reg[5]  ( .D(n40), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[5]) );
  DFFRX2 \PCplus4_regI_reg[17]  ( .D(n52), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[17]) );
  DFFRX2 \PCplus4_regI_reg[15]  ( .D(n50), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[15]) );
  DFFRX2 \PCplus4_regI_reg[21]  ( .D(n56), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[21]) );
  DFFRX2 \PCplus4_regI_reg[13]  ( .D(n48), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[13]) );
  DFFRX2 \PCplus4_regI_reg[11]  ( .D(n46), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[11]) );
  DFFRX2 \PCplus4_regI_reg[10]  ( .D(n45), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[10]) );
  DFFRX2 \PCplus4_regI_reg[8]  ( .D(n43), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[8]) );
  DFFRX2 \PCplus4_regI_reg[12]  ( .D(n47), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[12]) );
  DFFRX2 \PCplus4_regI_reg[14]  ( .D(n49), .CK(clk), .RN(n133), .Q(
        PCplus4_regI[14]) );
  DFFRX2 \PCplus4_regI_reg[0]  ( .D(n35), .CK(clk), .RN(n132), .Q(
        PCplus4_regI[0]) );
  DFFRX2 \PCplus4_regI_reg[3]  ( .D(n38), .CK(clk), .RN(n132), .Q(
        PCplus4_regI[3]) );
  DFFRX2 \PCplus4_regI_reg[18]  ( .D(n53), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[18]) );
  DFFRX2 \PCplus4_regI_reg[19]  ( .D(n54), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[19]) );
  DFFRX2 \PCplus4_regI_reg[20]  ( .D(n55), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[20]) );
  DFFRX2 \PCplus4_regI_reg[22]  ( .D(n57), .CK(clk), .RN(n134), .Q(
        PCplus4_regI[22]) );
  DFFRX2 \instruction_regI_reg[11]  ( .D(n14), .CK(clk), .RN(n130), .Q(Rd[0])
         );
  BUFX20 U2 ( .A(n1), .Y(n145) );
  BUFX20 U3 ( .A(n145), .Y(n144) );
  AO22XL U4 ( .A0(instruction_next[11]), .A1(n149), .B0(Rd[0]), .B1(n141), .Y(
        n14) );
  AO22X1 U5 ( .A0(instruction_next[0]), .A1(n148), .B0(funct[0]), .B1(n140), 
        .Y(n3) );
  AO22X2 U6 ( .A0(instruction_next[4]), .A1(n149), .B0(funct[4]), .B1(n141), 
        .Y(n7) );
  AO22X2 U7 ( .A0(instruction_next[2]), .A1(n148), .B0(funct[2]), .B1(n140), 
        .Y(n5) );
  AO22X2 U8 ( .A0(instruction_next[5]), .A1(n149), .B0(funct[5]), .B1(n141), 
        .Y(n8) );
  CLKBUFX2 U9 ( .A(rst_n), .Y(n137) );
  CLKBUFX2 U10 ( .A(rst_n), .Y(n136) );
  CLKAND2X6 U11 ( .A(n153), .B(n152), .Y(n1) );
  AO22X1 U12 ( .A0(instruction_next[27]), .A1(n150), .B0(opcode[1]), .B1(n142), 
        .Y(n30) );
  AO22X4 U13 ( .A0(instruction_next[31]), .A1(n151), .B0(opcode[5]), .B1(n143), 
        .Y(n34) );
  AO22X4 U14 ( .A0(instruction_next[28]), .A1(n151), .B0(opcode[2]), .B1(n143), 
        .Y(n31) );
  BUFX20 U15 ( .A(n144), .Y(n151) );
  AO22X4 U16 ( .A0(instruction_next[10]), .A1(n149), .B0(shamt[4]), .B1(n141), 
        .Y(n13) );
  AO22X4 U17 ( .A0(instruction_next[8]), .A1(n149), .B0(shamt[2]), .B1(n141), 
        .Y(n11) );
  AO22X4 U18 ( .A0(instruction_next[9]), .A1(n149), .B0(shamt[3]), .B1(n141), 
        .Y(n12) );
  AO22X4 U19 ( .A0(instruction_next[7]), .A1(n149), .B0(shamt[1]), .B1(n141), 
        .Y(n10) );
  AO22X4 U20 ( .A0(instruction_next[13]), .A1(n149), .B0(Rd[2]), .B1(n141), 
        .Y(n16) );
  AO22X4 U21 ( .A0(instruction_next[15]), .A1(n149), .B0(Rd[4]), .B1(n141), 
        .Y(n18) );
  AO22X4 U22 ( .A0(instruction_next[6]), .A1(n149), .B0(shamt[0]), .B1(n141), 
        .Y(n9) );
  AO22X4 U23 ( .A0(instruction_next[14]), .A1(n149), .B0(Rd[3]), .B1(n141), 
        .Y(n17) );
  AO22X4 U24 ( .A0(instruction_next[3]), .A1(n148), .B0(funct[3]), .B1(n140), 
        .Y(n6) );
  AO22X4 U25 ( .A0(PCplus4[4]), .A1(n146), .B0(PCplus4_regI[4]), .B1(n138), 
        .Y(n39) );
  AO22X4 U26 ( .A0(PCplus4[2]), .A1(n146), .B0(PCplus4_regI[2]), .B1(n138), 
        .Y(n37) );
  AO22X4 U27 ( .A0(PCplus4[1]), .A1(n146), .B0(PCplus4_regI[1]), .B1(n138), 
        .Y(n36) );
  AO22X4 U28 ( .A0(PCplus4[16]), .A1(n147), .B0(PCplus4_regI[16]), .B1(n139), 
        .Y(n51) );
  BUFX20 U29 ( .A(n144), .Y(n150) );
  BUFX20 U30 ( .A(n141), .Y(n142) );
  BUFX20 U31 ( .A(n144), .Y(n146) );
  AO22X4 U32 ( .A0(PCplus4[30]), .A1(n148), .B0(PCplus4_regI[30]), .B1(n140), 
        .Y(n65) );
  AO22X4 U33 ( .A0(PCplus4[24]), .A1(n148), .B0(PCplus4_regI[24]), .B1(n140), 
        .Y(n59) );
  AO22X4 U34 ( .A0(PCplus4[26]), .A1(n148), .B0(PCplus4_regI[26]), .B1(n140), 
        .Y(n61) );
  AO22X4 U35 ( .A0(PCplus4[27]), .A1(n148), .B0(PCplus4_regI[27]), .B1(n140), 
        .Y(n62) );
  AO22X4 U36 ( .A0(PCplus4[25]), .A1(n148), .B0(PCplus4_regI[25]), .B1(n140), 
        .Y(n60) );
  AO22X4 U37 ( .A0(PCplus4[31]), .A1(n148), .B0(PCplus4_regI[31]), .B1(n140), 
        .Y(n66) );
  AO22X4 U38 ( .A0(PCplus4[28]), .A1(n148), .B0(PCplus4_regI[28]), .B1(n140), 
        .Y(n63) );
  AO22X4 U39 ( .A0(instruction_next[1]), .A1(n148), .B0(funct[1]), .B1(n140), 
        .Y(n4) );
  BUFX20 U40 ( .A(n145), .Y(n148) );
  BUFX20 U41 ( .A(n141), .Y(n143) );
  BUFX20 U42 ( .A(n144), .Y(n147) );
  BUFX20 U43 ( .A(n140), .Y(n138) );
  AO22X4 U44 ( .A0(PCplus4[0]), .A1(n146), .B0(PCplus4_regI[0]), .B1(n138), 
        .Y(n35) );
  AO22X4 U45 ( .A0(PCplus4[8]), .A1(n146), .B0(PCplus4_regI[8]), .B1(n138), 
        .Y(n43) );
  BUFX20 U46 ( .A(n145), .Y(n149) );
  AO22XL U47 ( .A0(instruction_next[12]), .A1(n149), .B0(Rd[1]), .B1(n141), 
        .Y(n15) );
  AO22X4 U48 ( .A0(PCplus4[3]), .A1(n146), .B0(PCplus4_regI[3]), .B1(n138), 
        .Y(n38) );
  AO22X4 U49 ( .A0(PCplus4[10]), .A1(n146), .B0(PCplus4_regI[10]), .B1(n138), 
        .Y(n45) );
  AO22X4 U50 ( .A0(PCplus4[11]), .A1(n146), .B0(PCplus4_regI[11]), .B1(n138), 
        .Y(n46) );
  AO22X4 U51 ( .A0(PCplus4[7]), .A1(n146), .B0(PCplus4_regI[7]), .B1(n138), 
        .Y(n42) );
  AO22X4 U52 ( .A0(PCplus4[9]), .A1(n146), .B0(PCplus4_regI[9]), .B1(n138), 
        .Y(n44) );
  AO22X4 U53 ( .A0(PCplus4[5]), .A1(n146), .B0(PCplus4_regI[5]), .B1(n138), 
        .Y(n40) );
  AO22X4 U54 ( .A0(PCplus4[6]), .A1(n146), .B0(PCplus4_regI[6]), .B1(n138), 
        .Y(n41) );
  BUFX20 U55 ( .A(n140), .Y(n139) );
  AO22X4 U56 ( .A0(PCplus4[12]), .A1(n147), .B0(PCplus4_regI[12]), .B1(n139), 
        .Y(n47) );
  BUFX20 U57 ( .A(n154), .Y(n141) );
  BUFX20 U58 ( .A(n154), .Y(n140) );
  AO22X4 U59 ( .A0(PCplus4[23]), .A1(n147), .B0(PCplus4_regI[23]), .B1(n139), 
        .Y(n58) );
  AO22X4 U60 ( .A0(PCplus4[13]), .A1(n147), .B0(PCplus4_regI[13]), .B1(n139), 
        .Y(n48) );
  AO22X4 U61 ( .A0(PCplus4[14]), .A1(n147), .B0(PCplus4_regI[14]), .B1(n139), 
        .Y(n49) );
  AO22X4 U62 ( .A0(PCplus4[15]), .A1(n147), .B0(PCplus4_regI[15]), .B1(n139), 
        .Y(n50) );
  AO22X4 U63 ( .A0(PCplus4[17]), .A1(n147), .B0(PCplus4_regI[17]), .B1(n139), 
        .Y(n52) );
  AO22X4 U64 ( .A0(PCplus4[18]), .A1(n147), .B0(PCplus4_regI[18]), .B1(n139), 
        .Y(n53) );
  AO22X4 U65 ( .A0(PCplus4[19]), .A1(n147), .B0(PCplus4_regI[19]), .B1(n139), 
        .Y(n54) );
  AO22X4 U66 ( .A0(PCplus4[20]), .A1(n147), .B0(PCplus4_regI[20]), .B1(n139), 
        .Y(n55) );
  AO22X4 U67 ( .A0(PCplus4[21]), .A1(n147), .B0(PCplus4_regI[21]), .B1(n139), 
        .Y(n56) );
  AO22X4 U68 ( .A0(PCplus4[22]), .A1(n147), .B0(PCplus4_regI[22]), .B1(n139), 
        .Y(n57) );
  AO22X4 U69 ( .A0(instruction_next[29]), .A1(n151), .B0(opcode[3]), .B1(n143), 
        .Y(n32) );
  CLKBUFX3 U70 ( .A(shamt[4]), .Y(instruction_regI[10]) );
  CLKBUFX3 U71 ( .A(Rd[0]), .Y(instruction_regI[11]) );
  CLKBUFX3 U72 ( .A(Rd[1]), .Y(instruction_regI[12]) );
  CLKBUFX3 U73 ( .A(Rd[2]), .Y(instruction_regI[13]) );
  CLKBUFX3 U74 ( .A(Rd[3]), .Y(instruction_regI[14]) );
  CLKBUFX3 U75 ( .A(Rd[4]), .Y(instruction_regI[15]) );
  CLKBUFX3 U76 ( .A(shamt[0]), .Y(instruction_regI[6]) );
  CLKBUFX3 U77 ( .A(shamt[1]), .Y(instruction_regI[7]) );
  CLKBUFX3 U78 ( .A(shamt[2]), .Y(instruction_regI[8]) );
  CLKBUFX3 U79 ( .A(shamt[3]), .Y(instruction_regI[9]) );
  CLKBUFX2 U80 ( .A(Rt[0]), .Y(instruction_regI[16]) );
  CLKBUFX2 U81 ( .A(Rt[1]), .Y(instruction_regI[17]) );
  CLKBUFX2 U82 ( .A(Rs[0]), .Y(instruction_regI[21]) );
  CLKBUFX2 U83 ( .A(opcode[4]), .Y(instruction_regI[30]) );
  CLKBUFX2 U84 ( .A(funct[3]), .Y(instruction_regI[3]) );
  CLKBUFX2 U85 ( .A(Rt[2]), .Y(instruction_regI[18]) );
  CLKBUFX2 U86 ( .A(Rt[3]), .Y(instruction_regI[19]) );
  CLKBUFX2 U87 ( .A(Rt[4]), .Y(instruction_regI[20]) );
  CLKBUFX2 U88 ( .A(Rs[2]), .Y(instruction_regI[23]) );
  CLKBUFX2 U89 ( .A(Rs[3]), .Y(instruction_regI[24]) );
  CLKBUFX2 U90 ( .A(opcode[0]), .Y(instruction_regI[26]) );
  CLKBUFX2 U91 ( .A(funct[1]), .Y(instruction_regI[1]) );
  CLKBUFX2 U92 ( .A(funct[4]), .Y(instruction_regI[4]) );
  CLKBUFX2 U93 ( .A(funct[2]), .Y(instruction_regI[2]) );
  CLKBUFX2 U94 ( .A(funct[5]), .Y(instruction_regI[5]) );
  CLKBUFX2 U95 ( .A(funct[0]), .Y(instruction_regI[0]) );
  CLKBUFX2 U96 ( .A(opcode[1]), .Y(instruction_regI[27]) );
  CLKBUFX2 U97 ( .A(opcode[3]), .Y(instruction_regI[29]) );
  CLKBUFX2 U98 ( .A(opcode[5]), .Y(instruction_regI[31]) );
  CLKBUFX2 U99 ( .A(opcode[2]), .Y(instruction_regI[28]) );
  CLKBUFX2 U100 ( .A(Rs[1]), .Y(instruction_regI[22]) );
  CLKBUFX2 U101 ( .A(Rs[4]), .Y(instruction_regI[25]) );
  INVX6 U102 ( .A(n153), .Y(n154) );
  INVX3 U103 ( .A(flush), .Y(n152) );
  CLKBUFX2 U104 ( .A(funct[1]), .Y(branchOffset[1]) );
  CLKBUFX2 U105 ( .A(funct[0]), .Y(immediate[0]) );
  CLKBUFX2 U106 ( .A(funct[0]), .Y(branchOffset[0]) );
  CLKBUFX3 U107 ( .A(n137), .Y(n130) );
  CLKBUFX3 U108 ( .A(n137), .Y(n131) );
  CLKBUFX3 U109 ( .A(n137), .Y(n132) );
  CLKBUFX3 U110 ( .A(n136), .Y(n133) );
  CLKBUFX3 U111 ( .A(n136), .Y(n134) );
  CLKBUFX3 U112 ( .A(n136), .Y(n135) );
  AO22X1 U113 ( .A0(instruction_next[16]), .A1(n150), .B0(Rt[0]), .B1(n142), 
        .Y(n19) );
  AO22X1 U114 ( .A0(instruction_next[17]), .A1(n150), .B0(Rt[1]), .B1(n142), 
        .Y(n20) );
  AO22X1 U115 ( .A0(instruction_next[18]), .A1(n150), .B0(Rt[2]), .B1(n142), 
        .Y(n21) );
  AO22X1 U116 ( .A0(instruction_next[19]), .A1(n150), .B0(Rt[3]), .B1(n142), 
        .Y(n22) );
  AO22X1 U117 ( .A0(instruction_next[20]), .A1(n150), .B0(Rt[4]), .B1(n142), 
        .Y(n23) );
  AO22X1 U118 ( .A0(instruction_next[21]), .A1(n150), .B0(Rs[0]), .B1(n142), 
        .Y(n24) );
  AO22X1 U119 ( .A0(instruction_next[22]), .A1(n150), .B0(Rs[1]), .B1(n142), 
        .Y(n25) );
  AO22X1 U120 ( .A0(instruction_next[23]), .A1(n150), .B0(Rs[2]), .B1(n142), 
        .Y(n26) );
  AO22X1 U121 ( .A0(instruction_next[24]), .A1(n150), .B0(Rs[3]), .B1(n142), 
        .Y(n27) );
  AO22X1 U122 ( .A0(instruction_next[25]), .A1(n150), .B0(Rs[4]), .B1(n142), 
        .Y(n28) );
  AO22XL U123 ( .A0(instruction_next[26]), .A1(n150), .B0(opcode[0]), .B1(n142), .Y(n29) );
  AO22XL U124 ( .A0(instruction_next[30]), .A1(n151), .B0(opcode[4]), .B1(n143), .Y(n33) );
  AO22XL U125 ( .A0(PCplus4[29]), .A1(n148), .B0(PCplus4_regI[29]), .B1(n140), 
        .Y(n64) );
  CLKBUFX3 U126 ( .A(funct[1]), .Y(immediate[1]) );
  CLKBUFX3 U127 ( .A(Rd[4]), .Y(immediate[15]) );
  CLKBUFX3 U128 ( .A(Rd[4]), .Y(branchOffset[15]) );
  CLKBUFX3 U129 ( .A(Rd[3]), .Y(immediate[14]) );
  CLKBUFX3 U130 ( .A(Rd[3]), .Y(branchOffset[14]) );
  CLKBUFX3 U131 ( .A(Rd[2]), .Y(immediate[13]) );
  CLKBUFX3 U132 ( .A(Rd[2]), .Y(branchOffset[13]) );
  CLKBUFX3 U133 ( .A(Rd[1]), .Y(immediate[12]) );
  CLKBUFX3 U134 ( .A(Rd[1]), .Y(branchOffset[12]) );
  CLKBUFX3 U135 ( .A(Rd[0]), .Y(immediate[11]) );
  CLKBUFX3 U136 ( .A(Rd[0]), .Y(branchOffset[11]) );
  CLKBUFX3 U137 ( .A(shamt[4]), .Y(immediate[10]) );
  CLKBUFX3 U138 ( .A(shamt[4]), .Y(branchOffset[10]) );
  CLKBUFX3 U139 ( .A(shamt[3]), .Y(immediate[9]) );
  CLKBUFX3 U140 ( .A(shamt[3]), .Y(branchOffset[9]) );
  CLKBUFX3 U141 ( .A(shamt[2]), .Y(immediate[8]) );
  CLKBUFX3 U142 ( .A(shamt[2]), .Y(branchOffset[8]) );
  CLKBUFX3 U143 ( .A(shamt[1]), .Y(immediate[7]) );
  CLKBUFX3 U144 ( .A(shamt[1]), .Y(branchOffset[7]) );
  CLKBUFX3 U145 ( .A(shamt[0]), .Y(immediate[6]) );
  CLKBUFX3 U146 ( .A(shamt[0]), .Y(branchOffset[6]) );
  CLKBUFX3 U147 ( .A(funct[5]), .Y(immediate[5]) );
  CLKBUFX3 U148 ( .A(funct[5]), .Y(branchOffset[5]) );
  CLKBUFX3 U149 ( .A(funct[4]), .Y(immediate[4]) );
  CLKBUFX3 U150 ( .A(funct[4]), .Y(branchOffset[4]) );
  CLKBUFX3 U151 ( .A(funct[3]), .Y(immediate[3]) );
  CLKBUFX3 U152 ( .A(funct[3]), .Y(branchOffset[3]) );
  CLKBUFX3 U153 ( .A(funct[2]), .Y(immediate[2]) );
  CLKBUFX3 U154 ( .A(funct[2]), .Y(branchOffset[2]) );
  OAI21X4 U155 ( .A0(stall_lw_use), .A1(stallcache), .B0(n152), .Y(n153) );
endmodule


module DEC_EX_regFile ( clk, rst_n, stallcache, MemtoReg, ALUOp, JumpReg, 
        MemRead, MemWrite, ALUsrc, RegWrite, Branch, PCplus4_regI, funct, 
        branchOffset_D, A, B, ExtOut, Rs, Rt, wsel, MemtoReg_regD, ALUOp_regD, 
        MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, funct_regD, 
        A_regD, B_regD, ExtOut_regD, Rs_regD, Rt_regD, wsel_regD, JumpReg_regD, 
        Branch_regD, PCplus4_regD, branchOffset_regD );
  input [1:0] MemtoReg;
  input [5:0] ALUOp;
  input [31:0] PCplus4_regI;
  input [5:0] funct;
  input [15:0] branchOffset_D;
  input [31:0] A;
  input [31:0] B;
  input [31:0] ExtOut;
  input [4:0] Rs;
  input [4:0] Rt;
  input [4:0] wsel;
  output [1:0] MemtoReg_regD;
  output [5:0] ALUOp_regD;
  output [5:0] funct_regD;
  output [31:0] A_regD;
  output [31:0] B_regD;
  output [31:0] ExtOut_regD;
  output [4:0] Rs_regD;
  output [4:0] Rt_regD;
  output [4:0] wsel_regD;
  output [31:0] PCplus4_regD;
  output [15:0] branchOffset_regD;
  input clk, rst_n, stallcache, JumpReg, MemRead, MemWrite, ALUsrc, RegWrite,
         Branch;
  output MemRead_regD, MemWrite_regD, ALUsrc_regD, RegWrite_regD, JumpReg_regD,
         Branch_regD;
  wire   n2, n3, n14, n15, n16, n18, n19, n23, n27, n29, n31, n32, n33, n34,
         n35, n37, n38, n39, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n81, n82, n83, n84, n85, n87, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n108,
         n113, n115, n116, n117, n118, n119, n122, n123, n124, n125, n126,
         n132, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n170, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n10, n13, n21, n25, n26, n28, n30, n36, n40, n41, n42,
         n43, n44, n45, n53, n66, n79, n80, n86, n88, n89, n90, n91, n92, n105,
         n106, n107, n109, n110, n111, n112, n114, n120, n121, n127, n128,
         n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140,
         n167, n168, n169, n171, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453;

  DFFRX4 \funct_regD_reg[4]  ( .D(n305), .CK(clk), .RN(n40), .Q(funct_regD[4]), 
        .QN(n126) );
  DFFRX4 \funct_regD_reg[3]  ( .D(n304), .CK(clk), .RN(n40), .Q(funct_regD[3]), 
        .QN(n125) );
  DFFRX4 \funct_regD_reg[2]  ( .D(n303), .CK(clk), .RN(n40), .Q(funct_regD[2]), 
        .QN(n124) );
  DFFRX4 \funct_regD_reg[1]  ( .D(n302), .CK(clk), .RN(n40), .Q(funct_regD[1]), 
        .QN(n123) );
  DFFRX4 \funct_regD_reg[0]  ( .D(n301), .CK(clk), .RN(n40), .Q(funct_regD[0]), 
        .QN(n122) );
  DFFRX4 \ALUOp_regD_reg[5]  ( .D(n298), .CK(clk), .RN(n40), .Q(ALUOp_regD[5]), 
        .QN(n119) );
  DFFRX4 \ALUOp_regD_reg[4]  ( .D(n297), .CK(clk), .RN(n40), .Q(ALUOp_regD[4]), 
        .QN(n118) );
  DFFRX4 \ALUOp_regD_reg[3]  ( .D(n296), .CK(clk), .RN(n40), .Q(ALUOp_regD[3]), 
        .QN(n117) );
  DFFRX4 \ALUOp_regD_reg[2]  ( .D(n295), .CK(clk), .RN(n30), .Q(ALUOp_regD[2]), 
        .QN(n116) );
  DFFRX4 \ALUOp_regD_reg[1]  ( .D(n294), .CK(clk), .RN(n36), .Q(ALUOp_regD[1]), 
        .QN(n115) );
  DFFRX4 MemRead_regD_reg ( .D(n292), .CK(clk), .RN(n36), .Q(MemRead_regD), 
        .QN(n113) );
  DFFRX4 \A_regD_reg[9]  ( .D(n266), .CK(clk), .RN(n41), .Q(A_regD[9]), .QN(
        n87) );
  DFFRX4 \A_regD_reg[7]  ( .D(n264), .CK(clk), .RN(n41), .Q(A_regD[7]), .QN(
        n85) );
  DFFRX4 \A_regD_reg[6]  ( .D(n263), .CK(clk), .RN(n41), .Q(A_regD[6]), .QN(
        n84) );
  DFFRX4 \A_regD_reg[5]  ( .D(n262), .CK(clk), .RN(n41), .Q(A_regD[5]), .QN(
        n83) );
  DFFRX4 \A_regD_reg[4]  ( .D(n261), .CK(clk), .RN(n41), .Q(A_regD[4]), .QN(
        n82) );
  DFFRX4 \A_regD_reg[3]  ( .D(n260), .CK(clk), .RN(n41), .Q(A_regD[3]), .QN(
        n81) );
  DFFRX4 \ExtOut_regD_reg[5]  ( .D(n198), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[5]), .QN(n19) );
  DFFRX4 \ExtOut_regD_reg[4]  ( .D(n197), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[4]), .QN(n18) );
  DFFRX4 \ExtOut_regD_reg[2]  ( .D(n195), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[2]), .QN(n16) );
  DFFRX4 \ExtOut_regD_reg[1]  ( .D(n194), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[1]), .QN(n15) );
  DFFRX4 JumpReg_regD_reg ( .D(n177), .CK(clk), .RN(n80), .Q(JumpReg_regD), 
        .QN(n3) );
  DFFRX4 Branch_regD_reg ( .D(n176), .CK(clk), .RN(n80), .Q(Branch_regD), .QN(
        n2) );
  DFFRX1 MemWrite_regD_reg ( .D(n291), .CK(clk), .RN(n36), .Q(MemWrite_regD)
         );
  DFFRX1 \wsel_regD_reg[4]  ( .D(n182), .CK(clk), .RN(n80), .Q(wsel_regD[4])
         );
  DFFRX1 \wsel_regD_reg[2]  ( .D(n180), .CK(clk), .RN(n80), .Q(wsel_regD[2])
         );
  DFFRX1 \wsel_regD_reg[0]  ( .D(n178), .CK(clk), .RN(n80), .Q(wsel_regD[0])
         );
  DFFRX1 \wsel_regD_reg[3]  ( .D(n181), .CK(clk), .RN(n80), .Q(wsel_regD[3])
         );
  DFFRX1 \wsel_regD_reg[1]  ( .D(n179), .CK(clk), .RN(n80), .Q(wsel_regD[1])
         );
  DFFRX1 \PCplus4_regD_reg[31]  ( .D(n354), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[31]), .QN(n175) );
  DFFRX1 \branchOffset_regD_reg[14]  ( .D(n321), .CK(clk), .RN(n30), .Q(
        branchOffset_regD[14]), .QN(n142) );
  DFFRX1 \branchOffset_regD_reg[10]  ( .D(n317), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[10]) );
  DFFRX1 \branchOffset_regD_reg[6]  ( .D(n313), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[6]) );
  DFFRX1 \branchOffset_regD_reg[8]  ( .D(n315), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[8]) );
  DFFRX1 \branchOffset_regD_reg[9]  ( .D(n316), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[9]) );
  DFFRX1 \branchOffset_regD_reg[15]  ( .D(n322), .CK(clk), .RN(n30), .Q(
        branchOffset_regD[15]), .QN(n143) );
  DFFRX1 \branchOffset_regD_reg[13]  ( .D(n320), .CK(clk), .RN(n30), .Q(
        branchOffset_regD[13]), .QN(n141) );
  DFFRX1 \branchOffset_regD_reg[12]  ( .D(n319), .CK(clk), .RN(n26), .Q(
        branchOffset_regD[12]) );
  DFFRX1 \branchOffset_regD_reg[7]  ( .D(n314), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[7]) );
  DFFRX1 \branchOffset_regD_reg[5]  ( .D(n312), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[5]) );
  DFFRX1 \branchOffset_regD_reg[2]  ( .D(n309), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[2]) );
  DFFRX1 \branchOffset_regD_reg[11]  ( .D(n318), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[11]) );
  DFFRX1 \branchOffset_regD_reg[3]  ( .D(n310), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[3]) );
  DFFRX1 \branchOffset_regD_reg[4]  ( .D(n311), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[4]), .QN(n132) );
  DFFRX1 \branchOffset_regD_reg[1]  ( .D(n308), .CK(clk), .RN(n28), .Q(
        branchOffset_regD[1]) );
  DFFRX1 \branchOffset_regD_reg[0]  ( .D(n307), .CK(clk), .RN(n36), .Q(
        branchOffset_regD[0]) );
  DFFRX1 \PCplus4_regD_reg[7]  ( .D(n330), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[7]), .QN(n151) );
  DFFRX1 \PCplus4_regD_reg[6]  ( .D(n329), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[6]), .QN(n150) );
  DFFRX1 \PCplus4_regD_reg[5]  ( .D(n328), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[5]), .QN(n149) );
  DFFRX1 \PCplus4_regD_reg[4]  ( .D(n327), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[4]), .QN(n148) );
  DFFRX1 \PCplus4_regD_reg[9]  ( .D(n332), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[9]), .QN(n153) );
  DFFRX1 \PCplus4_regD_reg[8]  ( .D(n331), .CK(clk), .RN(n28), .Q(
        PCplus4_regD[8]), .QN(n152) );
  DFFRX1 \PCplus4_regD_reg[16]  ( .D(n339), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[16]), .QN(n160) );
  DFFRX1 \PCplus4_regD_reg[11]  ( .D(n334), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[11]), .QN(n155) );
  DFFRX1 \PCplus4_regD_reg[27]  ( .D(n350), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[27]) );
  DFFRX1 \PCplus4_regD_reg[26]  ( .D(n349), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[26]), .QN(n170) );
  DFFRX1 \PCplus4_regD_reg[25]  ( .D(n348), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[25]) );
  DFFRX1 \PCplus4_regD_reg[24]  ( .D(n347), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[24]) );
  DFFRX1 \PCplus4_regD_reg[23]  ( .D(n346), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[23]) );
  DFFRX1 \PCplus4_regD_reg[22]  ( .D(n345), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[22]), .QN(n166) );
  DFFRX1 \PCplus4_regD_reg[21]  ( .D(n344), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[21]), .QN(n165) );
  DFFRX1 \PCplus4_regD_reg[20]  ( .D(n343), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[20]), .QN(n164) );
  DFFRX1 \PCplus4_regD_reg[19]  ( .D(n342), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[19]), .QN(n163) );
  DFFRX1 \PCplus4_regD_reg[18]  ( .D(n341), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[18]), .QN(n162) );
  DFFRX1 \PCplus4_regD_reg[17]  ( .D(n340), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[17]), .QN(n161) );
  DFFRX1 \PCplus4_regD_reg[15]  ( .D(n338), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[15]), .QN(n159) );
  DFFRX1 \PCplus4_regD_reg[14]  ( .D(n337), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[14]), .QN(n158) );
  DFFRX1 \PCplus4_regD_reg[1]  ( .D(n324), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[1]), .QN(n145) );
  DFFRX1 \PCplus4_regD_reg[0]  ( .D(n323), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[0]), .QN(n144) );
  DFFRX1 \PCplus4_regD_reg[10]  ( .D(n333), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[10]), .QN(n154) );
  DFFRX1 \PCplus4_regD_reg[12]  ( .D(n335), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[12]), .QN(n156) );
  DFFRX1 \PCplus4_regD_reg[13]  ( .D(n336), .CK(clk), .RN(n25), .Q(
        PCplus4_regD[13]), .QN(n157) );
  DFFRX1 \PCplus4_regD_reg[3]  ( .D(n326), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[3]), .QN(n147) );
  DFFRX1 \PCplus4_regD_reg[2]  ( .D(n325), .CK(clk), .RN(n30), .Q(
        PCplus4_regD[2]), .QN(n146) );
  DFFRX1 \PCplus4_regD_reg[30]  ( .D(n353), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[30]), .QN(n174) );
  DFFRX1 \PCplus4_regD_reg[29]  ( .D(n352), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[29]), .QN(n173) );
  DFFRX1 \PCplus4_regD_reg[28]  ( .D(n351), .CK(clk), .RN(n26), .Q(
        PCplus4_regD[28]), .QN(n172) );
  DFFRX1 \B_regD_reg[19]  ( .D(n244), .CK(clk), .RN(n43), .Q(B_regD[19]), .QN(
        n65) );
  DFFRX1 \B_regD_reg[27]  ( .D(n252), .CK(clk), .RN(n44), .Q(B_regD[27]), .QN(
        n73) );
  DFFRX1 \B_regD_reg[29]  ( .D(n254), .CK(clk), .RN(n44), .Q(B_regD[29]), .QN(
        n75) );
  DFFRX1 \B_regD_reg[30]  ( .D(n255), .CK(clk), .RN(n44), .Q(B_regD[30]), .QN(
        n76) );
  DFFRX1 \B_regD_reg[23]  ( .D(n248), .CK(clk), .RN(n44), .Q(B_regD[23]), .QN(
        n69) );
  DFFRX1 \B_regD_reg[15]  ( .D(n240), .CK(clk), .RN(n43), .Q(B_regD[15]), .QN(
        n61) );
  DFFRX1 \B_regD_reg[12]  ( .D(n237), .CK(clk), .RN(n43), .Q(B_regD[12]), .QN(
        n58) );
  DFFRX1 \B_regD_reg[26]  ( .D(n251), .CK(clk), .RN(n44), .Q(B_regD[26]), .QN(
        n72) );
  DFFRX1 \B_regD_reg[22]  ( .D(n247), .CK(clk), .RN(n42), .Q(B_regD[22]), .QN(
        n68) );
  DFFRX1 \B_regD_reg[10]  ( .D(n235), .CK(clk), .RN(n45), .Q(B_regD[10]), .QN(
        n56) );
  DFFRX1 \B_regD_reg[14]  ( .D(n239), .CK(clk), .RN(n43), .Q(B_regD[14]), .QN(
        n60) );
  DFFRX1 \B_regD_reg[24]  ( .D(n249), .CK(clk), .RN(n44), .Q(B_regD[24]), .QN(
        n70) );
  DFFRX1 \B_regD_reg[6]  ( .D(n231), .CK(clk), .RN(n53), .Q(B_regD[6]), .QN(
        n52) );
  DFFRX1 \B_regD_reg[13]  ( .D(n238), .CK(clk), .RN(n43), .Q(B_regD[13]), .QN(
        n59) );
  DFFRX1 \B_regD_reg[18]  ( .D(n243), .CK(clk), .RN(n43), .Q(B_regD[18]), .QN(
        n64) );
  DFFRX1 \B_regD_reg[25]  ( .D(n250), .CK(clk), .RN(n44), .Q(B_regD[25]), .QN(
        n71) );
  DFFRX1 \B_regD_reg[17]  ( .D(n242), .CK(clk), .RN(n43), .Q(B_regD[17]), .QN(
        n63) );
  DFFRX1 \B_regD_reg[9]  ( .D(n234), .CK(clk), .RN(n53), .Q(B_regD[9]), .QN(
        n55) );
  DFFRX1 \B_regD_reg[21]  ( .D(n246), .CK(clk), .RN(n43), .Q(B_regD[21]), .QN(
        n67) );
  DFFRX1 \B_regD_reg[11]  ( .D(n236), .CK(clk), .RN(n43), .Q(B_regD[11]), .QN(
        n57) );
  DFFRX1 \A_regD_reg[23]  ( .D(n280), .CK(clk), .RN(n42), .Q(A_regD[23]), .QN(
        n101) );
  DFFRX1 \B_regD_reg[16]  ( .D(n241), .CK(clk), .RN(n43), .Q(B_regD[16]), .QN(
        n62) );
  DFFRX1 \A_regD_reg[19]  ( .D(n276), .CK(clk), .RN(n42), .Q(A_regD[19]), .QN(
        n97) );
  DFFRX1 \B_regD_reg[8]  ( .D(n233), .CK(clk), .RN(n53), .Q(B_regD[8]), .QN(
        n54) );
  DFFRX1 \A_regD_reg[24]  ( .D(n281), .CK(clk), .RN(n42), .Q(A_regD[24]), .QN(
        n102) );
  DFFRX1 \A_regD_reg[22]  ( .D(n279), .CK(clk), .RN(n42), .Q(A_regD[22]), .QN(
        n100) );
  DFFRX1 \A_regD_reg[20]  ( .D(n277), .CK(clk), .RN(n42), .Q(A_regD[20]), .QN(
        n98) );
  DFFRX1 \A_regD_reg[15]  ( .D(n272), .CK(clk), .RN(n42), .Q(A_regD[15]), .QN(
        n93) );
  DFFRX1 \A_regD_reg[18]  ( .D(n275), .CK(clk), .RN(n42), .Q(A_regD[18]), .QN(
        n96) );
  DFFRX1 \A_regD_reg[0]  ( .D(n257), .CK(clk), .RN(n44), .Q(A_regD[0]), .QN(
        n78) );
  DFFRX1 \A_regD_reg[21]  ( .D(n278), .CK(clk), .RN(n42), .Q(A_regD[21]), .QN(
        n99) );
  DFFRX1 \A_regD_reg[17]  ( .D(n274), .CK(clk), .RN(n42), .Q(A_regD[17]), .QN(
        n95) );
  DFFRX1 \A_regD_reg[16]  ( .D(n273), .CK(clk), .RN(n42), .Q(A_regD[16]), .QN(
        n94) );
  DFFRX1 \B_regD_reg[2]  ( .D(n227), .CK(clk), .RN(n53), .Q(B_regD[2]), .QN(
        n48) );
  DFFRX1 \B_regD_reg[1]  ( .D(n226), .CK(clk), .RN(n53), .Q(B_regD[1]), .QN(
        n47) );
  DFFRX1 \ExtOut_regD_reg[0]  ( .D(n193), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[0]), .QN(n14) );
  DFFRX1 \ExtOut_regD_reg[24]  ( .D(n217), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[24]), .QN(n38) );
  DFFRX1 \ExtOut_regD_reg[13]  ( .D(n206), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[13]), .QN(n27) );
  DFFRX1 \ExtOut_regD_reg[25]  ( .D(n218), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[25]), .QN(n39) );
  DFFRX1 \ExtOut_regD_reg[15]  ( .D(n208), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[15]), .QN(n29) );
  DFFRX1 \ExtOut_regD_reg[17]  ( .D(n210), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[17]), .QN(n31) );
  DFFRX1 \ExtOut_regD_reg[9]  ( .D(n202), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[9]), .QN(n23) );
  DFFRX1 \ExtOut_regD_reg[20]  ( .D(n213), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[20]), .QN(n34) );
  DFFRX1 \ExtOut_regD_reg[21]  ( .D(n214), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[21]), .QN(n35) );
  DFFRX1 \A_regD_reg[25]  ( .D(n282), .CK(clk), .RN(n42), .Q(A_regD[25]), .QN(
        n103) );
  DFFRX1 \B_regD_reg[5]  ( .D(n230), .CK(clk), .RN(n53), .Q(B_regD[5]), .QN(
        n51) );
  DFFRX1 \B_regD_reg[4]  ( .D(n229), .CK(clk), .RN(n53), .Q(B_regD[4]), .QN(
        n50) );
  DFFRX1 \B_regD_reg[3]  ( .D(n228), .CK(clk), .RN(n53), .Q(B_regD[3]), .QN(
        n49) );
  DFFRX1 \ExtOut_regD_reg[18]  ( .D(n211), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[18]), .QN(n32) );
  DFFRX1 \ExtOut_regD_reg[23]  ( .D(n216), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[23]), .QN(n37) );
  DFFRX2 \B_regD_reg[31]  ( .D(n256), .CK(clk), .RN(n44), .Q(B_regD[31]), .QN(
        n77) );
  DFFRX2 \B_regD_reg[28]  ( .D(n253), .CK(clk), .RN(n44), .Q(B_regD[28]), .QN(
        n74) );
  DFFRX2 \A_regD_reg[30]  ( .D(n287), .CK(clk), .RN(n36), .Q(A_regD[30]), .QN(
        n108) );
  DFFRX2 \A_regD_reg[26]  ( .D(n283), .CK(clk), .RN(n41), .Q(A_regD[26]), .QN(
        n104) );
  DFFRHQX8 \Rs_regD_reg[4]  ( .D(n192), .CK(clk), .RN(n66), .Q(Rs_regD[4]) );
  DFFRX2 \ExtOut_regD_reg[19]  ( .D(n212), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[19]), .QN(n33) );
  DFFRHQX8 \Rt_regD_reg[0]  ( .D(n183), .CK(clk), .RN(n80), .Q(Rt_regD[0]) );
  DFFRHQX8 \Rt_regD_reg[3]  ( .D(n186), .CK(clk), .RN(n80), .Q(Rt_regD[3]) );
  DFFRHQX8 \Rt_regD_reg[1]  ( .D(n184), .CK(clk), .RN(n80), .Q(Rt_regD[1]) );
  DFFRHQX8 \Rt_regD_reg[4]  ( .D(n187), .CK(clk), .RN(n79), .Q(Rt_regD[4]) );
  DFFRHQX8 \Rs_regD_reg[2]  ( .D(n190), .CK(clk), .RN(n66), .Q(Rs_regD[2]) );
  DFFRHQX8 \Rt_regD_reg[2]  ( .D(n185), .CK(clk), .RN(n80), .Q(Rt_regD[2]) );
  DFFRHQX8 \Rs_regD_reg[1]  ( .D(n189), .CK(clk), .RN(n66), .Q(Rs_regD[1]) );
  DFFRHQX8 \Rs_regD_reg[3]  ( .D(n191), .CK(clk), .RN(rst_n), .Q(Rs_regD[3])
         );
  DFFRX4 \B_regD_reg[0]  ( .D(n225), .CK(clk), .RN(n53), .Q(B_regD[0]), .QN(
        n46) );
  DFFRHQX8 \Rs_regD_reg[0]  ( .D(n188), .CK(clk), .RN(n66), .Q(Rs_regD[0]) );
  DFFRX1 \ExtOut_regD_reg[22]  ( .D(n215), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[22]) );
  DFFRX1 \ExtOut_regD_reg[16]  ( .D(n209), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[16]) );
  DFFRX1 \ExtOut_regD_reg[14]  ( .D(n207), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[14]) );
  DFFRX1 \A_regD_reg[1]  ( .D(n258), .CK(clk), .RN(n44), .Q(A_regD[1]) );
  DFFRX1 \ExtOut_regD_reg[26]  ( .D(n219), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[26]) );
  DFFRX1 \A_regD_reg[31]  ( .D(n288), .CK(clk), .RN(n36), .Q(A_regD[31]) );
  DFFRX1 \A_regD_reg[29]  ( .D(n286), .CK(clk), .RN(n36), .Q(A_regD[29]) );
  DFFRX1 \A_regD_reg[28]  ( .D(n285), .CK(clk), .RN(n36), .Q(A_regD[28]) );
  DFFRX1 \A_regD_reg[27]  ( .D(n284), .CK(clk), .RN(n36), .Q(A_regD[27]) );
  DFFRX1 \ExtOut_regD_reg[12]  ( .D(n205), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[12]) );
  DFFRX1 \ExtOut_regD_reg[11]  ( .D(n204), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[11]) );
  DFFRX1 \ExtOut_regD_reg[10]  ( .D(n203), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[10]) );
  DFFRX1 \ExtOut_regD_reg[8]  ( .D(n201), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[8]) );
  DFFRX1 \ExtOut_regD_reg[7]  ( .D(n200), .CK(clk), .RN(n79), .Q(
        ExtOut_regD[7]) );
  DFFRX1 \ExtOut_regD_reg[6]  ( .D(n199), .CK(clk), .RN(n53), .Q(
        ExtOut_regD[6]) );
  DFFRX1 \ExtOut_regD_reg[3]  ( .D(n196), .CK(clk), .RN(n66), .Q(
        ExtOut_regD[3]) );
  DFFRX1 \B_regD_reg[20]  ( .D(n245), .CK(clk), .RN(n43), .Q(B_regD[20]) );
  DFFRX1 \B_regD_reg[7]  ( .D(n232), .CK(clk), .RN(n53), .Q(B_regD[7]) );
  DFFRX1 \A_regD_reg[14]  ( .D(n271), .CK(clk), .RN(n40), .Q(A_regD[14]) );
  DFFRX1 \A_regD_reg[13]  ( .D(n270), .CK(clk), .RN(n41), .Q(A_regD[13]) );
  DFFRX1 \A_regD_reg[12]  ( .D(n269), .CK(clk), .RN(n41), .Q(A_regD[12]) );
  DFFRX1 \A_regD_reg[11]  ( .D(n268), .CK(clk), .RN(n41), .Q(A_regD[11]) );
  DFFRX1 \A_regD_reg[10]  ( .D(n267), .CK(clk), .RN(n41), .Q(A_regD[10]) );
  DFFRX1 \A_regD_reg[8]  ( .D(n265), .CK(clk), .RN(n41), .Q(A_regD[8]) );
  DFFRX1 \A_regD_reg[2]  ( .D(n259), .CK(clk), .RN(n43), .Q(A_regD[2]) );
  DFFRX1 \MemtoReg_regD_reg[0]  ( .D(n299), .CK(clk), .RN(n40), .Q(
        MemtoReg_regD[0]) );
  DFFRX1 \MemtoReg_regD_reg[1]  ( .D(n300), .CK(clk), .RN(n40), .Q(
        MemtoReg_regD[1]) );
  DFFRX1 \ExtOut_regD_reg[31]  ( .D(n224), .CK(clk), .RN(n53), .Q(
        ExtOut_regD[31]) );
  DFFRX1 \ExtOut_regD_reg[30]  ( .D(n223), .CK(clk), .RN(n44), .Q(
        ExtOut_regD[30]) );
  DFFRX1 \ExtOut_regD_reg[28]  ( .D(n221), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[28]) );
  DFFRX1 \ExtOut_regD_reg[27]  ( .D(n220), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[27]) );
  DFFSRHQX4 \ALUOp_regD_reg[0]  ( .D(n293), .CK(clk), .SN(1'b1), .RN(n36), .Q(
        ALUOp_regD[0]) );
  DFFSRHQX4 \funct_regD_reg[5]  ( .D(n306), .CK(clk), .SN(1'b1), .RN(n40), .Q(
        funct_regD[5]) );
  DFFSRHQX4 ALUsrc_regD_reg ( .D(n289), .CK(clk), .SN(1'b1), .RN(n36), .Q(
        ALUsrc_regD) );
  DFFRX4 \ExtOut_regD_reg[29]  ( .D(n222), .CK(clk), .RN(n45), .Q(
        ExtOut_regD[29]) );
  DFFRX2 RegWrite_regD_reg ( .D(n290), .CK(clk), .RN(n36), .Q(RegWrite_regD)
         );
  BUFX20 U2 ( .A(n112), .Y(n106) );
  CLKBUFX2 U3 ( .A(n127), .Y(n114) );
  BUFX16 U4 ( .A(n120), .Y(n92) );
  BUFX4 U5 ( .A(n128), .Y(n110) );
  BUFX4 U6 ( .A(stallcache), .Y(n127) );
  CLKBUFX2 U7 ( .A(rst_n), .Y(n89) );
  CLKBUFX2 U8 ( .A(rst_n), .Y(n86) );
  CLKBUFX2 U9 ( .A(rst_n), .Y(n90) );
  BUFX4 U10 ( .A(n121), .Y(n120) );
  CLKBUFX2 U11 ( .A(rst_n), .Y(n88) );
  BUFX6 U12 ( .A(n120), .Y(n91) );
  CLKMX2X4 U13 ( .A(branchOffset_D[8]), .B(branchOffset_regD[8]), .S0(n91), 
        .Y(n315) );
  CLKMX2X3 U14 ( .A(MemWrite), .B(MemWrite_regD), .S0(n92), .Y(n291) );
  CLKMX2X2 U18 ( .A(Rs[4]), .B(Rs_regD[4]), .S0(n92), .Y(n192) );
  INVXL U19 ( .A(Rt_regD[2]), .Y(n10) );
  INVXL U20 ( .A(Rt_regD[4]), .Y(n13) );
  INVXL U21 ( .A(Rt_regD[3]), .Y(n21) );
  CLKBUFX3 U22 ( .A(n112), .Y(n107) );
  CLKBUFX3 U23 ( .A(stallcache), .Y(n128) );
  CLKBUFX2 U24 ( .A(stallcache), .Y(n121) );
  CLKMX2X2 U25 ( .A(funct[5]), .B(funct_regD[5]), .S0(n106), .Y(n306) );
  MX2XL U26 ( .A(ExtOut[27]), .B(ExtOut_regD[27]), .S0(n107), .Y(n220) );
  MX2XL U27 ( .A(ExtOut[28]), .B(ExtOut_regD[28]), .S0(n107), .Y(n221) );
  MX2XL U28 ( .A(ExtOut[29]), .B(ExtOut_regD[29]), .S0(n107), .Y(n222) );
  MX2XL U29 ( .A(ExtOut[30]), .B(ExtOut_regD[30]), .S0(n107), .Y(n223) );
  MX2XL U30 ( .A(ExtOut[31]), .B(ExtOut_regD[31]), .S0(n107), .Y(n224) );
  MX2XL U31 ( .A(ExtOut[15]), .B(n384), .S0(n106), .Y(n208) );
  MX2XL U32 ( .A(ExtOut[16]), .B(ExtOut_regD[16]), .S0(n106), .Y(n209) );
  MX2XL U33 ( .A(ExtOut[17]), .B(n385), .S0(n106), .Y(n210) );
  MX2XL U34 ( .A(ExtOut[19]), .B(n387), .S0(n106), .Y(n212) );
  MX2XL U35 ( .A(ExtOut[20]), .B(n388), .S0(n106), .Y(n213) );
  MX2XL U36 ( .A(ExtOut[21]), .B(n389), .S0(n106), .Y(n214) );
  MX2XL U37 ( .A(ExtOut[22]), .B(ExtOut_regD[22]), .S0(n106), .Y(n215) );
  MX2XL U38 ( .A(ExtOut[23]), .B(n390), .S0(n106), .Y(n216) );
  MX2XL U39 ( .A(ExtOut[24]), .B(n391), .S0(n106), .Y(n217) );
  MX2XL U40 ( .A(ExtOut[25]), .B(n392), .S0(n106), .Y(n218) );
  MX2XL U41 ( .A(ExtOut[14]), .B(ExtOut_regD[14]), .S0(n106), .Y(n207) );
  CLKMX2X2 U42 ( .A(ExtOut[3]), .B(ExtOut_regD[3]), .S0(n105), .Y(n196) );
  CLKMX2X2 U43 ( .A(ExtOut[6]), .B(ExtOut_regD[6]), .S0(n105), .Y(n199) );
  CLKMX2X2 U44 ( .A(ExtOut[7]), .B(ExtOut_regD[7]), .S0(n105), .Y(n200) );
  CLKMX2X2 U45 ( .A(ExtOut[8]), .B(ExtOut_regD[8]), .S0(n105), .Y(n201) );
  CLKMX2X2 U46 ( .A(ExtOut[9]), .B(n382), .S0(n105), .Y(n202) );
  CLKMX2X2 U47 ( .A(ExtOut[10]), .B(ExtOut_regD[10]), .S0(n105), .Y(n203) );
  CLKMX2X2 U48 ( .A(ExtOut[11]), .B(ExtOut_regD[11]), .S0(n105), .Y(n204) );
  CLKMX2X2 U49 ( .A(ExtOut[12]), .B(ExtOut_regD[12]), .S0(n105), .Y(n205) );
  MX2XL U50 ( .A(branchOffset_D[0]), .B(branchOffset_regD[0]), .S0(n91), .Y(
        n307) );
  MX2XL U51 ( .A(branchOffset_D[13]), .B(n130), .S0(n106), .Y(n320) );
  MX2XL U52 ( .A(PCplus4_regI[10]), .B(n171), .S0(n92), .Y(n333) );
  CLKBUFX3 U53 ( .A(n121), .Y(n109) );
  CLKBUFX3 U54 ( .A(n128), .Y(n111) );
  CLKBUFX3 U55 ( .A(n114), .Y(n105) );
  CLKBUFX3 U56 ( .A(n90), .Y(n79) );
  CLKBUFX3 U57 ( .A(n90), .Y(n53) );
  CLKBUFX3 U58 ( .A(n89), .Y(n45) );
  CLKBUFX3 U59 ( .A(n90), .Y(n44) );
  CLKBUFX3 U60 ( .A(n89), .Y(n43) );
  CLKBUFX3 U61 ( .A(n89), .Y(n42) );
  CLKBUFX3 U62 ( .A(n88), .Y(n41) );
  CLKBUFX3 U63 ( .A(n86), .Y(n40) );
  CLKBUFX3 U64 ( .A(n88), .Y(n36) );
  CLKBUFX3 U65 ( .A(n88), .Y(n30) );
  CLKBUFX3 U66 ( .A(n86), .Y(n28) );
  CLKBUFX3 U67 ( .A(n86), .Y(n26) );
  CLKBUFX3 U68 ( .A(n89), .Y(n80) );
  CLKBUFX3 U69 ( .A(n90), .Y(n66) );
  CLKBUFX3 U70 ( .A(n127), .Y(n112) );
  CLKBUFX3 U71 ( .A(n86), .Y(n25) );
  CLKMX2X2 U72 ( .A(MemRead), .B(n448), .S0(n92), .Y(n292) );
  INVX1 U73 ( .A(n113), .Y(n448) );
  CLKMX2X2 U74 ( .A(Branch), .B(n372), .S0(n92), .Y(n176) );
  INVX1 U75 ( .A(n2), .Y(n372) );
  CLKMX2X2 U76 ( .A(JumpReg), .B(n373), .S0(n106), .Y(n177) );
  INVX1 U77 ( .A(n3), .Y(n373) );
  CLKMX2X2 U78 ( .A(RegWrite), .B(RegWrite_regD), .S0(n110), .Y(n290) );
  CLKMX2X2 U79 ( .A(funct[0]), .B(n443), .S0(n106), .Y(n301) );
  CLKINVX1 U80 ( .A(n122), .Y(n443) );
  CLKMX2X2 U81 ( .A(funct[1]), .B(n444), .S0(n110), .Y(n302) );
  CLKINVX1 U82 ( .A(n123), .Y(n444) );
  CLKMX2X2 U83 ( .A(funct[2]), .B(n445), .S0(n106), .Y(n303) );
  CLKINVX1 U84 ( .A(n124), .Y(n445) );
  CLKMX2X2 U85 ( .A(funct[3]), .B(n446), .S0(n106), .Y(n304) );
  CLKINVX1 U86 ( .A(n125), .Y(n446) );
  CLKMX2X2 U87 ( .A(funct[4]), .B(n447), .S0(n106), .Y(n305) );
  CLKINVX1 U88 ( .A(n126), .Y(n447) );
  MX2XL U89 ( .A(MemtoReg[1]), .B(MemtoReg_regD[1]), .S0(n120), .Y(n300) );
  CLKMX2X2 U90 ( .A(ALUOp[0]), .B(ALUOp_regD[0]), .S0(n92), .Y(n293) );
  CLKMX2X2 U91 ( .A(ALUOp[1]), .B(n449), .S0(n92), .Y(n294) );
  CLKINVX1 U92 ( .A(n115), .Y(n449) );
  CLKMX2X2 U93 ( .A(ALUOp[2]), .B(n450), .S0(n92), .Y(n295) );
  CLKINVX1 U94 ( .A(n116), .Y(n450) );
  CLKMX2X2 U95 ( .A(ALUOp[3]), .B(n451), .S0(n92), .Y(n296) );
  CLKINVX1 U96 ( .A(n117), .Y(n451) );
  CLKMX2X2 U97 ( .A(ALUOp[4]), .B(n452), .S0(n92), .Y(n297) );
  CLKINVX1 U98 ( .A(n118), .Y(n452) );
  CLKMX2X2 U99 ( .A(ALUOp[5]), .B(n453), .S0(n92), .Y(n298) );
  CLKINVX1 U100 ( .A(n119), .Y(n453) );
  MX2XL U101 ( .A(MemtoReg[0]), .B(MemtoReg_regD[0]), .S0(n106), .Y(n299) );
  MX2XL U102 ( .A(Rs[2]), .B(Rs_regD[2]), .S0(n106), .Y(n190) );
  MX2XL U103 ( .A(Rs[0]), .B(Rs_regD[0]), .S0(n120), .Y(n188) );
  MX2XL U104 ( .A(Rs[1]), .B(Rs_regD[1]), .S0(n106), .Y(n189) );
  MX2XL U105 ( .A(Rs[3]), .B(Rs_regD[3]), .S0(n110), .Y(n191) );
  MX2XL U106 ( .A(wsel[0]), .B(wsel_regD[0]), .S0(n106), .Y(n178) );
  MX2XL U107 ( .A(wsel[1]), .B(wsel_regD[1]), .S0(n92), .Y(n179) );
  MX2XL U108 ( .A(wsel[2]), .B(wsel_regD[2]), .S0(n120), .Y(n180) );
  MX2XL U109 ( .A(wsel[3]), .B(wsel_regD[3]), .S0(n120), .Y(n181) );
  MX2XL U110 ( .A(wsel[4]), .B(wsel_regD[4]), .S0(n106), .Y(n182) );
  CLKMX2X2 U111 ( .A(Rt[0]), .B(Rt_regD[0]), .S0(n92), .Y(n183) );
  CLKMX2X2 U112 ( .A(Rt[1]), .B(Rt_regD[1]), .S0(n106), .Y(n184) );
  CLKMX2X2 U113 ( .A(Rt[2]), .B(n374), .S0(n92), .Y(n185) );
  CLKINVX1 U114 ( .A(n10), .Y(n374) );
  CLKMX2X2 U115 ( .A(Rt[3]), .B(n375), .S0(n106), .Y(n186) );
  CLKINVX1 U116 ( .A(n21), .Y(n375) );
  CLKMX2X2 U117 ( .A(Rt[4]), .B(n376), .S0(n92), .Y(n187) );
  CLKINVX1 U118 ( .A(n13), .Y(n376) );
  CLKMX2X2 U119 ( .A(ExtOut[0]), .B(n377), .S0(n105), .Y(n193) );
  CLKINVX1 U120 ( .A(n14), .Y(n377) );
  CLKMX2X2 U121 ( .A(ExtOut[1]), .B(n378), .S0(n105), .Y(n194) );
  CLKINVX1 U122 ( .A(n15), .Y(n378) );
  CLKMX2X2 U123 ( .A(ExtOut[2]), .B(n379), .S0(n105), .Y(n195) );
  CLKINVX1 U124 ( .A(n16), .Y(n379) );
  CLKMX2X2 U125 ( .A(ExtOut[4]), .B(n380), .S0(n105), .Y(n197) );
  CLKINVX1 U126 ( .A(n18), .Y(n380) );
  CLKMX2X2 U127 ( .A(ExtOut[5]), .B(n381), .S0(n105), .Y(n198) );
  CLKINVX1 U128 ( .A(n19), .Y(n381) );
  CLKINVX1 U129 ( .A(n23), .Y(n382) );
  CLKMX2X2 U130 ( .A(ExtOut[13]), .B(n383), .S0(n106), .Y(n206) );
  CLKINVX1 U131 ( .A(n27), .Y(n383) );
  CLKINVX1 U132 ( .A(n29), .Y(n384) );
  CLKINVX1 U133 ( .A(n31), .Y(n385) );
  MX2XL U134 ( .A(ExtOut[18]), .B(n386), .S0(n106), .Y(n211) );
  CLKINVX1 U135 ( .A(n32), .Y(n386) );
  CLKINVX1 U136 ( .A(n33), .Y(n387) );
  CLKINVX1 U137 ( .A(n34), .Y(n388) );
  CLKINVX1 U138 ( .A(n35), .Y(n389) );
  CLKINVX1 U139 ( .A(n37), .Y(n390) );
  CLKINVX1 U140 ( .A(n38), .Y(n391) );
  CLKINVX1 U141 ( .A(n39), .Y(n392) );
  CLKMX2X2 U142 ( .A(ExtOut[26]), .B(ExtOut_regD[26]), .S0(n107), .Y(n219) );
  MX2XL U143 ( .A(B[0]), .B(n393), .S0(n107), .Y(n225) );
  CLKINVX1 U144 ( .A(n46), .Y(n393) );
  MX2XL U145 ( .A(B[1]), .B(n394), .S0(n107), .Y(n226) );
  CLKINVX1 U146 ( .A(n47), .Y(n394) );
  MX2XL U147 ( .A(B[2]), .B(n395), .S0(n107), .Y(n227) );
  CLKINVX1 U148 ( .A(n48), .Y(n395) );
  MX2XL U149 ( .A(B[3]), .B(n396), .S0(n107), .Y(n228) );
  CLKINVX1 U150 ( .A(n49), .Y(n396) );
  MX2XL U151 ( .A(B[4]), .B(n397), .S0(n107), .Y(n229) );
  CLKINVX1 U152 ( .A(n50), .Y(n397) );
  MX2XL U153 ( .A(B[5]), .B(n398), .S0(n107), .Y(n230) );
  CLKINVX1 U154 ( .A(n51), .Y(n398) );
  MX2XL U155 ( .A(B[6]), .B(n399), .S0(n107), .Y(n231) );
  CLKINVX1 U156 ( .A(n52), .Y(n399) );
  CLKMX2X2 U157 ( .A(B[7]), .B(B_regD[7]), .S0(n92), .Y(n232) );
  MX2XL U158 ( .A(B[8]), .B(n400), .S0(n106), .Y(n233) );
  CLKINVX1 U159 ( .A(n54), .Y(n400) );
  MX2XL U160 ( .A(B[9]), .B(n401), .S0(n106), .Y(n234) );
  CLKINVX1 U161 ( .A(n55), .Y(n401) );
  MX2XL U162 ( .A(B[10]), .B(n402), .S0(n106), .Y(n235) );
  CLKINVX1 U163 ( .A(n56), .Y(n402) );
  MX2XL U164 ( .A(B[11]), .B(n403), .S0(n106), .Y(n236) );
  CLKINVX1 U165 ( .A(n57), .Y(n403) );
  MX2XL U166 ( .A(B[12]), .B(n404), .S0(n106), .Y(n237) );
  CLKINVX1 U167 ( .A(n58), .Y(n404) );
  MX2XL U168 ( .A(B[13]), .B(n405), .S0(n106), .Y(n238) );
  CLKINVX1 U169 ( .A(n59), .Y(n405) );
  MX2XL U170 ( .A(B[14]), .B(n406), .S0(n106), .Y(n239) );
  CLKINVX1 U171 ( .A(n60), .Y(n406) );
  MX2XL U172 ( .A(B[15]), .B(n407), .S0(n106), .Y(n240) );
  CLKINVX1 U173 ( .A(n61), .Y(n407) );
  MX2XL U174 ( .A(B[16]), .B(n408), .S0(n106), .Y(n241) );
  CLKINVX1 U175 ( .A(n62), .Y(n408) );
  MX2XL U176 ( .A(B[17]), .B(n409), .S0(n106), .Y(n242) );
  CLKINVX1 U177 ( .A(n63), .Y(n409) );
  MX2XL U178 ( .A(B[18]), .B(n410), .S0(n106), .Y(n243) );
  CLKINVX1 U179 ( .A(n64), .Y(n410) );
  MX2XL U180 ( .A(B[19]), .B(n411), .S0(n106), .Y(n244) );
  CLKINVX1 U181 ( .A(n65), .Y(n411) );
  CLKMX2X2 U182 ( .A(B[20]), .B(B_regD[20]), .S0(n109), .Y(n245) );
  MX2XL U183 ( .A(B[21]), .B(n412), .S0(n109), .Y(n246) );
  CLKINVX1 U184 ( .A(n67), .Y(n412) );
  MX2XL U185 ( .A(B[22]), .B(n413), .S0(n109), .Y(n247) );
  CLKINVX1 U186 ( .A(n68), .Y(n413) );
  MX2XL U187 ( .A(B[23]), .B(n414), .S0(n109), .Y(n248) );
  CLKINVX1 U188 ( .A(n69), .Y(n414) );
  MX2XL U189 ( .A(B[24]), .B(n415), .S0(n109), .Y(n249) );
  CLKINVX1 U190 ( .A(n70), .Y(n415) );
  MX2XL U191 ( .A(B[25]), .B(n416), .S0(n109), .Y(n250) );
  CLKINVX1 U192 ( .A(n71), .Y(n416) );
  MX2XL U193 ( .A(B[26]), .B(n417), .S0(n109), .Y(n251) );
  CLKINVX1 U194 ( .A(n72), .Y(n417) );
  MX2XL U195 ( .A(B[27]), .B(n418), .S0(n109), .Y(n252) );
  CLKINVX1 U196 ( .A(n73), .Y(n418) );
  MX2XL U197 ( .A(B[28]), .B(n419), .S0(n109), .Y(n253) );
  CLKINVX1 U198 ( .A(n74), .Y(n419) );
  MX2XL U199 ( .A(B[29]), .B(n420), .S0(n109), .Y(n254) );
  CLKINVX1 U200 ( .A(n75), .Y(n420) );
  MX2XL U201 ( .A(B[30]), .B(n421), .S0(n109), .Y(n255) );
  CLKINVX1 U202 ( .A(n76), .Y(n421) );
  MX2XL U203 ( .A(B[31]), .B(n422), .S0(n109), .Y(n256) );
  CLKINVX1 U204 ( .A(n77), .Y(n422) );
  MX2XL U205 ( .A(A[0]), .B(n423), .S0(n109), .Y(n257) );
  CLKINVX1 U206 ( .A(n78), .Y(n423) );
  CLKMX2X2 U207 ( .A(A[1]), .B(A_regD[1]), .S0(n110), .Y(n258) );
  MX2XL U208 ( .A(A[2]), .B(A_regD[2]), .S0(n110), .Y(n259) );
  CLKMX2X2 U209 ( .A(A[3]), .B(n424), .S0(n110), .Y(n260) );
  CLKINVX1 U210 ( .A(n81), .Y(n424) );
  CLKMX2X2 U211 ( .A(A[4]), .B(n425), .S0(n110), .Y(n261) );
  CLKINVX1 U212 ( .A(n82), .Y(n425) );
  CLKMX2X2 U213 ( .A(A[5]), .B(n426), .S0(n110), .Y(n262) );
  CLKINVX1 U214 ( .A(n83), .Y(n426) );
  CLKMX2X2 U215 ( .A(A[6]), .B(n427), .S0(n110), .Y(n263) );
  CLKINVX1 U216 ( .A(n84), .Y(n427) );
  CLKMX2X2 U217 ( .A(A[7]), .B(n428), .S0(n110), .Y(n264) );
  CLKINVX1 U218 ( .A(n85), .Y(n428) );
  MX2XL U219 ( .A(A[8]), .B(A_regD[8]), .S0(n110), .Y(n265) );
  CLKMX2X2 U220 ( .A(A[9]), .B(n429), .S0(n110), .Y(n266) );
  CLKINVX1 U221 ( .A(n87), .Y(n429) );
  MX2XL U222 ( .A(A[10]), .B(A_regD[10]), .S0(n110), .Y(n267) );
  MX2XL U223 ( .A(A[11]), .B(A_regD[11]), .S0(n110), .Y(n268) );
  MX2XL U224 ( .A(A[12]), .B(A_regD[12]), .S0(n110), .Y(n269) );
  MX2XL U225 ( .A(A[13]), .B(A_regD[13]), .S0(n110), .Y(n270) );
  CLKMX2X2 U226 ( .A(A[14]), .B(A_regD[14]), .S0(n111), .Y(n271) );
  MX2XL U227 ( .A(A[15]), .B(n430), .S0(n111), .Y(n272) );
  CLKINVX1 U228 ( .A(n93), .Y(n430) );
  MX2XL U229 ( .A(A[16]), .B(n431), .S0(n111), .Y(n273) );
  CLKINVX1 U230 ( .A(n94), .Y(n431) );
  MX2XL U231 ( .A(A[17]), .B(n432), .S0(n111), .Y(n274) );
  CLKINVX1 U232 ( .A(n95), .Y(n432) );
  MX2XL U233 ( .A(A[18]), .B(n433), .S0(n111), .Y(n275) );
  CLKINVX1 U234 ( .A(n96), .Y(n433) );
  MX2XL U235 ( .A(A[19]), .B(n434), .S0(n111), .Y(n276) );
  CLKINVX1 U236 ( .A(n97), .Y(n434) );
  MX2XL U237 ( .A(A[20]), .B(n435), .S0(n111), .Y(n277) );
  CLKINVX1 U238 ( .A(n98), .Y(n435) );
  MX2XL U239 ( .A(A[21]), .B(n436), .S0(n111), .Y(n278) );
  CLKINVX1 U240 ( .A(n99), .Y(n436) );
  MX2XL U241 ( .A(A[22]), .B(n437), .S0(n111), .Y(n279) );
  CLKINVX1 U242 ( .A(n100), .Y(n437) );
  MX2XL U243 ( .A(A[23]), .B(n438), .S0(n111), .Y(n280) );
  CLKINVX1 U244 ( .A(n101), .Y(n438) );
  MX2XL U245 ( .A(A[24]), .B(n439), .S0(n111), .Y(n281) );
  CLKINVX1 U246 ( .A(n102), .Y(n439) );
  MX2XL U247 ( .A(A[25]), .B(n440), .S0(n111), .Y(n282) );
  CLKINVX1 U248 ( .A(n103), .Y(n440) );
  MX2XL U249 ( .A(A[26]), .B(n441), .S0(n111), .Y(n283) );
  CLKINVX1 U250 ( .A(n104), .Y(n441) );
  MX2XL U251 ( .A(branchOffset_D[1]), .B(branchOffset_regD[1]), .S0(n91), .Y(
        n308) );
  MX2XL U252 ( .A(branchOffset_D[2]), .B(branchOffset_regD[2]), .S0(n91), .Y(
        n309) );
  MX2XL U253 ( .A(branchOffset_D[3]), .B(branchOffset_regD[3]), .S0(n91), .Y(
        n310) );
  MX2XL U254 ( .A(branchOffset_D[4]), .B(n129), .S0(n91), .Y(n311) );
  CLKINVX1 U255 ( .A(n132), .Y(n129) );
  MX2XL U256 ( .A(branchOffset_D[5]), .B(branchOffset_regD[5]), .S0(n91), .Y(
        n312) );
  MX2XL U257 ( .A(branchOffset_D[6]), .B(branchOffset_regD[6]), .S0(n91), .Y(
        n313) );
  MX2XL U258 ( .A(branchOffset_D[7]), .B(branchOffset_regD[7]), .S0(n91), .Y(
        n314) );
  MX2XL U259 ( .A(branchOffset_D[9]), .B(branchOffset_regD[9]), .S0(n91), .Y(
        n316) );
  MX2XL U260 ( .A(branchOffset_D[10]), .B(branchOffset_regD[10]), .S0(n91), 
        .Y(n317) );
  MX2XL U261 ( .A(branchOffset_D[11]), .B(branchOffset_regD[11]), .S0(n91), 
        .Y(n318) );
  MX2XL U262 ( .A(branchOffset_D[12]), .B(branchOffset_regD[12]), .S0(n91), 
        .Y(n319) );
  CLKINVX1 U263 ( .A(n141), .Y(n130) );
  MX2XL U264 ( .A(branchOffset_D[14]), .B(n131), .S0(n92), .Y(n321) );
  CLKINVX1 U265 ( .A(n142), .Y(n131) );
  MX2XL U266 ( .A(branchOffset_D[15]), .B(n133), .S0(n92), .Y(n322) );
  CLKINVX1 U267 ( .A(n143), .Y(n133) );
  MX2XL U268 ( .A(PCplus4_regI[0]), .B(n134), .S0(n92), .Y(n323) );
  CLKINVX1 U269 ( .A(n144), .Y(n134) );
  MX2XL U270 ( .A(PCplus4_regI[1]), .B(n135), .S0(n92), .Y(n324) );
  CLKINVX1 U271 ( .A(n145), .Y(n135) );
  MX2XL U272 ( .A(PCplus4_regI[2]), .B(n136), .S0(n106), .Y(n325) );
  CLKINVX1 U273 ( .A(n146), .Y(n136) );
  MX2XL U274 ( .A(PCplus4_regI[3]), .B(n137), .S0(n92), .Y(n326) );
  CLKINVX1 U275 ( .A(n147), .Y(n137) );
  MX2XL U276 ( .A(PCplus4_regI[4]), .B(n138), .S0(n92), .Y(n327) );
  CLKINVX1 U277 ( .A(n148), .Y(n138) );
  MX2XL U278 ( .A(PCplus4_regI[5]), .B(n139), .S0(n106), .Y(n328) );
  CLKINVX1 U279 ( .A(n149), .Y(n139) );
  MX2XL U280 ( .A(PCplus4_regI[6]), .B(n140), .S0(n92), .Y(n329) );
  CLKINVX1 U281 ( .A(n150), .Y(n140) );
  MX2XL U282 ( .A(PCplus4_regI[7]), .B(n167), .S0(n92), .Y(n330) );
  CLKINVX1 U283 ( .A(n151), .Y(n167) );
  MX2XL U284 ( .A(PCplus4_regI[8]), .B(n168), .S0(n106), .Y(n331) );
  CLKINVX1 U285 ( .A(n152), .Y(n168) );
  MX2XL U286 ( .A(PCplus4_regI[9]), .B(n169), .S0(n92), .Y(n332) );
  CLKINVX1 U287 ( .A(n153), .Y(n169) );
  CLKINVX1 U288 ( .A(n154), .Y(n171) );
  MX2XL U289 ( .A(PCplus4_regI[11]), .B(n355), .S0(n92), .Y(n334) );
  CLKINVX1 U290 ( .A(n155), .Y(n355) );
  MX2XL U291 ( .A(PCplus4_regI[12]), .B(n356), .S0(n92), .Y(n335) );
  CLKINVX1 U292 ( .A(n156), .Y(n356) );
  MX2XL U293 ( .A(PCplus4_regI[13]), .B(n357), .S0(n92), .Y(n336) );
  CLKINVX1 U294 ( .A(n157), .Y(n357) );
  MX2XL U295 ( .A(PCplus4_regI[14]), .B(n358), .S0(n92), .Y(n337) );
  CLKINVX1 U296 ( .A(n158), .Y(n358) );
  MX2XL U297 ( .A(PCplus4_regI[15]), .B(n359), .S0(n92), .Y(n338) );
  CLKINVX1 U298 ( .A(n159), .Y(n359) );
  MX2XL U299 ( .A(PCplus4_regI[16]), .B(n360), .S0(n92), .Y(n339) );
  CLKINVX1 U300 ( .A(n160), .Y(n360) );
  MX2XL U301 ( .A(PCplus4_regI[17]), .B(n361), .S0(n92), .Y(n340) );
  CLKINVX1 U302 ( .A(n161), .Y(n361) );
  MX2XL U303 ( .A(PCplus4_regI[18]), .B(n362), .S0(n92), .Y(n341) );
  CLKINVX1 U304 ( .A(n162), .Y(n362) );
  MX2XL U305 ( .A(PCplus4_regI[19]), .B(n363), .S0(n92), .Y(n342) );
  CLKINVX1 U306 ( .A(n163), .Y(n363) );
  MX2XL U307 ( .A(PCplus4_regI[20]), .B(n364), .S0(n92), .Y(n343) );
  CLKINVX1 U308 ( .A(n164), .Y(n364) );
  MX2XL U309 ( .A(PCplus4_regI[21]), .B(n365), .S0(n92), .Y(n344) );
  CLKINVX1 U310 ( .A(n165), .Y(n365) );
  MX2XL U311 ( .A(PCplus4_regI[22]), .B(n366), .S0(n92), .Y(n345) );
  CLKINVX1 U312 ( .A(n166), .Y(n366) );
  MX2XL U313 ( .A(PCplus4_regI[23]), .B(PCplus4_regD[23]), .S0(n92), .Y(n346)
         );
  MX2XL U314 ( .A(PCplus4_regI[24]), .B(PCplus4_regD[24]), .S0(n92), .Y(n347)
         );
  MX2XL U315 ( .A(PCplus4_regI[25]), .B(PCplus4_regD[25]), .S0(n92), .Y(n348)
         );
  MX2XL U316 ( .A(PCplus4_regI[26]), .B(n367), .S0(n92), .Y(n349) );
  CLKINVX1 U317 ( .A(n170), .Y(n367) );
  MX2XL U318 ( .A(PCplus4_regI[27]), .B(PCplus4_regD[27]), .S0(n92), .Y(n350)
         );
  MX2XL U319 ( .A(PCplus4_regI[28]), .B(n368), .S0(n106), .Y(n351) );
  CLKINVX1 U320 ( .A(n172), .Y(n368) );
  MX2XL U321 ( .A(PCplus4_regI[29]), .B(n369), .S0(n92), .Y(n352) );
  CLKINVX1 U322 ( .A(n173), .Y(n369) );
  MX2XL U323 ( .A(PCplus4_regI[30]), .B(n370), .S0(n92), .Y(n353) );
  CLKINVX1 U324 ( .A(n174), .Y(n370) );
  MX2XL U325 ( .A(PCplus4_regI[31]), .B(n371), .S0(n106), .Y(n354) );
  CLKINVX1 U326 ( .A(n175), .Y(n371) );
  MX2XL U327 ( .A(A[27]), .B(A_regD[27]), .S0(n110), .Y(n284) );
  MX2XL U328 ( .A(A[28]), .B(A_regD[28]), .S0(n110), .Y(n285) );
  MX2XL U329 ( .A(A[29]), .B(A_regD[29]), .S0(n110), .Y(n286) );
  MX2XL U330 ( .A(A[30]), .B(n442), .S0(n110), .Y(n287) );
  CLKINVX1 U331 ( .A(n108), .Y(n442) );
  MX2XL U332 ( .A(A[31]), .B(A_regD[31]), .S0(n110), .Y(n288) );
  CLKMX2X2 U333 ( .A(ALUsrc), .B(ALUsrc_regD), .S0(n106), .Y(n289) );
endmodule


module EX_MEM_regFile ( clk, rst_n, stallcache, MemtoReg_regD, MemRead_regD, 
        MemWrite_regD, RegWrite_regD, B_regD, wsel_regD, ALUout, MemtoReg_regE, 
        MemRead_regE, MemWrite_regE, RegWrite_regE, B_regE, wsel_regE, 
        ALUout_regE );
  input [1:0] MemtoReg_regD;
  input [31:0] B_regD;
  input [4:0] wsel_regD;
  input [31:0] ALUout;
  output [1:0] MemtoReg_regE;
  output [31:0] B_regE;
  output [4:0] wsel_regE;
  output [31:0] ALUout_regE;
  input clk, rst_n, stallcache, MemRead_regD, MemWrite_regD, RegWrite_regD;
  output MemRead_regE, MemWrite_regE, RegWrite_regE;
  wire   n253, n254, n255, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n35, n39, n40, n41, n42, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n1, n33, n34, n36, n37, n38, n43,
         n44, n63, n64, n67, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n167, n168, n206, n208, n210, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n245, n246, n248, n249, n250;

  DFFRX4 \ALUout_regE_reg[31]  ( .D(n144), .CK(clk), .RN(n218), .QN(n70) );
  DFFRX4 \ALUout_regE_reg[26]  ( .D(n139), .CK(clk), .RN(n217), .QN(n65) );
  DFFRX4 \ALUout_regE_reg[21]  ( .D(n134), .CK(clk), .RN(n217), .QN(n60) );
  DFFRX4 \ALUout_regE_reg[11]  ( .D(n124), .CK(clk), .RN(n216), .QN(n50) );
  DFFRX4 \ALUout_regE_reg[9]  ( .D(n122), .CK(clk), .RN(n216), .Q(
        ALUout_regE[9]), .QN(n48) );
  DFFRX4 \ALUout_regE_reg[7]  ( .D(n120), .CK(clk), .RN(n216), .Q(
        ALUout_regE[7]), .QN(n46) );
  DFFRX4 \ALUout_regE_reg[6]  ( .D(n119), .CK(clk), .RN(n216), .Q(
        ALUout_regE[6]), .QN(n45) );
  DFFRX4 \ALUout_regE_reg[3]  ( .D(n116), .CK(clk), .RN(n215), .Q(
        ALUout_regE[3]), .QN(n42) );
  DFFRX4 \ALUout_regE_reg[2]  ( .D(n115), .CK(clk), .RN(n215), .Q(
        ALUout_regE[2]), .QN(n41) );
  DFFRX4 MemWrite_regE_reg ( .D(n104), .CK(clk), .RN(n214), .QN(n35) );
  DFFRX4 \ALUout_regE_reg[5]  ( .D(n118), .CK(clk), .RN(rst_n), .Q(
        ALUout_regE[5]) );
  DFFRX4 \ALUout_regE_reg[4]  ( .D(n117), .CK(clk), .RN(n215), .Q(
        ALUout_regE[4]) );
  DFFRX4 \ALUout_regE_reg[28]  ( .D(n141), .CK(clk), .RN(n217), .Q(n253), .QN(
        n206) );
  DFFRX4 \ALUout_regE_reg[25]  ( .D(n138), .CK(clk), .RN(n217), .Q(n254), .QN(
        n208) );
  DFFRX4 \ALUout_regE_reg[24]  ( .D(n137), .CK(clk), .RN(n217), .Q(n255), .QN(
        n210) );
  DFFRX1 \ALUout_regE_reg[30]  ( .D(n143), .CK(clk), .RN(n218), .Q(
        ALUout_regE[30]), .QN(n69) );
  DFFRX1 \ALUout_regE_reg[29]  ( .D(n142), .CK(clk), .RN(n217), .Q(
        ALUout_regE[29]), .QN(n68) );
  DFFRX1 \ALUout_regE_reg[27]  ( .D(n140), .CK(clk), .RN(n217), .Q(
        ALUout_regE[27]), .QN(n66) );
  DFFRX1 \ALUout_regE_reg[23]  ( .D(n136), .CK(clk), .RN(n217), .Q(
        ALUout_regE[23]), .QN(n62) );
  DFFRX1 \ALUout_regE_reg[19]  ( .D(n132), .CK(clk), .RN(n217), .Q(
        ALUout_regE[19]), .QN(n58) );
  DFFRX1 \ALUout_regE_reg[18]  ( .D(n131), .CK(clk), .RN(n217), .Q(
        ALUout_regE[18]), .QN(n57) );
  DFFRX1 \ALUout_regE_reg[15]  ( .D(n128), .CK(clk), .RN(n216), .Q(
        ALUout_regE[15]), .QN(n54) );
  DFFRX1 \ALUout_regE_reg[13]  ( .D(n126), .CK(clk), .RN(n216), .Q(
        ALUout_regE[13]), .QN(n52) );
  DFFRX1 \ALUout_regE_reg[12]  ( .D(n125), .CK(clk), .RN(n216), .Q(
        ALUout_regE[12]), .QN(n51) );
  DFFRX1 \ALUout_regE_reg[10]  ( .D(n123), .CK(clk), .RN(n216), .Q(
        ALUout_regE[10]), .QN(n49) );
  DFFRX1 \ALUout_regE_reg[22]  ( .D(n135), .CK(clk), .RN(n217), .Q(
        ALUout_regE[22]), .QN(n61) );
  DFFRX1 \ALUout_regE_reg[20]  ( .D(n133), .CK(clk), .RN(n217), .Q(
        ALUout_regE[20]), .QN(n59) );
  DFFRX1 \ALUout_regE_reg[17]  ( .D(n130), .CK(clk), .RN(n216), .Q(
        ALUout_regE[17]), .QN(n56) );
  DFFRX1 \ALUout_regE_reg[16]  ( .D(n129), .CK(clk), .RN(n216), .Q(
        ALUout_regE[16]), .QN(n55) );
  DFFRX1 \ALUout_regE_reg[14]  ( .D(n127), .CK(clk), .RN(n216), .Q(
        ALUout_regE[14]), .QN(n53) );
  DFFRX1 \ALUout_regE_reg[8]  ( .D(n121), .CK(clk), .RN(n216), .Q(
        ALUout_regE[8]), .QN(n47) );
  DFFRX1 \ALUout_regE_reg[0]  ( .D(n113), .CK(clk), .RN(n215), .Q(
        ALUout_regE[0]), .QN(n39) );
  DFFRX1 \ALUout_regE_reg[1]  ( .D(n114), .CK(clk), .RN(n215), .Q(
        ALUout_regE[1]), .QN(n40) );
  DFFRX2 \B_regE_reg[16]  ( .D(n87), .CK(clk), .RN(n213), .Q(n165), .QN(n18)
         );
  DFFRX2 \B_regE_reg[13]  ( .D(n84), .CK(clk), .RN(n213), .Q(n163), .QN(n15)
         );
  DFFRX2 \B_regE_reg[22]  ( .D(n93), .CK(clk), .RN(n213), .Q(n148), .QN(n24)
         );
  DFFRX2 \B_regE_reg[23]  ( .D(n94), .CK(clk), .RN(n213), .Q(n149), .QN(n25)
         );
  DFFRX2 \B_regE_reg[21]  ( .D(n92), .CK(clk), .RN(n213), .Q(n147), .QN(n23)
         );
  DFFRX2 \B_regE_reg[14]  ( .D(n85), .CK(clk), .RN(n213), .Q(n164), .QN(n16)
         );
  DFFRX2 \B_regE_reg[15]  ( .D(n86), .CK(clk), .RN(n213), .Q(n64), .QN(n17) );
  DFFRX2 \B_regE_reg[17]  ( .D(n88), .CK(clk), .RN(n213), .Q(n34), .QN(n19) );
  DFFRX2 \B_regE_reg[18]  ( .D(n89), .CK(clk), .RN(n213), .Q(n67), .QN(n20) );
  DFFRX2 \B_regE_reg[19]  ( .D(n90), .CK(clk), .RN(n213), .Q(n145), .QN(n21)
         );
  DFFRX2 \B_regE_reg[20]  ( .D(n91), .CK(clk), .RN(n213), .Q(n146), .QN(n22)
         );
  DFFRX2 \B_regE_reg[9]  ( .D(n80), .CK(clk), .RN(n212), .Q(n159), .QN(n11) );
  DFFRX2 \B_regE_reg[10]  ( .D(n81), .CK(clk), .RN(n212), .Q(n160), .QN(n12)
         );
  DFFRX2 \B_regE_reg[11]  ( .D(n82), .CK(clk), .RN(n212), .Q(n161), .QN(n13)
         );
  DFFRX2 \B_regE_reg[12]  ( .D(n83), .CK(clk), .RN(n213), .Q(n162), .QN(n14)
         );
  DFFRX2 \B_regE_reg[24]  ( .D(n95), .CK(clk), .RN(n214), .Q(n150), .QN(n26)
         );
  DFFRX2 \B_regE_reg[8]  ( .D(n79), .CK(clk), .RN(n212), .Q(n158), .QN(n10) );
  DFFRX2 \B_regE_reg[27]  ( .D(n98), .CK(clk), .RN(n214), .Q(n153), .QN(n29)
         );
  DFFRX2 \B_regE_reg[28]  ( .D(n99), .CK(clk), .RN(n214), .Q(n43), .QN(n30) );
  DFFRX2 \B_regE_reg[29]  ( .D(n100), .CK(clk), .RN(n214), .Q(n44), .QN(n31)
         );
  DFFRX2 \B_regE_reg[30]  ( .D(n101), .CK(clk), .RN(n214), .Q(n63), .QN(n32)
         );
  DFFRX2 \B_regE_reg[26]  ( .D(n97), .CK(clk), .RN(n214), .Q(n152), .QN(n28)
         );
  DFFRX2 \B_regE_reg[25]  ( .D(n96), .CK(clk), .RN(n214), .Q(n151), .QN(n27)
         );
  DFFRX2 \B_regE_reg[0]  ( .D(n71), .CK(clk), .RN(n212), .Q(n36), .QN(n2) );
  DFFRX2 \B_regE_reg[6]  ( .D(n77), .CK(clk), .RN(n212), .Q(n156), .QN(n8) );
  DFFRX2 \B_regE_reg[7]  ( .D(n78), .CK(clk), .RN(n212), .Q(n157), .QN(n9) );
  DFFRX2 \B_regE_reg[5]  ( .D(n76), .CK(clk), .RN(n212), .Q(n33), .QN(n7) );
  DFFRX2 \B_regE_reg[2]  ( .D(n73), .CK(clk), .RN(n212), .Q(n154), .QN(n4) );
  DFFRX2 \B_regE_reg[3]  ( .D(n74), .CK(clk), .RN(n212), .Q(n38), .QN(n5) );
  DFFRX2 \B_regE_reg[4]  ( .D(n75), .CK(clk), .RN(n212), .Q(n155), .QN(n6) );
  DFFRX2 \B_regE_reg[1]  ( .D(n72), .CK(clk), .RN(n212), .Q(n37), .QN(n3) );
  DFFRHQX8 \wsel_regE_reg[1]  ( .D(n109), .CK(clk), .RN(n215), .Q(wsel_regE[1]) );
  DFFRHQX8 \wsel_regE_reg[3]  ( .D(n111), .CK(clk), .RN(n215), .Q(wsel_regE[3]) );
  DFFRHQX8 \wsel_regE_reg[2]  ( .D(n110), .CK(clk), .RN(n215), .Q(wsel_regE[2]) );
  DFFRHQX8 \wsel_regE_reg[4]  ( .D(n112), .CK(clk), .RN(n215), .Q(wsel_regE[4]) );
  DFFRHQX8 \wsel_regE_reg[0]  ( .D(n108), .CK(clk), .RN(n215), .Q(wsel_regE[0]) );
  DFFRHQX8 RegWrite_regE_reg ( .D(n103), .CK(clk), .RN(n214), .Q(RegWrite_regE) );
  DFFRX1 MemRead_regE_reg ( .D(n105), .CK(clk), .RN(rst_n), .Q(MemRead_regE)
         );
  DFFRX1 \MemtoReg_regE_reg[1]  ( .D(n107), .CK(clk), .RN(n215), .Q(
        MemtoReg_regE[1]) );
  DFFRX1 \MemtoReg_regE_reg[0]  ( .D(n106), .CK(clk), .RN(n214), .Q(
        MemtoReg_regE[0]) );
  DFFRX2 \B_regE_reg[31]  ( .D(n102), .CK(clk), .RN(rst_n), .QN(n1) );
  MX2XL U2 ( .A(ALUout[20]), .B(n243), .S0(n224), .Y(n133) );
  MX2XL U3 ( .A(ALUout[7]), .B(n230), .S0(stallcache), .Y(n120) );
  INVX20 U4 ( .A(n210), .Y(ALUout_regE[24]) );
  INVX16 U5 ( .A(n208), .Y(ALUout_regE[25]) );
  INVX16 U6 ( .A(n206), .Y(ALUout_regE[28]) );
  CLKMX2X2 U7 ( .A(ALUout[24]), .B(n255), .S0(n224), .Y(n137) );
  CLKBUFX3 U8 ( .A(stallcache), .Y(n223) );
  CLKBUFX2 U9 ( .A(rst_n), .Y(n219) );
  CLKBUFX2 U10 ( .A(rst_n), .Y(n220) );
  CLKBUFX3 U11 ( .A(stallcache), .Y(n224) );
  CLKBUFX3 U12 ( .A(stallcache), .Y(n222) );
  BUFX2 U13 ( .A(n222), .Y(n221) );
  INVX16 U14 ( .A(n1), .Y(B_regE[31]) );
  CLKMX2X2 U15 ( .A(wsel_regD[0]), .B(wsel_regE[0]), .S0(stallcache), .Y(n108)
         );
  INVXL U16 ( .A(wsel_regE[1]), .Y(n167) );
  CLKINVX1 U17 ( .A(n167), .Y(n168) );
  MX2XL U18 ( .A(wsel_regD[4]), .B(wsel_regE[4]), .S0(stallcache), .Y(n112) );
  CLKMX2X2 U19 ( .A(wsel_regD[1]), .B(n168), .S0(stallcache), .Y(n109) );
  MX2XL U20 ( .A(ALUout[26]), .B(ALUout_regE[26]), .S0(stallcache), .Y(n139)
         );
  MX2XL U21 ( .A(ALUout[11]), .B(ALUout_regE[11]), .S0(stallcache), .Y(n124)
         );
  CLKMX2X2 U22 ( .A(ALUout[17]), .B(n240), .S0(n224), .Y(n130) );
  MX2XL U23 ( .A(B_regD[5]), .B(n33), .S0(n223), .Y(n76) );
  MX2XL U24 ( .A(B_regD[17]), .B(n34), .S0(n221), .Y(n88) );
  MX2XL U25 ( .A(ALUout[21]), .B(ALUout_regE[21]), .S0(n224), .Y(n134) );
  MX2XL U26 ( .A(B_regD[0]), .B(n36), .S0(stallcache), .Y(n71) );
  CLKMX2X2 U27 ( .A(ALUout[4]), .B(ALUout_regE[4]), .S0(stallcache), .Y(n117)
         );
  CLKMX2X2 U28 ( .A(ALUout[6]), .B(n229), .S0(stallcache), .Y(n119) );
  MX2XL U29 ( .A(B_regD[1]), .B(n37), .S0(stallcache), .Y(n72) );
  CLKMX2X2 U30 ( .A(B_regD[31]), .B(B_regE[31]), .S0(n221), .Y(n102) );
  INVX12 U31 ( .A(n3), .Y(B_regE[1]) );
  INVX12 U32 ( .A(n6), .Y(B_regE[4]) );
  INVX12 U33 ( .A(n5), .Y(B_regE[3]) );
  INVX12 U34 ( .A(n4), .Y(B_regE[2]) );
  INVX12 U35 ( .A(n7), .Y(B_regE[5]) );
  INVX12 U36 ( .A(n9), .Y(B_regE[7]) );
  INVX12 U37 ( .A(n8), .Y(B_regE[6]) );
  INVX12 U38 ( .A(n2), .Y(B_regE[0]) );
  INVX12 U39 ( .A(n27), .Y(B_regE[25]) );
  INVX12 U40 ( .A(n28), .Y(B_regE[26]) );
  INVX12 U41 ( .A(n32), .Y(B_regE[30]) );
  INVX12 U42 ( .A(n31), .Y(B_regE[29]) );
  INVX12 U43 ( .A(n30), .Y(B_regE[28]) );
  INVX12 U44 ( .A(n29), .Y(B_regE[27]) );
  INVX12 U45 ( .A(n10), .Y(B_regE[8]) );
  INVX12 U46 ( .A(n26), .Y(B_regE[24]) );
  INVX12 U47 ( .A(n14), .Y(B_regE[12]) );
  INVX12 U48 ( .A(n13), .Y(B_regE[11]) );
  INVX12 U49 ( .A(n12), .Y(B_regE[10]) );
  INVX12 U50 ( .A(n11), .Y(B_regE[9]) );
  INVX12 U51 ( .A(n22), .Y(B_regE[20]) );
  INVX12 U52 ( .A(n21), .Y(B_regE[19]) );
  INVX12 U53 ( .A(n20), .Y(B_regE[18]) );
  INVX12 U54 ( .A(n19), .Y(B_regE[17]) );
  INVX12 U55 ( .A(n17), .Y(B_regE[15]) );
  INVX12 U56 ( .A(n16), .Y(B_regE[14]) );
  INVX12 U57 ( .A(n23), .Y(B_regE[21]) );
  INVX12 U58 ( .A(n25), .Y(B_regE[23]) );
  INVX12 U59 ( .A(n24), .Y(B_regE[22]) );
  INVX12 U60 ( .A(n15), .Y(B_regE[13]) );
  INVX12 U61 ( .A(n18), .Y(B_regE[16]) );
  INVX20 U62 ( .A(n35), .Y(MemWrite_regE) );
  INVX20 U63 ( .A(n65), .Y(ALUout_regE[26]) );
  INVX20 U64 ( .A(n60), .Y(ALUout_regE[21]) );
  MX2XL U65 ( .A(ALUout[22]), .B(n245), .S0(n224), .Y(n135) );
  MX2XL U66 ( .A(MemRead_regD), .B(MemRead_regE), .S0(n221), .Y(n105) );
  CLKBUFX3 U67 ( .A(n219), .Y(n213) );
  CLKBUFX3 U68 ( .A(n219), .Y(n214) );
  CLKBUFX3 U69 ( .A(n219), .Y(n216) );
  CLKBUFX3 U70 ( .A(n220), .Y(n217) );
  CLKBUFX3 U71 ( .A(n218), .Y(n215) );
  CLKBUFX3 U72 ( .A(n220), .Y(n218) );
  CLKBUFX3 U73 ( .A(n220), .Y(n212) );
  MX2XL U74 ( .A(ALUout[31]), .B(ALUout_regE[31]), .S0(stallcache), .Y(n144)
         );
  CLKINVX1 U75 ( .A(n46), .Y(n230) );
  CLKINVX1 U76 ( .A(n47), .Y(n231) );
  MX2XL U77 ( .A(ALUout[28]), .B(n253), .S0(stallcache), .Y(n141) );
  CLKINVX1 U78 ( .A(n55), .Y(n239) );
  MX2XL U79 ( .A(wsel_regD[2]), .B(wsel_regE[2]), .S0(stallcache), .Y(n110) );
  CLKINVX1 U80 ( .A(n59), .Y(n243) );
  MX2XL U81 ( .A(ALUout[12]), .B(n235), .S0(n224), .Y(n125) );
  CLKINVX1 U82 ( .A(n51), .Y(n235) );
  MX2XL U83 ( .A(B_regD[3]), .B(n38), .S0(n223), .Y(n74) );
  MX2XL U84 ( .A(ALUout[13]), .B(n236), .S0(n224), .Y(n126) );
  CLKINVX1 U85 ( .A(n52), .Y(n236) );
  CLKINVX1 U86 ( .A(n61), .Y(n245) );
  MX2XL U87 ( .A(ALUout[23]), .B(n246), .S0(n224), .Y(n136) );
  CLKINVX1 U88 ( .A(n62), .Y(n246) );
  MX2XL U89 ( .A(wsel_regD[3]), .B(wsel_regE[3]), .S0(stallcache), .Y(n111) );
  MX2XL U90 ( .A(ALUout[9]), .B(n232), .S0(stallcache), .Y(n122) );
  CLKINVX1 U91 ( .A(n48), .Y(n232) );
  CLKINVX1 U92 ( .A(n56), .Y(n240) );
  MX2XL U93 ( .A(B_regD[28]), .B(n43), .S0(n221), .Y(n99) );
  MX2XL U94 ( .A(B_regD[29]), .B(n44), .S0(n221), .Y(n100) );
  MX2XL U95 ( .A(B_regD[30]), .B(n63), .S0(n221), .Y(n101) );
  CLKMX2X2 U96 ( .A(RegWrite_regD), .B(RegWrite_regE), .S0(n221), .Y(n103) );
  CLKMX2X2 U97 ( .A(MemWrite_regD), .B(MemWrite_regE), .S0(n221), .Y(n104) );
  MX2XL U98 ( .A(MemtoReg_regD[0]), .B(MemtoReg_regE[0]), .S0(n221), .Y(n106)
         );
  MX2XL U99 ( .A(MemtoReg_regD[1]), .B(MemtoReg_regE[1]), .S0(n221), .Y(n107)
         );
  MX2XL U100 ( .A(ALUout[14]), .B(n237), .S0(n224), .Y(n127) );
  CLKINVX1 U101 ( .A(n53), .Y(n237) );
  MX2XL U102 ( .A(ALUout[15]), .B(n238), .S0(n224), .Y(n128) );
  CLKINVX1 U103 ( .A(n54), .Y(n238) );
  MX2XL U104 ( .A(ALUout[18]), .B(n241), .S0(n224), .Y(n131) );
  CLKINVX1 U105 ( .A(n57), .Y(n241) );
  MX2XL U106 ( .A(ALUout[19]), .B(n242), .S0(n224), .Y(n132) );
  CLKINVX1 U107 ( .A(n58), .Y(n242) );
  MX2XL U108 ( .A(ALUout[1]), .B(n226), .S0(n224), .Y(n114) );
  CLKINVX1 U109 ( .A(n40), .Y(n226) );
  MX2XL U110 ( .A(ALUout[3]), .B(n228), .S0(stallcache), .Y(n116) );
  CLKINVX1 U111 ( .A(n42), .Y(n228) );
  MX2XL U112 ( .A(ALUout[5]), .B(ALUout_regE[5]), .S0(stallcache), .Y(n118) );
  MX2XL U113 ( .A(ALUout[2]), .B(n227), .S0(stallcache), .Y(n115) );
  CLKINVX1 U114 ( .A(n41), .Y(n227) );
  MX2XL U115 ( .A(ALUout[0]), .B(n225), .S0(stallcache), .Y(n113) );
  CLKINVX1 U116 ( .A(n39), .Y(n225) );
  CLKINVX1 U117 ( .A(n45), .Y(n229) );
  MX2XL U118 ( .A(ALUout[10]), .B(n233), .S0(stallcache), .Y(n123) );
  CLKINVX1 U119 ( .A(n49), .Y(n233) );
  MX2XL U120 ( .A(B_regD[15]), .B(n64), .S0(n222), .Y(n86) );
  MX2XL U121 ( .A(B_regD[18]), .B(n67), .S0(n222), .Y(n89) );
  MX2XL U122 ( .A(B_regD[19]), .B(n145), .S0(n222), .Y(n90) );
  MX2XL U123 ( .A(B_regD[20]), .B(n146), .S0(n223), .Y(n91) );
  MX2XL U124 ( .A(B_regD[21]), .B(n147), .S0(n222), .Y(n92) );
  MX2XL U125 ( .A(B_regD[22]), .B(n148), .S0(n223), .Y(n93) );
  MX2XL U126 ( .A(B_regD[23]), .B(n149), .S0(stallcache), .Y(n94) );
  MX2XL U127 ( .A(B_regD[24]), .B(n150), .S0(n223), .Y(n95) );
  MX2XL U128 ( .A(B_regD[25]), .B(n151), .S0(n222), .Y(n96) );
  MX2XL U129 ( .A(B_regD[26]), .B(n152), .S0(stallcache), .Y(n97) );
  MX2XL U130 ( .A(B_regD[27]), .B(n153), .S0(stallcache), .Y(n98) );
  MX2XL U131 ( .A(B_regD[2]), .B(n154), .S0(n223), .Y(n73) );
  MX2XL U132 ( .A(B_regD[4]), .B(n155), .S0(n223), .Y(n75) );
  MX2XL U133 ( .A(B_regD[6]), .B(n156), .S0(n223), .Y(n77) );
  MX2XL U134 ( .A(B_regD[7]), .B(n157), .S0(n223), .Y(n78) );
  MX2XL U135 ( .A(B_regD[8]), .B(n158), .S0(n223), .Y(n79) );
  MX2XL U136 ( .A(B_regD[9]), .B(n159), .S0(n224), .Y(n80) );
  MX2XL U137 ( .A(B_regD[10]), .B(n160), .S0(n224), .Y(n81) );
  MX2XL U138 ( .A(B_regD[11]), .B(n161), .S0(n223), .Y(n82) );
  MX2XL U139 ( .A(B_regD[12]), .B(n162), .S0(n224), .Y(n83) );
  MX2XL U140 ( .A(B_regD[13]), .B(n163), .S0(n224), .Y(n84) );
  MX2XL U141 ( .A(B_regD[14]), .B(n164), .S0(n222), .Y(n85) );
  MX2XL U142 ( .A(ALUout[27]), .B(n248), .S0(n223), .Y(n140) );
  CLKINVX1 U143 ( .A(n66), .Y(n248) );
  MX2XL U144 ( .A(ALUout[29]), .B(n249), .S0(n223), .Y(n142) );
  CLKINVX1 U145 ( .A(n68), .Y(n249) );
  MX2XL U146 ( .A(ALUout[30]), .B(n250), .S0(stallcache), .Y(n143) );
  CLKINVX1 U147 ( .A(n69), .Y(n250) );
  INVX20 U148 ( .A(n70), .Y(ALUout_regE[31]) );
  INVX20 U149 ( .A(n50), .Y(ALUout_regE[11]) );
  MX2XL U150 ( .A(ALUout[8]), .B(n231), .S0(stallcache), .Y(n121) );
  CLKMX2X2 U151 ( .A(ALUout[16]), .B(n239), .S0(n224), .Y(n129) );
  MX2XL U152 ( .A(B_regD[16]), .B(n165), .S0(stallcache), .Y(n87) );
  MX2XL U153 ( .A(ALUout[25]), .B(n254), .S0(n224), .Y(n138) );
endmodule


module MEM_WB_regFile ( clk, rst_n, stallcache, MemtoReg_regE, RegWrite_regE, 
        ALUout_regE, wsel_regE, dataOut, MemtoReg_regM, RegWrite_regM, 
        ALUout_regM, wsel_regM, dataOut_regM );
  input [1:0] MemtoReg_regE;
  input [31:0] ALUout_regE;
  input [4:0] wsel_regE;
  input [31:0] dataOut;
  output [1:0] MemtoReg_regM;
  output [31:0] ALUout_regM;
  output [4:0] wsel_regM;
  output [31:0] dataOut_regM;
  input clk, rst_n, stallcache, RegWrite_regE;
  output RegWrite_regM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n37, n39, n49, n50, n60, n61, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n64, n65, n66, n67, n68,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n154, n155, n157, n158, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197;

  DFFRX1 \dataOut_regM_reg[23]  ( .D(n132), .CK(clk), .RN(n141), .Q(
        dataOut_regM[23]), .QN(n60) );
  DFFRX1 \dataOut_regM_reg[13]  ( .D(n122), .CK(clk), .RN(n68), .Q(
        dataOut_regM[13]), .QN(n50) );
  DFFRX1 \dataOut_regM_reg[12]  ( .D(n121), .CK(clk), .RN(n68), .Q(
        dataOut_regM[12]), .QN(n49) );
  DFFRX1 \dataOut_regM_reg[2]  ( .D(n111), .CK(clk), .RN(n67), .Q(
        dataOut_regM[2]), .QN(n39) );
  DFFRX1 \ALUout_regM_reg[28]  ( .D(n97), .CK(clk), .RN(n66), .Q(
        ALUout_regM[28]), .QN(n30) );
  DFFRX1 \ALUout_regM_reg[26]  ( .D(n95), .CK(clk), .RN(n66), .Q(
        ALUout_regM[26]), .QN(n28) );
  DFFRX1 \ALUout_regM_reg[25]  ( .D(n94), .CK(clk), .RN(n66), .Q(
        ALUout_regM[25]), .QN(n27) );
  DFFRX1 \ALUout_regM_reg[2]  ( .D(n71), .CK(clk), .RN(n64), .Q(ALUout_regM[2]), .QN(n4) );
  DFFRX1 \ALUout_regM_reg[1]  ( .D(n70), .CK(clk), .RN(n64), .Q(ALUout_regM[1]), .QN(n3) );
  DFFRX1 \dataOut_regM_reg[0]  ( .D(n109), .CK(clk), .RN(n67), .Q(
        dataOut_regM[0]), .QN(n37) );
  DFFRX1 \ALUout_regM_reg[29]  ( .D(n98), .CK(clk), .RN(n66), .Q(
        ALUout_regM[29]), .QN(n31) );
  DFFRX1 \ALUout_regM_reg[27]  ( .D(n96), .CK(clk), .RN(n66), .Q(
        ALUout_regM[27]), .QN(n29) );
  DFFRX1 \ALUout_regM_reg[30]  ( .D(n99), .CK(clk), .RN(n66), .Q(
        ALUout_regM[30]), .QN(n32) );
  DFFRX1 \ALUout_regM_reg[23]  ( .D(n92), .CK(clk), .RN(n65), .Q(
        ALUout_regM[23]), .QN(n25) );
  DFFRX1 \ALUout_regM_reg[19]  ( .D(n88), .CK(clk), .RN(n65), .Q(
        ALUout_regM[19]), .QN(n21) );
  DFFRX1 \ALUout_regM_reg[24]  ( .D(n93), .CK(clk), .RN(n66), .Q(
        ALUout_regM[24]), .QN(n26) );
  DFFRX1 \ALUout_regM_reg[15]  ( .D(n84), .CK(clk), .RN(n65), .Q(
        ALUout_regM[15]), .QN(n17) );
  DFFRX1 \ALUout_regM_reg[22]  ( .D(n91), .CK(clk), .RN(n65), .Q(
        ALUout_regM[22]), .QN(n24) );
  DFFRX1 \ALUout_regM_reg[13]  ( .D(n82), .CK(clk), .RN(n65), .Q(
        ALUout_regM[13]), .QN(n15) );
  DFFRX1 \ALUout_regM_reg[12]  ( .D(n81), .CK(clk), .RN(n65), .Q(
        ALUout_regM[12]), .QN(n14) );
  DFFRX1 \ALUout_regM_reg[20]  ( .D(n89), .CK(clk), .RN(n65), .Q(
        ALUout_regM[20]), .QN(n22) );
  DFFRX1 \ALUout_regM_reg[14]  ( .D(n83), .CK(clk), .RN(n65), .Q(
        ALUout_regM[14]), .QN(n16) );
  DFFRX1 \ALUout_regM_reg[18]  ( .D(n87), .CK(clk), .RN(n65), .Q(
        ALUout_regM[18]), .QN(n20) );
  DFFRX1 \ALUout_regM_reg[21]  ( .D(n90), .CK(clk), .RN(n65), .Q(
        ALUout_regM[21]), .QN(n23) );
  DFFRX1 \ALUout_regM_reg[10]  ( .D(n79), .CK(clk), .RN(n64), .Q(
        ALUout_regM[10]), .QN(n12) );
  DFFRX1 \ALUout_regM_reg[17]  ( .D(n86), .CK(clk), .RN(n65), .Q(
        ALUout_regM[17]), .QN(n19) );
  DFFRX1 \ALUout_regM_reg[11]  ( .D(n80), .CK(clk), .RN(n64), .Q(
        ALUout_regM[11]), .QN(n13) );
  DFFRX1 \ALUout_regM_reg[16]  ( .D(n85), .CK(clk), .RN(n65), .Q(
        ALUout_regM[16]), .QN(n18) );
  DFFRX1 \ALUout_regM_reg[8]  ( .D(n77), .CK(clk), .RN(n64), .Q(ALUout_regM[8]), .QN(n10) );
  DFFRX1 \ALUout_regM_reg[31]  ( .D(n100), .CK(clk), .RN(n66), .Q(
        ALUout_regM[31]), .QN(n33) );
  DFFRX1 \ALUout_regM_reg[0]  ( .D(n69), .CK(clk), .RN(n64), .Q(ALUout_regM[0]), .QN(n2) );
  DFFRX1 \ALUout_regM_reg[9]  ( .D(n78), .CK(clk), .RN(n64), .Q(ALUout_regM[9]), .QN(n11) );
  DFFRX1 \ALUout_regM_reg[7]  ( .D(n76), .CK(clk), .RN(n64), .Q(ALUout_regM[7]), .QN(n9) );
  DFFRX1 \ALUout_regM_reg[6]  ( .D(n75), .CK(clk), .RN(n64), .Q(ALUout_regM[6]), .QN(n8) );
  DFFRX1 \ALUout_regM_reg[5]  ( .D(n74), .CK(clk), .RN(n64), .Q(ALUout_regM[5]), .QN(n7) );
  DFFRX1 \ALUout_regM_reg[4]  ( .D(n73), .CK(clk), .RN(n64), .Q(ALUout_regM[4]), .QN(n6) );
  DFFRHQX8 \wsel_regM_reg[1]  ( .D(n105), .CK(clk), .RN(n67), .Q(wsel_regM[1])
         );
  DFFRHQX8 \wsel_regM_reg[4]  ( .D(n108), .CK(clk), .RN(n67), .Q(wsel_regM[4])
         );
  DFFRHQX8 \wsel_regM_reg[0]  ( .D(n104), .CK(clk), .RN(n66), .Q(wsel_regM[0])
         );
  DFFRHQX8 \wsel_regM_reg[3]  ( .D(n107), .CK(clk), .RN(n67), .Q(wsel_regM[3])
         );
  DFFRHQX8 \wsel_regM_reg[2]  ( .D(n106), .CK(clk), .RN(n67), .Q(wsel_regM[2])
         );
  DFFRHQX8 \MemtoReg_regM_reg[0]  ( .D(n102), .CK(clk), .RN(n66), .Q(
        MemtoReg_regM[0]) );
  DFFRHQX8 \MemtoReg_regM_reg[1]  ( .D(n103), .CK(clk), .RN(n66), .Q(
        MemtoReg_regM[1]) );
  DFFRHQX8 RegWrite_regM_reg ( .D(n101), .CK(clk), .RN(rst_n), .Q(
        RegWrite_regM) );
  DFFRX4 \ALUout_regM_reg[3]  ( .D(n72), .CK(clk), .RN(n64), .Q(ALUout_regM[3]), .QN(n5) );
  DFFRX1 \dataOut_regM_reg[3]  ( .D(n112), .CK(clk), .RN(n67), .Q(
        dataOut_regM[3]) );
  DFFRX1 \dataOut_regM_reg[19]  ( .D(n128), .CK(clk), .RN(n68), .Q(
        dataOut_regM[19]) );
  DFFRX1 \dataOut_regM_reg[31]  ( .D(n140), .CK(clk), .RN(n141), .Q(
        dataOut_regM[31]) );
  DFFRX1 \dataOut_regM_reg[30]  ( .D(n139), .CK(clk), .RN(n141), .Q(
        dataOut_regM[30]) );
  DFFRX1 \dataOut_regM_reg[28]  ( .D(n137), .CK(clk), .RN(n141), .Q(
        dataOut_regM[28]) );
  DFFRX1 \dataOut_regM_reg[27]  ( .D(n136), .CK(clk), .RN(n141), .Q(
        dataOut_regM[27]) );
  DFFSRHQX4 \dataOut_regM_reg[22]  ( .D(n131), .CK(clk), .SN(1'b1), .RN(n141), 
        .Q(dataOut_regM[22]) );
  DFFSRHQX4 \dataOut_regM_reg[21]  ( .D(n130), .CK(clk), .SN(1'b1), .RN(n141), 
        .Q(dataOut_regM[21]) );
  DFFSRHQX4 \dataOut_regM_reg[20]  ( .D(n129), .CK(clk), .SN(1'b1), .RN(n141), 
        .Q(dataOut_regM[20]) );
  DFFSRHQX4 \dataOut_regM_reg[18]  ( .D(n127), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[18]) );
  DFFSRHQX4 \dataOut_regM_reg[17]  ( .D(n126), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[17]) );
  DFFSRHQX4 \dataOut_regM_reg[16]  ( .D(n125), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[16]) );
  DFFSRHQX4 \dataOut_regM_reg[15]  ( .D(n124), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[15]) );
  DFFSRHQX4 \dataOut_regM_reg[14]  ( .D(n123), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[14]) );
  DFFSRHQX4 \dataOut_regM_reg[11]  ( .D(n120), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[11]) );
  DFFSRHQX4 \dataOut_regM_reg[10]  ( .D(n119), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[10]) );
  DFFSRHQX4 \dataOut_regM_reg[9]  ( .D(n118), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[9]) );
  DFFSRHQX4 \dataOut_regM_reg[8]  ( .D(n117), .CK(clk), .SN(1'b1), .RN(n68), 
        .Q(dataOut_regM[8]) );
  DFFSRHQX4 \dataOut_regM_reg[7]  ( .D(n116), .CK(clk), .SN(1'b1), .RN(n67), 
        .Q(dataOut_regM[7]) );
  DFFSRHQX4 \dataOut_regM_reg[6]  ( .D(n115), .CK(clk), .SN(1'b1), .RN(n67), 
        .Q(dataOut_regM[6]) );
  DFFSRHQX4 \dataOut_regM_reg[5]  ( .D(n114), .CK(clk), .SN(1'b1), .RN(n67), 
        .Q(dataOut_regM[5]) );
  DFFSRHQX4 \dataOut_regM_reg[4]  ( .D(n113), .CK(clk), .SN(1'b1), .RN(n67), 
        .Q(dataOut_regM[4]) );
  DFFSRHQX4 \dataOut_regM_reg[1]  ( .D(n110), .CK(clk), .SN(1'b1), .RN(n67), 
        .Q(dataOut_regM[1]) );
  DFFRX2 \dataOut_regM_reg[25]  ( .D(n134), .CK(clk), .RN(n141), .Q(
        dataOut_regM[25]) );
  DFFRX2 \dataOut_regM_reg[26]  ( .D(n135), .CK(clk), .RN(n141), .Q(
        dataOut_regM[26]) );
  DFFRX2 \dataOut_regM_reg[29]  ( .D(n138), .CK(clk), .RN(n141), .Q(
        dataOut_regM[29]) );
  DFFRX4 \dataOut_regM_reg[24]  ( .D(n133), .CK(clk), .RN(n141), .Q(
        dataOut_regM[24]), .QN(n61) );
  BUFX20 U2 ( .A(n149), .Y(n147) );
  BUFX20 U3 ( .A(n150), .Y(n146) );
  CLKMX2X2 U4 ( .A(dataOut[25]), .B(dataOut_regM[25]), .S0(n146), .Y(n134) );
  CLKMX2X2 U5 ( .A(dataOut[14]), .B(dataOut_regM[14]), .S0(n147), .Y(n123) );
  CLKMX2X2 U6 ( .A(dataOut[18]), .B(dataOut_regM[18]), .S0(n146), .Y(n127) );
  CLKMX2X2 U7 ( .A(dataOut[0]), .B(n151), .S0(n144), .Y(n109) );
  CLKMX2X2 U8 ( .A(dataOut[2]), .B(n152), .S0(n144), .Y(n111) );
  CLKMX2X2 U9 ( .A(dataOut[12]), .B(n154), .S0(n144), .Y(n121) );
  CLKMX2X2 U10 ( .A(dataOut[13]), .B(n155), .S0(n147), .Y(n122) );
  CLKMX2X2 U11 ( .A(dataOut[23]), .B(n157), .S0(n146), .Y(n132) );
  CLKBUFX2 U12 ( .A(rst_n), .Y(n143) );
  CLKBUFX2 U13 ( .A(rst_n), .Y(n142) );
  MX2X1 U14 ( .A(dataOut[24]), .B(n158), .S0(n146), .Y(n133) );
  MX2X1 U15 ( .A(dataOut[10]), .B(dataOut_regM[10]), .S0(n144), .Y(n119) );
  MX2X1 U16 ( .A(dataOut[17]), .B(dataOut_regM[17]), .S0(n146), .Y(n126) );
  CLKMX2X2 U17 ( .A(dataOut[21]), .B(dataOut_regM[21]), .S0(n147), .Y(n130) );
  CLKMX2X2 U18 ( .A(dataOut[22]), .B(dataOut_regM[22]), .S0(n146), .Y(n131) );
  CLKMX2X2 U19 ( .A(dataOut[7]), .B(dataOut_regM[7]), .S0(n144), .Y(n116) );
  CLKMX2X2 U20 ( .A(dataOut[20]), .B(dataOut_regM[20]), .S0(n147), .Y(n129) );
  CLKMX2X2 U21 ( .A(dataOut[4]), .B(dataOut_regM[4]), .S0(n144), .Y(n113) );
  CLKMX2X2 U22 ( .A(dataOut[15]), .B(dataOut_regM[15]), .S0(n146), .Y(n124) );
  CLKMX2X2 U23 ( .A(dataOut[1]), .B(dataOut_regM[1]), .S0(n144), .Y(n110) );
  CLKMX2X2 U24 ( .A(dataOut[16]), .B(dataOut_regM[16]), .S0(n147), .Y(n125) );
  CLKMX2X2 U25 ( .A(dataOut[8]), .B(dataOut_regM[8]), .S0(n144), .Y(n117) );
  CLKMX2X2 U26 ( .A(dataOut[11]), .B(dataOut_regM[11]), .S0(n144), .Y(n120) );
  CLKMX2X2 U27 ( .A(dataOut[9]), .B(dataOut_regM[9]), .S0(n144), .Y(n118) );
  CLKMX2X2 U28 ( .A(dataOut[6]), .B(dataOut_regM[6]), .S0(n144), .Y(n115) );
  MX2X1 U29 ( .A(dataOut[31]), .B(dataOut_regM[31]), .S0(n145), .Y(n140) );
  MX2X1 U30 ( .A(dataOut[28]), .B(dataOut_regM[28]), .S0(n145), .Y(n137) );
  MX2X2 U31 ( .A(dataOut[29]), .B(dataOut_regM[29]), .S0(n145), .Y(n138) );
  MX2X2 U32 ( .A(dataOut[26]), .B(dataOut_regM[26]), .S0(n145), .Y(n135) );
  MX2X2 U50 ( .A(dataOut[5]), .B(dataOut_regM[5]), .S0(n144), .Y(n114) );
  MX2X1 U51 ( .A(dataOut[3]), .B(dataOut_regM[3]), .S0(n144), .Y(n112) );
  MX2X1 U52 ( .A(dataOut[19]), .B(dataOut_regM[19]), .S0(n147), .Y(n128) );
  CLKBUFX2 U53 ( .A(n149), .Y(n148) );
  CLKBUFX3 U54 ( .A(n150), .Y(n145) );
  MX2XL U55 ( .A(ALUout_regE[30]), .B(n196), .S0(n148), .Y(n99) );
  MX2XL U56 ( .A(ALUout_regE[31]), .B(n197), .S0(n148), .Y(n100) );
  MX2XL U57 ( .A(ALUout_regE[2]), .B(n168), .S0(n146), .Y(n71) );
  MX2XL U58 ( .A(ALUout_regE[27]), .B(n193), .S0(n147), .Y(n96) );
  MX2XL U59 ( .A(ALUout_regE[12]), .B(n178), .S0(n146), .Y(n81) );
  MX2XL U60 ( .A(ALUout_regE[18]), .B(n184), .S0(n147), .Y(n87) );
  MX2XL U61 ( .A(ALUout_regE[20]), .B(n186), .S0(n147), .Y(n89) );
  MX2XL U62 ( .A(ALUout_regE[13]), .B(n179), .S0(n146), .Y(n82) );
  MX2XL U63 ( .A(ALUout_regE[15]), .B(n181), .S0(n147), .Y(n84) );
  MX2XL U64 ( .A(ALUout_regE[16]), .B(n182), .S0(n147), .Y(n85) );
  MX2XL U65 ( .A(ALUout_regE[11]), .B(n177), .S0(n146), .Y(n80) );
  MX2XL U66 ( .A(ALUout_regE[0]), .B(n166), .S0(n145), .Y(n69) );
  MX2XL U67 ( .A(ALUout_regE[1]), .B(n167), .S0(n145), .Y(n70) );
  CLKBUFX3 U68 ( .A(stallcache), .Y(n144) );
  CLKBUFX3 U69 ( .A(n143), .Y(n64) );
  CLKBUFX3 U70 ( .A(n143), .Y(n65) );
  CLKBUFX3 U71 ( .A(n142), .Y(n67) );
  CLKBUFX3 U72 ( .A(n143), .Y(n68) );
  CLKBUFX3 U73 ( .A(n142), .Y(n141) );
  CLKBUFX3 U74 ( .A(n142), .Y(n66) );
  CLKBUFX3 U75 ( .A(stallcache), .Y(n150) );
  CLKBUFX3 U76 ( .A(stallcache), .Y(n149) );
  CLKINVX1 U77 ( .A(n21), .Y(n185) );
  CLKINVX1 U78 ( .A(n24), .Y(n188) );
  CLKINVX1 U79 ( .A(n10), .Y(n174) );
  CLKINVX1 U80 ( .A(n12), .Y(n176) );
  CLKINVX1 U81 ( .A(n16), .Y(n180) );
  CLKINVX1 U82 ( .A(n11), .Y(n175) );
  CLKINVX1 U83 ( .A(n31), .Y(n195) );
  MX2XL U84 ( .A(ALUout_regE[28]), .B(n194), .S0(n148), .Y(n97) );
  CLKINVX1 U85 ( .A(n30), .Y(n194) );
  MX2XL U86 ( .A(ALUout_regE[25]), .B(n191), .S0(n147), .Y(n94) );
  CLKINVX1 U87 ( .A(n27), .Y(n191) );
  MX2XL U88 ( .A(ALUout_regE[24]), .B(n190), .S0(n147), .Y(n93) );
  CLKINVX1 U89 ( .A(n26), .Y(n190) );
  MX2XL U90 ( .A(ALUout_regE[21]), .B(n187), .S0(n147), .Y(n90) );
  CLKINVX1 U91 ( .A(n23), .Y(n187) );
  MX2XL U92 ( .A(ALUout_regE[26]), .B(n192), .S0(n147), .Y(n95) );
  CLKINVX1 U93 ( .A(n28), .Y(n192) );
  MX2XL U94 ( .A(wsel_regE[1]), .B(wsel_regM[1]), .S0(n145), .Y(n105) );
  CLKINVX1 U95 ( .A(n18), .Y(n182) );
  MX2XL U96 ( .A(ALUout_regE[3]), .B(n169), .S0(n146), .Y(n72) );
  CLKINVX1 U97 ( .A(n5), .Y(n169) );
  CLKINVX1 U98 ( .A(n13), .Y(n177) );
  MX2XL U99 ( .A(wsel_regE[4]), .B(wsel_regM[4]), .S0(n145), .Y(n108) );
  CLKINVX1 U100 ( .A(n4), .Y(n168) );
  CLKINVX1 U101 ( .A(n15), .Y(n179) );
  CLKINVX1 U102 ( .A(n14), .Y(n178) );
  CLKINVX1 U103 ( .A(n17), .Y(n181) );
  CLKINVX1 U104 ( .A(n22), .Y(n186) );
  CLKINVX1 U105 ( .A(n20), .Y(n184) );
  CLKINVX1 U106 ( .A(n29), .Y(n193) );
  MX2XL U107 ( .A(ALUout_regE[23]), .B(n189), .S0(n147), .Y(n92) );
  CLKINVX1 U108 ( .A(n25), .Y(n189) );
  MX2XL U109 ( .A(ALUout_regE[7]), .B(n173), .S0(n146), .Y(n76) );
  CLKINVX1 U110 ( .A(n9), .Y(n173) );
  MX2XL U111 ( .A(ALUout_regE[17]), .B(n183), .S0(n147), .Y(n86) );
  CLKINVX1 U112 ( .A(n19), .Y(n183) );
  CLKINVX1 U113 ( .A(n32), .Y(n196) );
  CLKINVX1 U114 ( .A(n33), .Y(n197) );
  MX2XL U115 ( .A(wsel_regE[3]), .B(wsel_regM[3]), .S0(n145), .Y(n107) );
  MX2XL U116 ( .A(RegWrite_regE), .B(RegWrite_regM), .S0(n148), .Y(n101) );
  MX2XL U117 ( .A(MemtoReg_regE[1]), .B(MemtoReg_regM[1]), .S0(n148), .Y(n103)
         );
  MX2XL U118 ( .A(MemtoReg_regE[0]), .B(MemtoReg_regM[0]), .S0(n148), .Y(n102)
         );
  MX2XL U119 ( .A(ALUout_regE[4]), .B(n170), .S0(n146), .Y(n73) );
  CLKINVX1 U120 ( .A(n6), .Y(n170) );
  MX2XL U121 ( .A(ALUout_regE[5]), .B(n171), .S0(n146), .Y(n74) );
  CLKINVX1 U122 ( .A(n7), .Y(n171) );
  MX2XL U123 ( .A(ALUout_regE[6]), .B(n172), .S0(n146), .Y(n75) );
  CLKINVX1 U124 ( .A(n8), .Y(n172) );
  MX2XL U125 ( .A(dataOut[27]), .B(dataOut_regM[27]), .S0(n145), .Y(n136) );
  MX2XL U126 ( .A(dataOut[30]), .B(dataOut_regM[30]), .S0(n145), .Y(n139) );
  CLKINVX1 U127 ( .A(n2), .Y(n166) );
  CLKINVX1 U128 ( .A(n3), .Y(n167) );
  CLKINVX1 U129 ( .A(n37), .Y(n151) );
  CLKINVX1 U130 ( .A(n39), .Y(n152) );
  CLKINVX1 U131 ( .A(n49), .Y(n154) );
  CLKINVX1 U132 ( .A(n50), .Y(n155) );
  CLKINVX1 U133 ( .A(n60), .Y(n157) );
  CLKINVX1 U134 ( .A(n61), .Y(n158) );
  MX2XL U135 ( .A(ALUout_regE[22]), .B(n188), .S0(n147), .Y(n91) );
  MX2XL U136 ( .A(ALUout_regE[19]), .B(n185), .S0(n147), .Y(n88) );
  MX2XL U137 ( .A(wsel_regE[0]), .B(wsel_regM[0]), .S0(n145), .Y(n104) );
  MX2XL U138 ( .A(wsel_regE[2]), .B(wsel_regM[2]), .S0(n145), .Y(n106) );
  MX2XL U139 ( .A(ALUout_regE[10]), .B(n176), .S0(n146), .Y(n79) );
  MX2X1 U140 ( .A(ALUout_regE[29]), .B(n195), .S0(n148), .Y(n98) );
  MX2XL U141 ( .A(ALUout_regE[8]), .B(n174), .S0(n146), .Y(n77) );
  MX2XL U142 ( .A(ALUout_regE[14]), .B(n180), .S0(n146), .Y(n83) );
  MX2XL U143 ( .A(ALUout_regE[9]), .B(n175), .S0(n146), .Y(n78) );
endmodule


module maincontrol ( opcode, funct, RegDst, MemtoReg, ALUOp, Branch, MemRead, 
        MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp );
  input [5:0] opcode;
  input [5:0] funct;
  output [1:0] RegDst;
  output [1:0] MemtoReg;
  output [5:0] ALUOp;
  output Branch, MemRead, MemWrite, ALUsrc, RegWrite, JumpReg, ExtOp;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n8, n9, n10, n31, n32, n33, n34, n35,
         n36, n37;

  NAND3X2 U3 ( .A(n35), .B(n34), .C(n12), .Y(n17) );
  NAND2X2 U4 ( .A(n10), .B(n17), .Y(RegDst[0]) );
  INVX2 U5 ( .A(opcode[3]), .Y(n34) );
  CLKINVX3 U6 ( .A(opcode[5]), .Y(n31) );
  NAND3X2 U7 ( .A(n10), .B(n15), .C(n19), .Y(MemtoReg[0]) );
  INVX8 U8 ( .A(opcode[1]), .Y(n35) );
  NOR2X4 U9 ( .A(n14), .B(ALUOp[4]), .Y(RegDst[1]) );
  NOR2XL U10 ( .A(ALUOp[4]), .B(n20), .Y(Branch) );
  NOR3XL U11 ( .A(n34), .B(ALUOp[4]), .C(n16), .Y(MemWrite) );
  NOR2XL U12 ( .A(ALUOp[4]), .B(n11), .Y(RegWrite) );
  AND3XL U13 ( .A(funct[3]), .B(n25), .C(n32), .Y(JumpReg) );
  NOR3XL U14 ( .A(n16), .B(ALUOp[4]), .C(opcode[3]), .Y(MemRead) );
  NAND4XL U15 ( .A(n10), .B(n26), .C(n20), .D(n14), .Y(ALUsrc) );
  CLKBUFX2 U16 ( .A(opcode[0]), .Y(ALUOp[0]) );
  CLKBUFX2 U17 ( .A(opcode[1]), .Y(ALUOp[1]) );
  CLKBUFX2 U18 ( .A(opcode[2]), .Y(ALUOp[2]) );
  CLKBUFX2 U19 ( .A(opcode[3]), .Y(ALUOp[3]) );
  CLKBUFX2 U20 ( .A(opcode[5]), .Y(ALUOp[5]) );
  NAND4X2 U21 ( .A(opcode[1]), .B(n24), .C(n34), .D(n31), .Y(n14) );
  NAND3XL U22 ( .A(opcode[2]), .B(n36), .C(n27), .Y(n20) );
  INVX3 U23 ( .A(n20), .Y(n33) );
  NAND3X2 U24 ( .A(n21), .B(n22), .C(funct[3]), .Y(n18) );
  INVX4 U25 ( .A(opcode[0]), .Y(n36) );
  BUFX8 U26 ( .A(opcode[4]), .Y(ALUOp[4]) );
  AOI211XL U27 ( .A0(n12), .A1(n35), .B0(n13), .C0(n8), .Y(n11) );
  INVXL U28 ( .A(n14), .Y(n8) );
  AOI2BB2XL U29 ( .B0(n36), .B1(opcode[3]), .A0N(opcode[1]), .A1N(n23), .Y(n15) );
  NAND3XL U30 ( .A(opcode[1]), .B(n24), .C(opcode[5]), .Y(n16) );
  NOR3XL U31 ( .A(ALUOp[4]), .B(funct[1]), .C(n37), .Y(n25) );
  CLKINVX1 U32 ( .A(n17), .Y(n32) );
  CLKBUFX3 U33 ( .A(RegDst[0]), .Y(ExtOp) );
  OAI31XL U34 ( .A0(n17), .A1(ALUOp[4]), .A2(n18), .B0(n9), .Y(MemtoReg[1]) );
  CLKINVX1 U35 ( .A(RegDst[1]), .Y(n9) );
  CLKINVX1 U36 ( .A(n21), .Y(n37) );
  OAI31XL U37 ( .A0(n37), .A1(funct[3]), .A2(n22), .B0(n32), .Y(n26) );
  NOR3X2 U38 ( .A(opcode[2]), .B(opcode[5]), .C(opcode[0]), .Y(n12) );
  OAI22XL U39 ( .A0(opcode[5]), .A1(n15), .B0(opcode[3]), .B1(n16), .Y(n13) );
  NOR3X1 U40 ( .A(funct[5]), .B(funct[4]), .C(funct[2]), .Y(n21) );
  NOR2X1 U41 ( .A(n36), .B(opcode[2]), .Y(n24) );
  NOR2BX1 U42 ( .AN(funct[0]), .B(funct[1]), .Y(n22) );
  NOR3XL U43 ( .A(opcode[1]), .B(opcode[5]), .C(opcode[3]), .Y(n27) );
  INVX1 U44 ( .A(n28), .Y(n10) );
  OAI221XL U45 ( .A0(n29), .A1(n35), .B0(n24), .B1(n31), .C0(n30), .Y(n28) );
  AOI31XL U46 ( .A0(n23), .A1(n35), .A2(opcode[0]), .B0(ALUOp[4]), .Y(n30) );
  AOI32X1 U47 ( .A0(opcode[0]), .A1(n31), .A2(opcode[3]), .B0(opcode[2]), .B1(
        n34), .Y(n29) );
  NAND2X1 U48 ( .A(opcode[3]), .B(opcode[2]), .Y(n23) );
  AOI221X1 U49 ( .A0(n12), .A1(opcode[1]), .B0(n32), .B1(n18), .C0(n33), .Y(
        n19) );
endmodule


module registerFile ( clk, rst_n, rsel1, rsel2, wsel, wen, wdata, rdata1, 
        rdata2 );
  input [4:0] rsel1;
  input [4:0] rsel2;
  input [4:0] wsel;
  input [31:0] wdata;
  output [31:0] rdata1;
  output [31:0] rdata2;
  input clk, rst_n, wen;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, \register[31][31] ,
         \register[31][30] , \register[31][29] , \register[31][28] ,
         \register[31][27] , \register[31][26] , \register[31][25] ,
         \register[31][24] , \register[31][23] , \register[31][22] ,
         \register[31][21] , \register[31][20] , \register[31][19] ,
         \register[31][18] , \register[31][17] , \register[31][16] ,
         \register[31][15] , \register[31][14] , \register[31][13] ,
         \register[31][12] , \register[31][11] , \register[31][10] ,
         \register[31][9] , \register[31][8] , \register[31][7] ,
         \register[31][6] , \register[31][5] , \register[31][4] ,
         \register[31][3] , \register[31][2] , \register[31][1] ,
         \register[31][0] , \register[30][31] , \register[30][30] ,
         \register[30][29] , \register[30][28] , \register[30][27] ,
         \register[30][26] , \register[30][25] , \register[30][24] ,
         \register[30][23] , \register[30][22] , \register[30][21] ,
         \register[30][20] , \register[30][19] , \register[30][18] ,
         \register[30][17] , \register[30][16] , \register[30][15] ,
         \register[30][14] , \register[30][13] , \register[30][12] ,
         \register[30][11] , \register[30][10] , \register[30][9] ,
         \register[30][8] , \register[30][7] , \register[30][6] ,
         \register[30][5] , \register[30][4] , \register[30][3] ,
         \register[30][2] , \register[30][1] , \register[30][0] ,
         \register[29][31] , \register[29][30] , \register[29][29] ,
         \register[29][28] , \register[29][27] , \register[29][26] ,
         \register[29][25] , \register[29][24] , \register[29][23] ,
         \register[29][22] , \register[29][21] , \register[29][20] ,
         \register[29][19] , \register[29][18] , \register[29][17] ,
         \register[29][16] , \register[29][15] , \register[29][14] ,
         \register[29][13] , \register[29][12] , \register[29][11] ,
         \register[29][10] , \register[29][9] , \register[29][8] ,
         \register[29][7] , \register[29][6] , \register[29][5] ,
         \register[29][4] , \register[29][3] , \register[29][2] ,
         \register[29][1] , \register[29][0] , \register[28][31] ,
         \register[28][30] , \register[28][29] , \register[28][28] ,
         \register[28][27] , \register[28][26] , \register[28][25] ,
         \register[28][24] , \register[28][23] , \register[28][22] ,
         \register[28][21] , \register[28][20] , \register[28][19] ,
         \register[28][18] , \register[28][17] , \register[28][16] ,
         \register[28][15] , \register[28][14] , \register[28][13] ,
         \register[28][12] , \register[28][11] , \register[28][10] ,
         \register[28][9] , \register[28][8] , \register[28][7] ,
         \register[28][6] , \register[28][5] , \register[28][4] ,
         \register[28][3] , \register[28][2] , \register[28][1] ,
         \register[28][0] , \register[27][31] , \register[27][30] ,
         \register[27][29] , \register[27][28] , \register[27][27] ,
         \register[27][26] , \register[27][25] , \register[27][24] ,
         \register[27][23] , \register[27][22] , \register[27][21] ,
         \register[27][20] , \register[27][19] , \register[27][18] ,
         \register[27][17] , \register[27][16] , \register[27][15] ,
         \register[27][14] , \register[27][13] , \register[27][12] ,
         \register[27][11] , \register[27][10] , \register[27][9] ,
         \register[27][8] , \register[27][7] , \register[27][6] ,
         \register[27][5] , \register[27][4] , \register[27][3] ,
         \register[27][2] , \register[27][1] , \register[27][0] ,
         \register[26][31] , \register[26][30] , \register[26][29] ,
         \register[26][28] , \register[26][27] , \register[26][26] ,
         \register[26][25] , \register[26][24] , \register[26][23] ,
         \register[26][22] , \register[26][21] , \register[26][20] ,
         \register[26][19] , \register[26][18] , \register[26][17] ,
         \register[26][16] , \register[26][15] , \register[26][14] ,
         \register[26][13] , \register[26][12] , \register[26][11] ,
         \register[26][10] , \register[26][9] , \register[26][8] ,
         \register[26][7] , \register[26][6] , \register[26][5] ,
         \register[26][4] , \register[26][3] , \register[26][2] ,
         \register[26][1] , \register[26][0] , \register[25][31] ,
         \register[25][30] , \register[25][29] , \register[25][28] ,
         \register[25][27] , \register[25][26] , \register[25][25] ,
         \register[25][24] , \register[25][23] , \register[25][22] ,
         \register[25][21] , \register[25][20] , \register[25][19] ,
         \register[25][18] , \register[25][17] , \register[25][16] ,
         \register[25][15] , \register[25][14] , \register[25][13] ,
         \register[25][12] , \register[25][11] , \register[25][10] ,
         \register[25][9] , \register[25][8] , \register[25][7] ,
         \register[25][6] , \register[25][5] , \register[25][4] ,
         \register[25][3] , \register[25][2] , \register[25][1] ,
         \register[25][0] , \register[24][31] , \register[24][30] ,
         \register[24][29] , \register[24][28] , \register[24][27] ,
         \register[24][26] , \register[24][25] , \register[24][24] ,
         \register[24][23] , \register[24][22] , \register[24][21] ,
         \register[24][20] , \register[24][19] , \register[24][18] ,
         \register[24][17] , \register[24][16] , \register[24][15] ,
         \register[24][14] , \register[24][13] , \register[24][12] ,
         \register[24][11] , \register[24][10] , \register[24][9] ,
         \register[24][8] , \register[24][7] , \register[24][6] ,
         \register[24][5] , \register[24][4] , \register[24][3] ,
         \register[24][2] , \register[24][1] , \register[24][0] ,
         \register[23][31] , \register[23][30] , \register[23][29] ,
         \register[23][28] , \register[23][27] , \register[23][26] ,
         \register[23][25] , \register[23][24] , \register[23][23] ,
         \register[23][22] , \register[23][21] , \register[23][20] ,
         \register[23][19] , \register[23][18] , \register[23][17] ,
         \register[23][16] , \register[23][15] , \register[23][14] ,
         \register[23][13] , \register[23][12] , \register[23][11] ,
         \register[23][10] , \register[23][9] , \register[23][8] ,
         \register[23][7] , \register[23][6] , \register[23][5] ,
         \register[23][4] , \register[23][3] , \register[23][2] ,
         \register[23][1] , \register[23][0] , \register[22][31] ,
         \register[22][30] , \register[22][29] , \register[22][28] ,
         \register[22][27] , \register[22][26] , \register[22][25] ,
         \register[22][24] , \register[22][23] , \register[22][22] ,
         \register[22][21] , \register[22][20] , \register[22][19] ,
         \register[22][18] , \register[22][17] , \register[22][16] ,
         \register[22][15] , \register[22][14] , \register[22][13] ,
         \register[22][12] , \register[22][11] , \register[22][10] ,
         \register[22][9] , \register[22][8] , \register[22][7] ,
         \register[22][6] , \register[22][5] , \register[22][4] ,
         \register[22][3] , \register[22][2] , \register[22][1] ,
         \register[22][0] , \register[21][31] , \register[21][30] ,
         \register[21][29] , \register[21][28] , \register[21][27] ,
         \register[21][26] , \register[21][25] , \register[21][24] ,
         \register[21][23] , \register[21][22] , \register[21][21] ,
         \register[21][20] , \register[21][19] , \register[21][18] ,
         \register[21][17] , \register[21][16] , \register[21][15] ,
         \register[21][14] , \register[21][13] , \register[21][12] ,
         \register[21][11] , \register[21][10] , \register[21][9] ,
         \register[21][8] , \register[21][7] , \register[21][6] ,
         \register[21][5] , \register[21][4] , \register[21][3] ,
         \register[21][2] , \register[21][1] , \register[21][0] ,
         \register[20][31] , \register[20][30] , \register[20][29] ,
         \register[20][28] , \register[20][27] , \register[20][26] ,
         \register[20][25] , \register[20][24] , \register[20][23] ,
         \register[20][22] , \register[20][21] , \register[20][20] ,
         \register[20][19] , \register[20][18] , \register[20][17] ,
         \register[20][16] , \register[20][15] , \register[20][14] ,
         \register[20][13] , \register[20][12] , \register[20][11] ,
         \register[20][10] , \register[20][9] , \register[20][8] ,
         \register[20][7] , \register[20][6] , \register[20][5] ,
         \register[20][4] , \register[20][3] , \register[20][2] ,
         \register[20][1] , \register[20][0] , \register[19][31] ,
         \register[19][30] , \register[19][29] , \register[19][28] ,
         \register[19][27] , \register[19][26] , \register[19][25] ,
         \register[19][24] , \register[19][23] , \register[19][22] ,
         \register[19][21] , \register[19][20] , \register[19][19] ,
         \register[19][18] , \register[19][17] , \register[19][16] ,
         \register[19][15] , \register[19][14] , \register[19][13] ,
         \register[19][12] , \register[19][11] , \register[19][10] ,
         \register[19][9] , \register[19][8] , \register[19][7] ,
         \register[19][6] , \register[19][5] , \register[19][4] ,
         \register[19][3] , \register[19][2] , \register[19][1] ,
         \register[19][0] , \register[18][31] , \register[18][30] ,
         \register[18][29] , \register[18][28] , \register[18][27] ,
         \register[18][26] , \register[18][25] , \register[18][24] ,
         \register[18][23] , \register[18][22] , \register[18][21] ,
         \register[18][20] , \register[18][19] , \register[18][18] ,
         \register[18][17] , \register[18][16] , \register[18][15] ,
         \register[18][14] , \register[18][13] , \register[18][12] ,
         \register[18][11] , \register[18][10] , \register[18][9] ,
         \register[18][8] , \register[18][7] , \register[18][6] ,
         \register[18][5] , \register[18][4] , \register[18][3] ,
         \register[18][2] , \register[18][1] , \register[18][0] ,
         \register[17][31] , \register[17][30] , \register[17][29] ,
         \register[17][28] , \register[17][27] , \register[17][26] ,
         \register[17][25] , \register[17][24] , \register[17][23] ,
         \register[17][22] , \register[17][21] , \register[17][20] ,
         \register[17][19] , \register[17][18] , \register[17][17] ,
         \register[17][16] , \register[17][15] , \register[17][14] ,
         \register[17][13] , \register[17][12] , \register[17][11] ,
         \register[17][10] , \register[17][9] , \register[17][8] ,
         \register[17][7] , \register[17][6] , \register[17][5] ,
         \register[17][4] , \register[17][3] , \register[17][2] ,
         \register[17][1] , \register[17][0] , \register[16][31] ,
         \register[16][30] , \register[16][29] , \register[16][28] ,
         \register[16][27] , \register[16][26] , \register[16][25] ,
         \register[16][24] , \register[16][23] , \register[16][22] ,
         \register[16][21] , \register[16][20] , \register[16][19] ,
         \register[16][18] , \register[16][17] , \register[16][16] ,
         \register[16][15] , \register[16][14] , \register[16][13] ,
         \register[16][12] , \register[16][11] , \register[16][10] ,
         \register[16][9] , \register[16][8] , \register[16][7] ,
         \register[16][6] , \register[16][5] , \register[16][4] ,
         \register[16][3] , \register[16][2] , \register[16][1] ,
         \register[16][0] , \register[15][31] , \register[15][30] ,
         \register[15][29] , \register[15][28] , \register[15][27] ,
         \register[15][26] , \register[15][25] , \register[15][24] ,
         \register[15][23] , \register[15][22] , \register[15][21] ,
         \register[15][20] , \register[15][19] , \register[15][18] ,
         \register[15][17] , \register[15][16] , \register[15][15] ,
         \register[15][14] , \register[15][13] , \register[15][12] ,
         \register[15][11] , \register[15][10] , \register[15][9] ,
         \register[15][8] , \register[15][7] , \register[15][6] ,
         \register[15][5] , \register[15][4] , \register[15][3] ,
         \register[15][2] , \register[15][1] , \register[15][0] ,
         \register[14][31] , \register[14][30] , \register[14][29] ,
         \register[14][28] , \register[14][27] , \register[14][26] ,
         \register[14][25] , \register[14][24] , \register[14][23] ,
         \register[14][22] , \register[14][21] , \register[14][20] ,
         \register[14][19] , \register[14][18] , \register[14][17] ,
         \register[14][16] , \register[14][15] , \register[14][14] ,
         \register[14][13] , \register[14][12] , \register[14][11] ,
         \register[14][10] , \register[14][9] , \register[14][8] ,
         \register[14][7] , \register[14][6] , \register[14][5] ,
         \register[14][4] , \register[14][3] , \register[14][2] ,
         \register[14][1] , \register[14][0] , \register[13][31] ,
         \register[13][30] , \register[13][29] , \register[13][28] ,
         \register[13][27] , \register[13][26] , \register[13][25] ,
         \register[13][24] , \register[13][23] , \register[13][22] ,
         \register[13][21] , \register[13][20] , \register[13][19] ,
         \register[13][18] , \register[13][17] , \register[13][16] ,
         \register[13][15] , \register[13][14] , \register[13][13] ,
         \register[13][12] , \register[13][11] , \register[13][10] ,
         \register[13][9] , \register[13][8] , \register[13][7] ,
         \register[13][6] , \register[13][5] , \register[13][4] ,
         \register[13][3] , \register[13][2] , \register[13][1] ,
         \register[13][0] , \register[12][31] , \register[12][30] ,
         \register[12][29] , \register[12][28] , \register[12][27] ,
         \register[12][26] , \register[12][25] , \register[12][24] ,
         \register[12][23] , \register[12][22] , \register[12][21] ,
         \register[12][20] , \register[12][19] , \register[12][18] ,
         \register[12][17] , \register[12][16] , \register[12][15] ,
         \register[12][14] , \register[12][13] , \register[12][12] ,
         \register[12][11] , \register[12][10] , \register[12][9] ,
         \register[12][8] , \register[12][7] , \register[12][6] ,
         \register[12][5] , \register[12][4] , \register[12][3] ,
         \register[12][2] , \register[12][1] , \register[12][0] ,
         \register[11][31] , \register[11][30] , \register[11][29] ,
         \register[11][28] , \register[11][27] , \register[11][26] ,
         \register[11][25] , \register[11][24] , \register[11][23] ,
         \register[11][22] , \register[11][21] , \register[11][20] ,
         \register[11][19] , \register[11][18] , \register[11][17] ,
         \register[11][16] , \register[11][15] , \register[11][14] ,
         \register[11][13] , \register[11][12] , \register[11][11] ,
         \register[11][10] , \register[11][9] , \register[11][8] ,
         \register[11][7] , \register[11][6] , \register[11][5] ,
         \register[11][4] , \register[11][3] , \register[11][2] ,
         \register[11][1] , \register[11][0] , \register[10][31] ,
         \register[10][30] , \register[10][29] , \register[10][28] ,
         \register[10][27] , \register[10][26] , \register[10][25] ,
         \register[10][24] , \register[10][23] , \register[10][22] ,
         \register[10][21] , \register[10][20] , \register[10][19] ,
         \register[10][18] , \register[10][17] , \register[10][16] ,
         \register[10][15] , \register[10][14] , \register[10][13] ,
         \register[10][12] , \register[10][11] , \register[10][10] ,
         \register[10][9] , \register[10][8] , \register[10][7] ,
         \register[10][6] , \register[10][5] , \register[10][4] ,
         \register[10][3] , \register[10][2] , \register[10][1] ,
         \register[10][0] , \register[9][31] , \register[9][30] ,
         \register[9][29] , \register[9][28] , \register[9][27] ,
         \register[9][26] , \register[9][25] , \register[9][24] ,
         \register[9][23] , \register[9][22] , \register[9][21] ,
         \register[9][20] , \register[9][19] , \register[9][18] ,
         \register[9][17] , \register[9][16] , \register[9][15] ,
         \register[9][14] , \register[9][13] , \register[9][12] ,
         \register[9][11] , \register[9][10] , \register[9][9] ,
         \register[9][8] , \register[9][7] , \register[9][6] ,
         \register[9][5] , \register[9][4] , \register[9][3] ,
         \register[9][2] , \register[9][1] , \register[9][0] ,
         \register[8][31] , \register[8][30] , \register[8][29] ,
         \register[8][28] , \register[8][27] , \register[8][26] ,
         \register[8][25] , \register[8][24] , \register[8][23] ,
         \register[8][22] , \register[8][21] , \register[8][20] ,
         \register[8][19] , \register[8][18] , \register[8][17] ,
         \register[8][16] , \register[8][15] , \register[8][14] ,
         \register[8][13] , \register[8][12] , \register[8][11] ,
         \register[8][10] , \register[8][9] , \register[8][8] ,
         \register[8][7] , \register[8][6] , \register[8][5] ,
         \register[8][4] , \register[8][3] , \register[8][2] ,
         \register[8][1] , \register[8][0] , \register[7][31] ,
         \register[7][30] , \register[7][29] , \register[7][28] ,
         \register[7][27] , \register[7][26] , \register[7][25] ,
         \register[7][24] , \register[7][23] , \register[7][22] ,
         \register[7][21] , \register[7][20] , \register[7][19] ,
         \register[7][18] , \register[7][17] , \register[7][16] ,
         \register[7][15] , \register[7][14] , \register[7][13] ,
         \register[7][12] , \register[7][11] , \register[7][10] ,
         \register[7][9] , \register[7][8] , \register[7][7] ,
         \register[7][6] , \register[7][5] , \register[7][4] ,
         \register[7][3] , \register[7][2] , \register[7][1] ,
         \register[7][0] , \register[6][31] , \register[6][30] ,
         \register[6][29] , \register[6][28] , \register[6][27] ,
         \register[6][26] , \register[6][25] , \register[6][24] ,
         \register[6][23] , \register[6][22] , \register[6][21] ,
         \register[6][20] , \register[6][19] , \register[6][18] ,
         \register[6][17] , \register[6][16] , \register[6][15] ,
         \register[6][14] , \register[6][13] , \register[6][12] ,
         \register[6][11] , \register[6][10] , \register[6][9] ,
         \register[6][8] , \register[6][7] , \register[6][6] ,
         \register[6][5] , \register[6][4] , \register[6][3] ,
         \register[6][2] , \register[6][1] , \register[6][0] ,
         \register[5][31] , \register[5][30] , \register[5][29] ,
         \register[5][28] , \register[5][27] , \register[5][26] ,
         \register[5][25] , \register[5][24] , \register[5][23] ,
         \register[5][22] , \register[5][21] , \register[5][20] ,
         \register[5][19] , \register[5][18] , \register[5][17] ,
         \register[5][16] , \register[5][15] , \register[5][14] ,
         \register[5][13] , \register[5][12] , \register[5][11] ,
         \register[5][10] , \register[5][9] , \register[5][8] ,
         \register[5][7] , \register[5][6] , \register[5][5] ,
         \register[5][4] , \register[5][3] , \register[5][2] ,
         \register[5][1] , \register[5][0] , \register[4][31] ,
         \register[4][30] , \register[4][29] , \register[4][28] ,
         \register[4][27] , \register[4][26] , \register[4][25] ,
         \register[4][24] , \register[4][23] , \register[4][22] ,
         \register[4][21] , \register[4][20] , \register[4][19] ,
         \register[4][18] , \register[4][17] , \register[4][16] ,
         \register[4][15] , \register[4][14] , \register[4][13] ,
         \register[4][12] , \register[4][11] , \register[4][10] ,
         \register[4][9] , \register[4][8] , \register[4][7] ,
         \register[4][6] , \register[4][5] , \register[4][4] ,
         \register[4][3] , \register[4][2] , \register[4][1] ,
         \register[4][0] , \register[3][31] , \register[3][30] ,
         \register[3][29] , \register[3][28] , \register[3][27] ,
         \register[3][26] , \register[3][25] , \register[3][24] ,
         \register[3][23] , \register[3][22] , \register[3][21] ,
         \register[3][20] , \register[3][19] , \register[3][18] ,
         \register[3][17] , \register[3][16] , \register[3][15] ,
         \register[3][14] , \register[3][13] , \register[3][12] ,
         \register[3][11] , \register[3][10] , \register[3][9] ,
         \register[3][8] , \register[3][7] , \register[3][6] ,
         \register[3][5] , \register[3][4] , \register[3][3] ,
         \register[3][2] , \register[3][1] , \register[3][0] ,
         \register[2][31] , \register[2][30] , \register[2][29] ,
         \register[2][28] , \register[2][27] , \register[2][26] ,
         \register[2][25] , \register[2][24] , \register[2][23] ,
         \register[2][22] , \register[2][21] , \register[2][20] ,
         \register[2][19] , \register[2][18] , \register[2][17] ,
         \register[2][16] , \register[2][15] , \register[2][14] ,
         \register[2][13] , \register[2][12] , \register[2][11] ,
         \register[2][10] , \register[2][9] , \register[2][8] ,
         \register[2][7] , \register[2][6] , \register[2][5] ,
         \register[2][4] , \register[2][3] , \register[2][2] ,
         \register[2][1] , \register[2][0] , \register[1][31] ,
         \register[1][30] , \register[1][29] , \register[1][28] ,
         \register[1][27] , \register[1][26] , \register[1][25] ,
         \register[1][24] , \register[1][23] , \register[1][22] ,
         \register[1][21] , \register[1][20] , \register[1][19] ,
         \register[1][18] , \register[1][17] , \register[1][16] ,
         \register[1][15] , \register[1][14] , \register[1][13] ,
         \register[1][12] , \register[1][11] , \register[1][10] ,
         \register[1][9] , \register[1][8] , \register[1][7] ,
         \register[1][6] , \register[1][5] , \register[1][4] ,
         \register[1][3] , \register[1][2] , \register[1][1] ,
         \register[1][0] , N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n68, n69, n70, n71, n72, n73, n75, n76, n77, n79,
         n80, n81, n82, n83, n84, n85, n86, n88, n90, n91, n92, n93, n94, n95,
         n97, n99, n100, n101, n102, n103, n104, n106, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n67, n74,
         n78, n87, n89, n96, n98, n105, n107, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620;
  assign N12 = rsel1[0];
  assign N13 = rsel1[1];
  assign N14 = rsel1[2];
  assign N15 = rsel1[3];
  assign N16 = rsel1[4];
  assign N17 = rsel2[0];
  assign N18 = rsel2[1];
  assign N19 = rsel2[2];
  assign N20 = rsel2[3];
  assign N21 = rsel2[4];

  DFFRX1 \register_reg[2][21]  ( .D(n161), .CK(clk), .RN(n2183), .Q(
        \register[2][21] ), .QN(n2572) );
  DFFRX1 \register_reg[2][20]  ( .D(n160), .CK(clk), .RN(n2183), .Q(
        \register[2][20] ), .QN(n2571) );
  DFFRX1 \register_reg[2][19]  ( .D(n159), .CK(clk), .RN(n2183), .Q(
        \register[2][19] ), .QN(n2570) );
  DFFRX1 \register_reg[2][18]  ( .D(n158), .CK(clk), .RN(n2183), .Q(
        \register[2][18] ), .QN(n2569) );
  DFFRX1 \register_reg[2][17]  ( .D(n157), .CK(clk), .RN(n2183), .Q(
        \register[2][17] ), .QN(n2568) );
  DFFRX1 \register_reg[2][15]  ( .D(n155), .CK(clk), .RN(n2182), .Q(
        \register[2][15] ), .QN(n2566) );
  DFFRX1 \register_reg[2][4]  ( .D(n144), .CK(clk), .RN(n2182), .Q(
        \register[2][4] ), .QN(n2555) );
  DFFRX1 \register_reg[2][2]  ( .D(n142), .CK(clk), .RN(n2188), .Q(
        \register[2][2] ), .QN(n2553) );
  DFFRX1 \register_reg[2][1]  ( .D(n141), .CK(clk), .RN(n2188), .Q(
        \register[2][1] ), .QN(n2552) );
  DFFRX1 \register_reg[2][0]  ( .D(n140), .CK(clk), .RN(n2188), .Q(
        \register[2][0] ), .QN(n2551) );
  DFFRX1 \register_reg[31][31]  ( .D(n1099), .CK(clk), .RN(n2252), .Q(
        \register[31][31] ) );
  DFFRX1 \register_reg[31][30]  ( .D(n1098), .CK(clk), .RN(n2252), .Q(
        \register[31][30] ) );
  DFFRX1 \register_reg[31][29]  ( .D(n1097), .CK(clk), .RN(n2252), .Q(
        \register[31][29] ) );
  DFFRX1 \register_reg[31][28]  ( .D(n1096), .CK(clk), .RN(n2252), .Q(
        \register[31][28] ) );
  DFFRX1 \register_reg[31][27]  ( .D(n1095), .CK(clk), .RN(n2252), .Q(
        \register[31][27] ) );
  DFFRX1 \register_reg[31][26]  ( .D(n1094), .CK(clk), .RN(n2252), .Q(
        \register[31][26] ) );
  DFFRX1 \register_reg[31][25]  ( .D(n1093), .CK(clk), .RN(n2252), .Q(
        \register[31][25] ) );
  DFFRX1 \register_reg[31][24]  ( .D(n1092), .CK(clk), .RN(n2252), .Q(
        \register[31][24] ) );
  DFFRX1 \register_reg[31][23]  ( .D(n1091), .CK(clk), .RN(n2251), .Q(
        \register[31][23] ) );
  DFFRX1 \register_reg[31][22]  ( .D(n1090), .CK(clk), .RN(n2251), .Q(
        \register[31][22] ) );
  DFFRX1 \register_reg[31][21]  ( .D(n1089), .CK(clk), .RN(n2251), .Q(
        \register[31][21] ) );
  DFFRX1 \register_reg[31][20]  ( .D(n1088), .CK(clk), .RN(n2251), .Q(
        \register[31][20] ) );
  DFFRX1 \register_reg[31][19]  ( .D(n1087), .CK(clk), .RN(n2251), .Q(
        \register[31][19] ) );
  DFFRX1 \register_reg[31][18]  ( .D(n1086), .CK(clk), .RN(n2251), .Q(
        \register[31][18] ) );
  DFFRX1 \register_reg[31][17]  ( .D(n1085), .CK(clk), .RN(n2251), .Q(
        \register[31][17] ) );
  DFFRX1 \register_reg[31][16]  ( .D(n1084), .CK(clk), .RN(n2251), .Q(
        \register[31][16] ) );
  DFFRX1 \register_reg[31][15]  ( .D(n1083), .CK(clk), .RN(n2251), .Q(
        \register[31][15] ) );
  DFFRX1 \register_reg[31][14]  ( .D(n1082), .CK(clk), .RN(n2251), .Q(
        \register[31][14] ) );
  DFFRX1 \register_reg[31][13]  ( .D(n1081), .CK(clk), .RN(n2251), .Q(
        \register[31][13] ) );
  DFFRX1 \register_reg[31][12]  ( .D(n1080), .CK(clk), .RN(n2251), .Q(
        \register[31][12] ) );
  DFFRX1 \register_reg[31][11]  ( .D(n1079), .CK(clk), .RN(n2250), .Q(
        \register[31][11] ) );
  DFFRX1 \register_reg[31][10]  ( .D(n1078), .CK(clk), .RN(n2250), .Q(
        \register[31][10] ) );
  DFFRX1 \register_reg[31][9]  ( .D(n1077), .CK(clk), .RN(n2250), .Q(
        \register[31][9] ) );
  DFFRX1 \register_reg[31][8]  ( .D(n1076), .CK(clk), .RN(n2250), .Q(
        \register[31][8] ) );
  DFFRX1 \register_reg[31][7]  ( .D(n1075), .CK(clk), .RN(n2250), .Q(
        \register[31][7] ) );
  DFFRX1 \register_reg[31][6]  ( .D(n1074), .CK(clk), .RN(n2250), .Q(
        \register[31][6] ) );
  DFFRX1 \register_reg[31][5]  ( .D(n1073), .CK(clk), .RN(n2250), .Q(
        \register[31][5] ) );
  DFFRX1 \register_reg[31][4]  ( .D(n1072), .CK(clk), .RN(n2250), .Q(
        \register[31][4] ) );
  DFFRX1 \register_reg[31][3]  ( .D(n1071), .CK(clk), .RN(n2250), .Q(
        \register[31][3] ) );
  DFFRX1 \register_reg[31][2]  ( .D(n1070), .CK(clk), .RN(n2250), .Q(
        \register[31][2] ) );
  DFFRX1 \register_reg[31][1]  ( .D(n1069), .CK(clk), .RN(n2250), .Q(
        \register[31][1] ) );
  DFFRX1 \register_reg[31][0]  ( .D(n1068), .CK(clk), .RN(n2250), .Q(
        \register[31][0] ) );
  DFFRX1 \register_reg[27][31]  ( .D(n971), .CK(clk), .RN(n2256), .Q(
        \register[27][31] ) );
  DFFRX1 \register_reg[27][30]  ( .D(n970), .CK(clk), .RN(n2256), .Q(
        \register[27][30] ) );
  DFFRX1 \register_reg[27][29]  ( .D(n969), .CK(clk), .RN(n2256), .Q(
        \register[27][29] ) );
  DFFRX1 \register_reg[27][28]  ( .D(n968), .CK(clk), .RN(n2256), .Q(
        \register[27][28] ) );
  DFFRX1 \register_reg[27][27]  ( .D(n967), .CK(clk), .RN(n2257), .Q(
        \register[27][27] ) );
  DFFRX1 \register_reg[27][26]  ( .D(n966), .CK(clk), .RN(n2257), .Q(
        \register[27][26] ) );
  DFFRX1 \register_reg[27][25]  ( .D(n965), .CK(clk), .RN(n2257), .Q(
        \register[27][25] ) );
  DFFRX1 \register_reg[27][24]  ( .D(n964), .CK(clk), .RN(n2257), .Q(
        \register[27][24] ) );
  DFFRX1 \register_reg[27][23]  ( .D(n963), .CK(clk), .RN(n2257), .Q(
        \register[27][23] ) );
  DFFRX1 \register_reg[27][22]  ( .D(n962), .CK(clk), .RN(n2257), .Q(
        \register[27][22] ) );
  DFFRX1 \register_reg[27][21]  ( .D(n961), .CK(clk), .RN(n2257), .Q(
        \register[27][21] ) );
  DFFRX1 \register_reg[27][20]  ( .D(n960), .CK(clk), .RN(n2257), .Q(
        \register[27][20] ) );
  DFFRX1 \register_reg[27][19]  ( .D(n959), .CK(clk), .RN(n2240), .Q(
        \register[27][19] ) );
  DFFRX1 \register_reg[27][18]  ( .D(n958), .CK(clk), .RN(n2240), .Q(
        \register[27][18] ) );
  DFFRX1 \register_reg[27][17]  ( .D(n957), .CK(clk), .RN(n2240), .Q(
        \register[27][17] ) );
  DFFRX1 \register_reg[27][16]  ( .D(n956), .CK(clk), .RN(n2240), .Q(
        \register[27][16] ) );
  DFFRX1 \register_reg[27][15]  ( .D(n955), .CK(clk), .RN(n2240), .Q(
        \register[27][15] ) );
  DFFRX1 \register_reg[27][14]  ( .D(n954), .CK(clk), .RN(n2240), .Q(
        \register[27][14] ) );
  DFFRX1 \register_reg[27][13]  ( .D(n953), .CK(clk), .RN(n2240), .Q(
        \register[27][13] ) );
  DFFRX1 \register_reg[27][12]  ( .D(n952), .CK(clk), .RN(n2240), .Q(
        \register[27][12] ) );
  DFFRX1 \register_reg[27][11]  ( .D(n951), .CK(clk), .RN(n2240), .Q(
        \register[27][11] ) );
  DFFRX1 \register_reg[27][10]  ( .D(n950), .CK(clk), .RN(n2240), .Q(
        \register[27][10] ) );
  DFFRX1 \register_reg[27][9]  ( .D(n949), .CK(clk), .RN(n2240), .Q(
        \register[27][9] ) );
  DFFRX1 \register_reg[27][8]  ( .D(n948), .CK(clk), .RN(n2240), .Q(
        \register[27][8] ) );
  DFFRX1 \register_reg[27][7]  ( .D(n947), .CK(clk), .RN(n2239), .Q(
        \register[27][7] ) );
  DFFRX1 \register_reg[27][6]  ( .D(n946), .CK(clk), .RN(n2239), .Q(
        \register[27][6] ) );
  DFFRX1 \register_reg[27][5]  ( .D(n945), .CK(clk), .RN(n2239), .Q(
        \register[27][5] ) );
  DFFRX1 \register_reg[27][4]  ( .D(n944), .CK(clk), .RN(n2239), .Q(
        \register[27][4] ) );
  DFFRX1 \register_reg[27][3]  ( .D(n943), .CK(clk), .RN(n2239), .Q(
        \register[27][3] ) );
  DFFRX1 \register_reg[27][2]  ( .D(n942), .CK(clk), .RN(n2239), .Q(
        \register[27][2] ) );
  DFFRX1 \register_reg[27][1]  ( .D(n941), .CK(clk), .RN(n2239), .Q(
        \register[27][1] ) );
  DFFRX1 \register_reg[27][0]  ( .D(n940), .CK(clk), .RN(n2239), .Q(
        \register[27][0] ) );
  DFFRX1 \register_reg[23][31]  ( .D(n843), .CK(clk), .RN(n2247), .Q(
        \register[23][31] ) );
  DFFRX1 \register_reg[23][30]  ( .D(n842), .CK(clk), .RN(n2247), .Q(
        \register[23][30] ) );
  DFFRX1 \register_reg[23][29]  ( .D(n841), .CK(clk), .RN(n2247), .Q(
        \register[23][29] ) );
  DFFRX1 \register_reg[23][28]  ( .D(n840), .CK(clk), .RN(n2247), .Q(
        \register[23][28] ) );
  DFFRX1 \register_reg[23][27]  ( .D(n839), .CK(clk), .RN(n2246), .Q(
        \register[23][27] ) );
  DFFRX1 \register_reg[23][26]  ( .D(n838), .CK(clk), .RN(n2246), .Q(
        \register[23][26] ) );
  DFFRX1 \register_reg[23][25]  ( .D(n837), .CK(clk), .RN(n2246), .Q(
        \register[23][25] ) );
  DFFRX1 \register_reg[23][24]  ( .D(n836), .CK(clk), .RN(n2246), .Q(
        \register[23][24] ) );
  DFFRX1 \register_reg[23][23]  ( .D(n835), .CK(clk), .RN(n2246), .Q(
        \register[23][23] ) );
  DFFRX1 \register_reg[23][22]  ( .D(n834), .CK(clk), .RN(n2246), .Q(
        \register[23][22] ) );
  DFFRX1 \register_reg[23][21]  ( .D(n833), .CK(clk), .RN(n2246), .Q(
        \register[23][21] ) );
  DFFRX1 \register_reg[23][20]  ( .D(n832), .CK(clk), .RN(n2246), .Q(
        \register[23][20] ) );
  DFFRX1 \register_reg[23][19]  ( .D(n831), .CK(clk), .RN(n2246), .Q(
        \register[23][19] ) );
  DFFRX1 \register_reg[23][18]  ( .D(n830), .CK(clk), .RN(n2246), .Q(
        \register[23][18] ) );
  DFFRX1 \register_reg[23][17]  ( .D(n829), .CK(clk), .RN(n2246), .Q(
        \register[23][17] ) );
  DFFRX1 \register_reg[23][16]  ( .D(n828), .CK(clk), .RN(n2246), .Q(
        \register[23][16] ) );
  DFFRX1 \register_reg[23][15]  ( .D(n827), .CK(clk), .RN(n2245), .Q(
        \register[23][15] ) );
  DFFRX1 \register_reg[23][14]  ( .D(n826), .CK(clk), .RN(n2245), .Q(
        \register[23][14] ) );
  DFFRX1 \register_reg[23][13]  ( .D(n825), .CK(clk), .RN(n2245), .Q(
        \register[23][13] ) );
  DFFRX1 \register_reg[23][12]  ( .D(n824), .CK(clk), .RN(n2245), .Q(
        \register[23][12] ) );
  DFFRX1 \register_reg[23][11]  ( .D(n823), .CK(clk), .RN(n2245), .Q(
        \register[23][11] ) );
  DFFRX1 \register_reg[23][10]  ( .D(n822), .CK(clk), .RN(n2245), .Q(
        \register[23][10] ) );
  DFFRX1 \register_reg[23][9]  ( .D(n821), .CK(clk), .RN(n2245), .Q(
        \register[23][9] ) );
  DFFRX1 \register_reg[23][8]  ( .D(n820), .CK(clk), .RN(n2245), .Q(
        \register[23][8] ) );
  DFFRX1 \register_reg[23][7]  ( .D(n819), .CK(clk), .RN(n2245), .Q(
        \register[23][7] ) );
  DFFRX1 \register_reg[23][6]  ( .D(n818), .CK(clk), .RN(n2245), .Q(
        \register[23][6] ) );
  DFFRX1 \register_reg[23][5]  ( .D(n817), .CK(clk), .RN(n2245), .Q(
        \register[23][5] ) );
  DFFRX1 \register_reg[23][4]  ( .D(n816), .CK(clk), .RN(n2245), .Q(
        \register[23][4] ) );
  DFFRX1 \register_reg[23][3]  ( .D(n815), .CK(clk), .RN(n2228), .Q(
        \register[23][3] ) );
  DFFRX1 \register_reg[23][2]  ( .D(n814), .CK(clk), .RN(n2228), .Q(
        \register[23][2] ) );
  DFFRX1 \register_reg[23][1]  ( .D(n813), .CK(clk), .RN(n2228), .Q(
        \register[23][1] ) );
  DFFRX1 \register_reg[23][0]  ( .D(n812), .CK(clk), .RN(n2228), .Q(
        \register[23][0] ) );
  DFFRX1 \register_reg[19][31]  ( .D(n715), .CK(clk), .RN(n2236), .Q(
        \register[19][31] ) );
  DFFRX1 \register_reg[19][30]  ( .D(n714), .CK(clk), .RN(n2236), .Q(
        \register[19][30] ) );
  DFFRX1 \register_reg[19][29]  ( .D(n713), .CK(clk), .RN(n2236), .Q(
        \register[19][29] ) );
  DFFRX1 \register_reg[19][28]  ( .D(n712), .CK(clk), .RN(n2236), .Q(
        \register[19][28] ) );
  DFFRX1 \register_reg[19][27]  ( .D(n711), .CK(clk), .RN(n2236), .Q(
        \register[19][27] ) );
  DFFRX1 \register_reg[19][26]  ( .D(n710), .CK(clk), .RN(n2236), .Q(
        \register[19][26] ) );
  DFFRX1 \register_reg[19][25]  ( .D(n709), .CK(clk), .RN(n2236), .Q(
        \register[19][25] ) );
  DFFRX1 \register_reg[19][24]  ( .D(n708), .CK(clk), .RN(n2236), .Q(
        \register[19][24] ) );
  DFFRX1 \register_reg[19][23]  ( .D(n707), .CK(clk), .RN(n2235), .Q(
        \register[19][23] ) );
  DFFRX1 \register_reg[19][22]  ( .D(n706), .CK(clk), .RN(n2235), .Q(
        \register[19][22] ) );
  DFFRX1 \register_reg[19][21]  ( .D(n705), .CK(clk), .RN(n2235), .Q(
        \register[19][21] ) );
  DFFRX1 \register_reg[19][20]  ( .D(n704), .CK(clk), .RN(n2235), .Q(
        \register[19][20] ) );
  DFFRX1 \register_reg[19][19]  ( .D(n703), .CK(clk), .RN(n2235), .Q(
        \register[19][19] ) );
  DFFRX1 \register_reg[19][18]  ( .D(n702), .CK(clk), .RN(n2235), .Q(
        \register[19][18] ) );
  DFFRX1 \register_reg[19][17]  ( .D(n701), .CK(clk), .RN(n2235), .Q(
        \register[19][17] ) );
  DFFRX1 \register_reg[19][16]  ( .D(n700), .CK(clk), .RN(n2235), .Q(
        \register[19][16] ) );
  DFFRX1 \register_reg[19][15]  ( .D(n699), .CK(clk), .RN(n2235), .Q(
        \register[19][15] ) );
  DFFRX1 \register_reg[19][14]  ( .D(n698), .CK(clk), .RN(n2235), .Q(
        \register[19][14] ) );
  DFFRX1 \register_reg[19][13]  ( .D(n697), .CK(clk), .RN(n2235), .Q(
        \register[19][13] ) );
  DFFRX1 \register_reg[19][12]  ( .D(n696), .CK(clk), .RN(n2235), .Q(
        \register[19][12] ) );
  DFFRX1 \register_reg[19][11]  ( .D(n695), .CK(clk), .RN(n2234), .Q(
        \register[19][11] ) );
  DFFRX1 \register_reg[19][10]  ( .D(n694), .CK(clk), .RN(n2234), .Q(
        \register[19][10] ) );
  DFFRX1 \register_reg[19][9]  ( .D(n693), .CK(clk), .RN(n2234), .Q(
        \register[19][9] ) );
  DFFRX1 \register_reg[19][8]  ( .D(n692), .CK(clk), .RN(n2234), .Q(
        \register[19][8] ) );
  DFFRX1 \register_reg[19][7]  ( .D(n691), .CK(clk), .RN(n2234), .Q(
        \register[19][7] ) );
  DFFRX1 \register_reg[19][6]  ( .D(n690), .CK(clk), .RN(n2234), .Q(
        \register[19][6] ) );
  DFFRX1 \register_reg[19][5]  ( .D(n689), .CK(clk), .RN(n2234), .Q(
        \register[19][5] ) );
  DFFRX1 \register_reg[19][4]  ( .D(n688), .CK(clk), .RN(n2234), .Q(
        \register[19][4] ) );
  DFFRX1 \register_reg[19][3]  ( .D(n687), .CK(clk), .RN(n2234), .Q(
        \register[19][3] ) );
  DFFRX1 \register_reg[19][2]  ( .D(n686), .CK(clk), .RN(n2234), .Q(
        \register[19][2] ) );
  DFFRX1 \register_reg[19][1]  ( .D(n685), .CK(clk), .RN(n2234), .Q(
        \register[19][1] ) );
  DFFRX1 \register_reg[19][0]  ( .D(n684), .CK(clk), .RN(n2234), .Q(
        \register[19][0] ) );
  DFFRX1 \register_reg[15][31]  ( .D(n587), .CK(clk), .RN(n2217), .Q(
        \register[15][31] ) );
  DFFRX1 \register_reg[15][30]  ( .D(n586), .CK(clk), .RN(n2217), .Q(
        \register[15][30] ) );
  DFFRX1 \register_reg[15][29]  ( .D(n585), .CK(clk), .RN(n2217), .Q(
        \register[15][29] ) );
  DFFRX1 \register_reg[15][28]  ( .D(n584), .CK(clk), .RN(n2217), .Q(
        \register[15][28] ) );
  DFFRX1 \register_reg[15][27]  ( .D(n583), .CK(clk), .RN(n2217), .Q(
        \register[15][27] ) );
  DFFRX1 \register_reg[15][26]  ( .D(n582), .CK(clk), .RN(n2217), .Q(
        \register[15][26] ) );
  DFFRX1 \register_reg[15][25]  ( .D(n581), .CK(clk), .RN(n2217), .Q(
        \register[15][25] ) );
  DFFRX1 \register_reg[15][24]  ( .D(n580), .CK(clk), .RN(n2217), .Q(
        \register[15][24] ) );
  DFFRX1 \register_reg[15][23]  ( .D(n579), .CK(clk), .RN(n2217), .Q(
        \register[15][23] ) );
  DFFRX1 \register_reg[15][22]  ( .D(n578), .CK(clk), .RN(n2217), .Q(
        \register[15][22] ) );
  DFFRX1 \register_reg[15][21]  ( .D(n577), .CK(clk), .RN(n2217), .Q(
        \register[15][21] ) );
  DFFRX1 \register_reg[15][20]  ( .D(n576), .CK(clk), .RN(n2217), .Q(
        \register[15][20] ) );
  DFFRX1 \register_reg[15][19]  ( .D(n575), .CK(clk), .RN(n2224), .Q(
        \register[15][19] ) );
  DFFRX1 \register_reg[15][18]  ( .D(n574), .CK(clk), .RN(n2224), .Q(
        \register[15][18] ) );
  DFFRX1 \register_reg[15][17]  ( .D(n573), .CK(clk), .RN(n2224), .Q(
        \register[15][17] ) );
  DFFRX1 \register_reg[15][16]  ( .D(n572), .CK(clk), .RN(n2224), .Q(
        \register[15][16] ) );
  DFFRX1 \register_reg[15][15]  ( .D(n571), .CK(clk), .RN(n2224), .Q(
        \register[15][15] ) );
  DFFRX1 \register_reg[15][14]  ( .D(n570), .CK(clk), .RN(n2224), .Q(
        \register[15][14] ) );
  DFFRX1 \register_reg[15][13]  ( .D(n569), .CK(clk), .RN(n2224), .Q(
        \register[15][13] ) );
  DFFRX1 \register_reg[15][12]  ( .D(n568), .CK(clk), .RN(n2224), .Q(
        \register[15][12] ) );
  DFFRX1 \register_reg[15][11]  ( .D(n567), .CK(clk), .RN(n2224), .Q(
        \register[15][11] ) );
  DFFRX1 \register_reg[15][10]  ( .D(n566), .CK(clk), .RN(n2224), .Q(
        \register[15][10] ) );
  DFFRX1 \register_reg[15][9]  ( .D(n565), .CK(clk), .RN(n2224), .Q(
        \register[15][9] ) );
  DFFRX1 \register_reg[15][8]  ( .D(n564), .CK(clk), .RN(n2224), .Q(
        \register[15][8] ) );
  DFFRX1 \register_reg[15][7]  ( .D(n563), .CK(clk), .RN(n2223), .Q(
        \register[15][7] ) );
  DFFRX1 \register_reg[15][6]  ( .D(n562), .CK(clk), .RN(n2223), .Q(
        \register[15][6] ) );
  DFFRX1 \register_reg[15][5]  ( .D(n561), .CK(clk), .RN(n2223), .Q(
        \register[15][5] ) );
  DFFRX1 \register_reg[15][4]  ( .D(n560), .CK(clk), .RN(n2223), .Q(
        \register[15][4] ) );
  DFFRX1 \register_reg[15][3]  ( .D(n559), .CK(clk), .RN(n2223), .Q(
        \register[15][3] ) );
  DFFRX1 \register_reg[15][2]  ( .D(n558), .CK(clk), .RN(n2223), .Q(
        \register[15][2] ) );
  DFFRX1 \register_reg[15][1]  ( .D(n557), .CK(clk), .RN(n2223), .Q(
        \register[15][1] ) );
  DFFRX1 \register_reg[15][0]  ( .D(n556), .CK(clk), .RN(n2223), .Q(
        \register[15][0] ) );
  DFFRX1 \register_reg[11][31]  ( .D(n459), .CK(clk), .RN(n2207), .Q(
        \register[11][31] ) );
  DFFRX1 \register_reg[11][30]  ( .D(n458), .CK(clk), .RN(n2207), .Q(
        \register[11][30] ) );
  DFFRX1 \register_reg[11][29]  ( .D(n457), .CK(clk), .RN(n2207), .Q(
        \register[11][29] ) );
  DFFRX1 \register_reg[11][28]  ( .D(n456), .CK(clk), .RN(n2207), .Q(
        \register[11][28] ) );
  DFFRX1 \register_reg[11][27]  ( .D(n455), .CK(clk), .RN(n2206), .Q(
        \register[11][27] ) );
  DFFRX1 \register_reg[11][26]  ( .D(n454), .CK(clk), .RN(n2206), .Q(
        \register[11][26] ) );
  DFFRX1 \register_reg[11][25]  ( .D(n453), .CK(clk), .RN(n2206), .Q(
        \register[11][25] ) );
  DFFRX1 \register_reg[11][24]  ( .D(n452), .CK(clk), .RN(n2206), .Q(
        \register[11][24] ) );
  DFFRX1 \register_reg[11][23]  ( .D(n451), .CK(clk), .RN(n2206), .Q(
        \register[11][23] ) );
  DFFRX1 \register_reg[11][22]  ( .D(n450), .CK(clk), .RN(n2206), .Q(
        \register[11][22] ) );
  DFFRX1 \register_reg[11][21]  ( .D(n449), .CK(clk), .RN(n2206), .Q(
        \register[11][21] ) );
  DFFRX1 \register_reg[11][20]  ( .D(n448), .CK(clk), .RN(n2206), .Q(
        \register[11][20] ) );
  DFFRX1 \register_reg[11][19]  ( .D(n447), .CK(clk), .RN(n2206), .Q(
        \register[11][19] ) );
  DFFRX1 \register_reg[11][18]  ( .D(n446), .CK(clk), .RN(n2206), .Q(
        \register[11][18] ) );
  DFFRX1 \register_reg[11][17]  ( .D(n445), .CK(clk), .RN(n2206), .Q(
        \register[11][17] ) );
  DFFRX1 \register_reg[11][16]  ( .D(n444), .CK(clk), .RN(n2206), .Q(
        \register[11][16] ) );
  DFFRX1 \register_reg[11][15]  ( .D(n443), .CK(clk), .RN(n2205), .Q(
        \register[11][15] ) );
  DFFRX1 \register_reg[11][14]  ( .D(n442), .CK(clk), .RN(n2205), .Q(
        \register[11][14] ) );
  DFFRX1 \register_reg[11][13]  ( .D(n441), .CK(clk), .RN(n2205), .Q(
        \register[11][13] ) );
  DFFRX1 \register_reg[11][12]  ( .D(n440), .CK(clk), .RN(n2205), .Q(
        \register[11][12] ) );
  DFFRX1 \register_reg[11][11]  ( .D(n439), .CK(clk), .RN(n2205), .Q(
        \register[11][11] ) );
  DFFRX1 \register_reg[11][10]  ( .D(n438), .CK(clk), .RN(n2205), .Q(
        \register[11][10] ) );
  DFFRX1 \register_reg[11][9]  ( .D(n437), .CK(clk), .RN(n2205), .Q(
        \register[11][9] ) );
  DFFRX1 \register_reg[11][8]  ( .D(n436), .CK(clk), .RN(n2205), .Q(
        \register[11][8] ) );
  DFFRX1 \register_reg[11][7]  ( .D(n435), .CK(clk), .RN(n2205), .Q(
        \register[11][7] ) );
  DFFRX1 \register_reg[11][6]  ( .D(n434), .CK(clk), .RN(n2205), .Q(
        \register[11][6] ) );
  DFFRX1 \register_reg[11][5]  ( .D(n433), .CK(clk), .RN(n2205), .Q(
        \register[11][5] ) );
  DFFRX1 \register_reg[11][4]  ( .D(n432), .CK(clk), .RN(n2205), .Q(
        \register[11][4] ) );
  DFFRX1 \register_reg[11][3]  ( .D(n431), .CK(clk), .RN(n2212), .Q(
        \register[11][3] ) );
  DFFRX1 \register_reg[11][2]  ( .D(n430), .CK(clk), .RN(n2212), .Q(
        \register[11][2] ) );
  DFFRX1 \register_reg[11][1]  ( .D(n429), .CK(clk), .RN(n2212), .Q(
        \register[11][1] ) );
  DFFRX1 \register_reg[11][0]  ( .D(n428), .CK(clk), .RN(n2212), .Q(
        \register[11][0] ) );
  DFFRX1 \register_reg[7][31]  ( .D(n331), .CK(clk), .RN(n2196), .Q(
        \register[7][31] ) );
  DFFRX1 \register_reg[7][30]  ( .D(n330), .CK(clk), .RN(n2196), .Q(
        \register[7][30] ) );
  DFFRX1 \register_reg[7][29]  ( .D(n329), .CK(clk), .RN(n2196), .Q(
        \register[7][29] ) );
  DFFRX1 \register_reg[7][28]  ( .D(n328), .CK(clk), .RN(n2196), .Q(
        \register[7][28] ) );
  DFFRX1 \register_reg[7][27]  ( .D(n327), .CK(clk), .RN(n2196), .Q(
        \register[7][27] ) );
  DFFRX1 \register_reg[7][26]  ( .D(n326), .CK(clk), .RN(n2196), .Q(
        \register[7][26] ) );
  DFFRX1 \register_reg[7][25]  ( .D(n325), .CK(clk), .RN(n2196), .Q(
        \register[7][25] ) );
  DFFRX1 \register_reg[7][24]  ( .D(n324), .CK(clk), .RN(n2196), .Q(
        \register[7][24] ) );
  DFFRX1 \register_reg[7][23]  ( .D(n323), .CK(clk), .RN(n2195), .Q(
        \register[7][23] ) );
  DFFRX1 \register_reg[7][22]  ( .D(n322), .CK(clk), .RN(n2195), .Q(
        \register[7][22] ) );
  DFFRX1 \register_reg[7][21]  ( .D(n321), .CK(clk), .RN(n2195), .Q(
        \register[7][21] ) );
  DFFRX1 \register_reg[7][20]  ( .D(n320), .CK(clk), .RN(n2195), .Q(
        \register[7][20] ) );
  DFFRX1 \register_reg[7][19]  ( .D(n319), .CK(clk), .RN(n2195), .Q(
        \register[7][19] ) );
  DFFRX1 \register_reg[7][18]  ( .D(n318), .CK(clk), .RN(n2195), .Q(
        \register[7][18] ) );
  DFFRX1 \register_reg[7][17]  ( .D(n317), .CK(clk), .RN(n2195), .Q(
        \register[7][17] ) );
  DFFRX1 \register_reg[7][16]  ( .D(n316), .CK(clk), .RN(n2195), .Q(
        \register[7][16] ) );
  DFFRX1 \register_reg[7][15]  ( .D(n315), .CK(clk), .RN(n2195), .Q(
        \register[7][15] ) );
  DFFRX1 \register_reg[7][14]  ( .D(n314), .CK(clk), .RN(n2195), .Q(
        \register[7][14] ) );
  DFFRX1 \register_reg[7][13]  ( .D(n313), .CK(clk), .RN(n2195), .Q(
        \register[7][13] ) );
  DFFRX1 \register_reg[7][12]  ( .D(n312), .CK(clk), .RN(n2195), .Q(
        \register[7][12] ) );
  DFFRX1 \register_reg[7][11]  ( .D(n311), .CK(clk), .RN(n2194), .Q(
        \register[7][11] ) );
  DFFRX1 \register_reg[7][10]  ( .D(n310), .CK(clk), .RN(n2194), .Q(
        \register[7][10] ) );
  DFFRX1 \register_reg[7][9]  ( .D(n309), .CK(clk), .RN(n2194), .Q(
        \register[7][9] ) );
  DFFRX1 \register_reg[7][8]  ( .D(n308), .CK(clk), .RN(n2194), .Q(
        \register[7][8] ) );
  DFFRX1 \register_reg[7][7]  ( .D(n307), .CK(clk), .RN(n2194), .Q(
        \register[7][7] ) );
  DFFRX1 \register_reg[7][6]  ( .D(n306), .CK(clk), .RN(n2194), .Q(
        \register[7][6] ) );
  DFFRX1 \register_reg[7][5]  ( .D(n305), .CK(clk), .RN(n2194), .Q(
        \register[7][5] ) );
  DFFRX1 \register_reg[7][4]  ( .D(n304), .CK(clk), .RN(n2194), .Q(
        \register[7][4] ) );
  DFFRX1 \register_reg[7][3]  ( .D(n303), .CK(clk), .RN(n2194), .Q(
        \register[7][3] ) );
  DFFRX1 \register_reg[7][2]  ( .D(n302), .CK(clk), .RN(n2194), .Q(
        \register[7][2] ) );
  DFFRX1 \register_reg[7][1]  ( .D(n301), .CK(clk), .RN(n2194), .Q(
        \register[7][1] ) );
  DFFRX1 \register_reg[7][0]  ( .D(n300), .CK(clk), .RN(n2194), .Q(
        \register[7][0] ) );
  DFFRX1 \register_reg[29][31]  ( .D(n1035), .CK(clk), .RN(n2255), .Q(
        \register[29][31] ) );
  DFFRX1 \register_reg[29][30]  ( .D(n1034), .CK(clk), .RN(n2255), .Q(
        \register[29][30] ) );
  DFFRX1 \register_reg[29][29]  ( .D(n1033), .CK(clk), .RN(n2255), .Q(
        \register[29][29] ) );
  DFFRX1 \register_reg[29][28]  ( .D(n1032), .CK(clk), .RN(n2255), .Q(
        \register[29][28] ) );
  DFFRX1 \register_reg[29][27]  ( .D(n1031), .CK(clk), .RN(n2253), .Q(
        \register[29][27] ) );
  DFFRX1 \register_reg[29][26]  ( .D(n1030), .CK(clk), .RN(n2253), .Q(
        \register[29][26] ) );
  DFFRX1 \register_reg[29][25]  ( .D(n1029), .CK(clk), .RN(n2253), .Q(
        \register[29][25] ) );
  DFFRX1 \register_reg[29][24]  ( .D(n1028), .CK(clk), .RN(n2253), .Q(
        \register[29][24] ) );
  DFFRX1 \register_reg[29][23]  ( .D(n1027), .CK(clk), .RN(n2254), .Q(
        \register[29][23] ) );
  DFFRX1 \register_reg[29][22]  ( .D(n1026), .CK(clk), .RN(n2254), .Q(
        \register[29][22] ) );
  DFFRX1 \register_reg[29][21]  ( .D(n1025), .CK(clk), .RN(n2254), .Q(
        \register[29][21] ) );
  DFFRX1 \register_reg[29][20]  ( .D(n1024), .CK(clk), .RN(n2254), .Q(
        \register[29][20] ) );
  DFFRX1 \register_reg[29][19]  ( .D(n1023), .CK(clk), .RN(n2254), .Q(
        \register[29][19] ) );
  DFFRX1 \register_reg[29][18]  ( .D(n1022), .CK(clk), .RN(n2254), .Q(
        \register[29][18] ) );
  DFFRX1 \register_reg[29][17]  ( .D(n1021), .CK(clk), .RN(n2254), .Q(
        \register[29][17] ) );
  DFFRX1 \register_reg[29][16]  ( .D(n1020), .CK(clk), .RN(n2254), .Q(
        \register[29][16] ) );
  DFFRX1 \register_reg[29][15]  ( .D(n1019), .CK(clk), .RN(n2252), .Q(
        \register[29][15] ) );
  DFFRX1 \register_reg[29][14]  ( .D(n1018), .CK(clk), .RN(n2252), .Q(
        \register[29][14] ) );
  DFFRX1 \register_reg[29][13]  ( .D(n1017), .CK(clk), .RN(n2252), .Q(
        \register[29][13] ) );
  DFFRX1 \register_reg[29][12]  ( .D(n1016), .CK(clk), .RN(n2252), .Q(
        \register[29][12] ) );
  DFFRX1 \register_reg[29][11]  ( .D(n1015), .CK(clk), .RN(n2253), .Q(
        \register[29][11] ) );
  DFFRX1 \register_reg[29][10]  ( .D(n1014), .CK(clk), .RN(n2253), .Q(
        \register[29][10] ) );
  DFFRX1 \register_reg[29][9]  ( .D(n1013), .CK(clk), .RN(n2253), .Q(
        \register[29][9] ) );
  DFFRX1 \register_reg[29][8]  ( .D(n1012), .CK(clk), .RN(n2253), .Q(
        \register[29][8] ) );
  DFFRX1 \register_reg[29][7]  ( .D(n1011), .CK(clk), .RN(n2253), .Q(
        \register[29][7] ) );
  DFFRX1 \register_reg[29][6]  ( .D(n1010), .CK(clk), .RN(n2253), .Q(
        \register[29][6] ) );
  DFFRX1 \register_reg[29][5]  ( .D(n1009), .CK(clk), .RN(n2253), .Q(
        \register[29][5] ) );
  DFFRX1 \register_reg[29][4]  ( .D(n1008), .CK(clk), .RN(n2253), .Q(
        \register[29][4] ) );
  DFFRX1 \register_reg[29][3]  ( .D(n1007), .CK(clk), .RN(n2259), .Q(
        \register[29][3] ) );
  DFFRX1 \register_reg[29][2]  ( .D(n1006), .CK(clk), .RN(n2259), .Q(
        \register[29][2] ) );
  DFFRX1 \register_reg[29][1]  ( .D(n1005), .CK(clk), .RN(n2259), .Q(
        \register[29][1] ) );
  DFFRX1 \register_reg[29][0]  ( .D(n1004), .CK(clk), .RN(n2259), .Q(
        \register[29][0] ) );
  DFFRX1 \register_reg[25][31]  ( .D(n907), .CK(clk), .RN(n2244), .Q(
        \register[25][31] ) );
  DFFRX1 \register_reg[25][30]  ( .D(n906), .CK(clk), .RN(n2244), .Q(
        \register[25][30] ) );
  DFFRX1 \register_reg[25][29]  ( .D(n905), .CK(clk), .RN(n2244), .Q(
        \register[25][29] ) );
  DFFRX1 \register_reg[25][28]  ( .D(n904), .CK(clk), .RN(n2244), .Q(
        \register[25][28] ) );
  DFFRX1 \register_reg[25][27]  ( .D(n903), .CK(clk), .RN(n2244), .Q(
        \register[25][27] ) );
  DFFRX1 \register_reg[25][26]  ( .D(n902), .CK(clk), .RN(n2244), .Q(
        \register[25][26] ) );
  DFFRX1 \register_reg[25][25]  ( .D(n901), .CK(clk), .RN(n2244), .Q(
        \register[25][25] ) );
  DFFRX1 \register_reg[25][24]  ( .D(n900), .CK(clk), .RN(n2244), .Q(
        \register[25][24] ) );
  DFFRX1 \register_reg[25][23]  ( .D(n899), .CK(clk), .RN(n2243), .Q(
        \register[25][23] ) );
  DFFRX1 \register_reg[25][22]  ( .D(n898), .CK(clk), .RN(n2243), .Q(
        \register[25][22] ) );
  DFFRX1 \register_reg[25][21]  ( .D(n897), .CK(clk), .RN(n2243), .Q(
        \register[25][21] ) );
  DFFRX1 \register_reg[25][20]  ( .D(n896), .CK(clk), .RN(n2243), .Q(
        \register[25][20] ) );
  DFFRX1 \register_reg[25][19]  ( .D(n895), .CK(clk), .RN(n2243), .Q(
        \register[25][19] ) );
  DFFRX1 \register_reg[25][18]  ( .D(n894), .CK(clk), .RN(n2243), .Q(
        \register[25][18] ) );
  DFFRX1 \register_reg[25][17]  ( .D(n893), .CK(clk), .RN(n2243), .Q(
        \register[25][17] ) );
  DFFRX1 \register_reg[25][16]  ( .D(n892), .CK(clk), .RN(n2243), .Q(
        \register[25][16] ) );
  DFFRX1 \register_reg[25][15]  ( .D(n891), .CK(clk), .RN(n2243), .Q(
        \register[25][15] ) );
  DFFRX1 \register_reg[25][14]  ( .D(n890), .CK(clk), .RN(n2243), .Q(
        \register[25][14] ) );
  DFFRX1 \register_reg[25][13]  ( .D(n889), .CK(clk), .RN(n2243), .Q(
        \register[25][13] ) );
  DFFRX1 \register_reg[25][12]  ( .D(n888), .CK(clk), .RN(n2243), .Q(
        \register[25][12] ) );
  DFFRX1 \register_reg[25][11]  ( .D(n887), .CK(clk), .RN(n2242), .Q(
        \register[25][11] ) );
  DFFRX1 \register_reg[25][10]  ( .D(n886), .CK(clk), .RN(n2242), .Q(
        \register[25][10] ) );
  DFFRX1 \register_reg[25][9]  ( .D(n885), .CK(clk), .RN(n2242), .Q(
        \register[25][9] ) );
  DFFRX1 \register_reg[25][8]  ( .D(n884), .CK(clk), .RN(n2242), .Q(
        \register[25][8] ) );
  DFFRX1 \register_reg[25][7]  ( .D(n883), .CK(clk), .RN(n2242), .Q(
        \register[25][7] ) );
  DFFRX1 \register_reg[25][6]  ( .D(n882), .CK(clk), .RN(n2242), .Q(
        \register[25][6] ) );
  DFFRX1 \register_reg[25][5]  ( .D(n881), .CK(clk), .RN(n2242), .Q(
        \register[25][5] ) );
  DFFRX1 \register_reg[25][4]  ( .D(n880), .CK(clk), .RN(n2242), .Q(
        \register[25][4] ) );
  DFFRX1 \register_reg[25][3]  ( .D(n879), .CK(clk), .RN(n2242), .Q(
        \register[25][3] ) );
  DFFRX1 \register_reg[25][2]  ( .D(n878), .CK(clk), .RN(n2242), .Q(
        \register[25][2] ) );
  DFFRX1 \register_reg[25][1]  ( .D(n877), .CK(clk), .RN(n2242), .Q(
        \register[25][1] ) );
  DFFRX1 \register_reg[25][0]  ( .D(n876), .CK(clk), .RN(n2242), .Q(
        \register[25][0] ) );
  DFFRX1 \register_reg[21][31]  ( .D(n779), .CK(clk), .RN(n2225), .Q(
        \register[21][31] ) );
  DFFRX1 \register_reg[21][30]  ( .D(n778), .CK(clk), .RN(n2225), .Q(
        \register[21][30] ) );
  DFFRX1 \register_reg[21][29]  ( .D(n777), .CK(clk), .RN(n2225), .Q(
        \register[21][29] ) );
  DFFRX1 \register_reg[21][28]  ( .D(n776), .CK(clk), .RN(n2225), .Q(
        \register[21][28] ) );
  DFFRX1 \register_reg[21][27]  ( .D(n775), .CK(clk), .RN(n2225), .Q(
        \register[21][27] ) );
  DFFRX1 \register_reg[21][26]  ( .D(n774), .CK(clk), .RN(n2225), .Q(
        \register[21][26] ) );
  DFFRX1 \register_reg[21][25]  ( .D(n773), .CK(clk), .RN(n2225), .Q(
        \register[21][25] ) );
  DFFRX1 \register_reg[21][24]  ( .D(n772), .CK(clk), .RN(n2225), .Q(
        \register[21][24] ) );
  DFFRX1 \register_reg[21][23]  ( .D(n771), .CK(clk), .RN(n2225), .Q(
        \register[21][23] ) );
  DFFRX1 \register_reg[21][22]  ( .D(n770), .CK(clk), .RN(n2225), .Q(
        \register[21][22] ) );
  DFFRX1 \register_reg[21][21]  ( .D(n769), .CK(clk), .RN(n2225), .Q(
        \register[21][21] ) );
  DFFRX1 \register_reg[21][20]  ( .D(n768), .CK(clk), .RN(n2225), .Q(
        \register[21][20] ) );
  DFFRX1 \register_reg[21][19]  ( .D(n767), .CK(clk), .RN(n2232), .Q(
        \register[21][19] ) );
  DFFRX1 \register_reg[21][18]  ( .D(n766), .CK(clk), .RN(n2232), .Q(
        \register[21][18] ) );
  DFFRX1 \register_reg[21][17]  ( .D(n765), .CK(clk), .RN(n2232), .Q(
        \register[21][17] ) );
  DFFRX1 \register_reg[21][16]  ( .D(n764), .CK(clk), .RN(n2232), .Q(
        \register[21][16] ) );
  DFFRX1 \register_reg[21][15]  ( .D(n763), .CK(clk), .RN(n2232), .Q(
        \register[21][15] ) );
  DFFRX1 \register_reg[21][14]  ( .D(n762), .CK(clk), .RN(n2232), .Q(
        \register[21][14] ) );
  DFFRX1 \register_reg[21][13]  ( .D(n761), .CK(clk), .RN(n2232), .Q(
        \register[21][13] ) );
  DFFRX1 \register_reg[21][12]  ( .D(n760), .CK(clk), .RN(n2232), .Q(
        \register[21][12] ) );
  DFFRX1 \register_reg[21][11]  ( .D(n759), .CK(clk), .RN(n2232), .Q(
        \register[21][11] ) );
  DFFRX1 \register_reg[21][10]  ( .D(n758), .CK(clk), .RN(n2232), .Q(
        \register[21][10] ) );
  DFFRX1 \register_reg[21][9]  ( .D(n757), .CK(clk), .RN(n2232), .Q(
        \register[21][9] ) );
  DFFRX1 \register_reg[21][8]  ( .D(n756), .CK(clk), .RN(n2232), .Q(
        \register[21][8] ) );
  DFFRX1 \register_reg[21][7]  ( .D(n755), .CK(clk), .RN(n2231), .Q(
        \register[21][7] ) );
  DFFRX1 \register_reg[21][6]  ( .D(n754), .CK(clk), .RN(n2231), .Q(
        \register[21][6] ) );
  DFFRX1 \register_reg[21][5]  ( .D(n753), .CK(clk), .RN(n2231), .Q(
        \register[21][5] ) );
  DFFRX1 \register_reg[21][4]  ( .D(n752), .CK(clk), .RN(n2231), .Q(
        \register[21][4] ) );
  DFFRX1 \register_reg[21][3]  ( .D(n751), .CK(clk), .RN(n2231), .Q(
        \register[21][3] ) );
  DFFRX1 \register_reg[21][2]  ( .D(n750), .CK(clk), .RN(n2231), .Q(
        \register[21][2] ) );
  DFFRX1 \register_reg[21][1]  ( .D(n749), .CK(clk), .RN(n2231), .Q(
        \register[21][1] ) );
  DFFRX1 \register_reg[21][0]  ( .D(n748), .CK(clk), .RN(n2231), .Q(
        \register[21][0] ) );
  DFFRX1 \register_reg[17][31]  ( .D(n651), .CK(clk), .RN(n2215), .Q(
        \register[17][31] ) );
  DFFRX1 \register_reg[17][30]  ( .D(n650), .CK(clk), .RN(n2215), .Q(
        \register[17][30] ) );
  DFFRX1 \register_reg[17][29]  ( .D(n649), .CK(clk), .RN(n2215), .Q(
        \register[17][29] ) );
  DFFRX1 \register_reg[17][28]  ( .D(n648), .CK(clk), .RN(n2215), .Q(
        \register[17][28] ) );
  DFFRX1 \register_reg[17][27]  ( .D(n647), .CK(clk), .RN(n2214), .Q(
        \register[17][27] ) );
  DFFRX1 \register_reg[17][26]  ( .D(n646), .CK(clk), .RN(n2214), .Q(
        \register[17][26] ) );
  DFFRX1 \register_reg[17][25]  ( .D(n645), .CK(clk), .RN(n2214), .Q(
        \register[17][25] ) );
  DFFRX1 \register_reg[17][24]  ( .D(n644), .CK(clk), .RN(n2214), .Q(
        \register[17][24] ) );
  DFFRX1 \register_reg[17][23]  ( .D(n643), .CK(clk), .RN(n2214), .Q(
        \register[17][23] ) );
  DFFRX1 \register_reg[17][22]  ( .D(n642), .CK(clk), .RN(n2214), .Q(
        \register[17][22] ) );
  DFFRX1 \register_reg[17][21]  ( .D(n641), .CK(clk), .RN(n2214), .Q(
        \register[17][21] ) );
  DFFRX1 \register_reg[17][20]  ( .D(n640), .CK(clk), .RN(n2214), .Q(
        \register[17][20] ) );
  DFFRX1 \register_reg[17][19]  ( .D(n639), .CK(clk), .RN(n2214), .Q(
        \register[17][19] ) );
  DFFRX1 \register_reg[17][18]  ( .D(n638), .CK(clk), .RN(n2214), .Q(
        \register[17][18] ) );
  DFFRX1 \register_reg[17][17]  ( .D(n637), .CK(clk), .RN(n2214), .Q(
        \register[17][17] ) );
  DFFRX1 \register_reg[17][16]  ( .D(n636), .CK(clk), .RN(n2214), .Q(
        \register[17][16] ) );
  DFFRX1 \register_reg[17][15]  ( .D(n635), .CK(clk), .RN(n2213), .Q(
        \register[17][15] ) );
  DFFRX1 \register_reg[17][14]  ( .D(n634), .CK(clk), .RN(n2213), .Q(
        \register[17][14] ) );
  DFFRX1 \register_reg[17][13]  ( .D(n633), .CK(clk), .RN(n2213), .Q(
        \register[17][13] ) );
  DFFRX1 \register_reg[17][12]  ( .D(n632), .CK(clk), .RN(n2213), .Q(
        \register[17][12] ) );
  DFFRX1 \register_reg[17][11]  ( .D(n631), .CK(clk), .RN(n2213), .Q(
        \register[17][11] ) );
  DFFRX1 \register_reg[17][10]  ( .D(n630), .CK(clk), .RN(n2213), .Q(
        \register[17][10] ) );
  DFFRX1 \register_reg[17][9]  ( .D(n629), .CK(clk), .RN(n2213), .Q(
        \register[17][9] ) );
  DFFRX1 \register_reg[17][8]  ( .D(n628), .CK(clk), .RN(n2213), .Q(
        \register[17][8] ) );
  DFFRX1 \register_reg[17][7]  ( .D(n627), .CK(clk), .RN(n2213), .Q(
        \register[17][7] ) );
  DFFRX1 \register_reg[17][6]  ( .D(n626), .CK(clk), .RN(n2213), .Q(
        \register[17][6] ) );
  DFFRX1 \register_reg[17][5]  ( .D(n625), .CK(clk), .RN(n2213), .Q(
        \register[17][5] ) );
  DFFRX1 \register_reg[17][4]  ( .D(n624), .CK(clk), .RN(n2213), .Q(
        \register[17][4] ) );
  DFFRX1 \register_reg[17][3]  ( .D(n623), .CK(clk), .RN(n2220), .Q(
        \register[17][3] ) );
  DFFRX1 \register_reg[17][2]  ( .D(n622), .CK(clk), .RN(n2220), .Q(
        \register[17][2] ) );
  DFFRX1 \register_reg[17][1]  ( .D(n621), .CK(clk), .RN(n2220), .Q(
        \register[17][1] ) );
  DFFRX1 \register_reg[17][0]  ( .D(n620), .CK(clk), .RN(n2220), .Q(
        \register[17][0] ) );
  DFFRX1 \register_reg[13][31]  ( .D(n523), .CK(clk), .RN(n2204), .Q(
        \register[13][31] ) );
  DFFRX1 \register_reg[13][30]  ( .D(n522), .CK(clk), .RN(n2204), .Q(
        \register[13][30] ) );
  DFFRX1 \register_reg[13][29]  ( .D(n521), .CK(clk), .RN(n2204), .Q(
        \register[13][29] ) );
  DFFRX1 \register_reg[13][28]  ( .D(n520), .CK(clk), .RN(n2204), .Q(
        \register[13][28] ) );
  DFFRX1 \register_reg[13][27]  ( .D(n519), .CK(clk), .RN(n2204), .Q(
        \register[13][27] ) );
  DFFRX1 \register_reg[13][26]  ( .D(n518), .CK(clk), .RN(n2204), .Q(
        \register[13][26] ) );
  DFFRX1 \register_reg[13][25]  ( .D(n517), .CK(clk), .RN(n2204), .Q(
        \register[13][25] ) );
  DFFRX1 \register_reg[13][24]  ( .D(n516), .CK(clk), .RN(n2204), .Q(
        \register[13][24] ) );
  DFFRX1 \register_reg[13][23]  ( .D(n515), .CK(clk), .RN(n2203), .Q(
        \register[13][23] ) );
  DFFRX1 \register_reg[13][22]  ( .D(n514), .CK(clk), .RN(n2203), .Q(
        \register[13][22] ) );
  DFFRX1 \register_reg[13][21]  ( .D(n513), .CK(clk), .RN(n2203), .Q(
        \register[13][21] ) );
  DFFRX1 \register_reg[13][20]  ( .D(n512), .CK(clk), .RN(n2203), .Q(
        \register[13][20] ) );
  DFFRX1 \register_reg[13][19]  ( .D(n511), .CK(clk), .RN(n2203), .Q(
        \register[13][19] ) );
  DFFRX1 \register_reg[13][18]  ( .D(n510), .CK(clk), .RN(n2203), .Q(
        \register[13][18] ) );
  DFFRX1 \register_reg[13][17]  ( .D(n509), .CK(clk), .RN(n2203), .Q(
        \register[13][17] ) );
  DFFRX1 \register_reg[13][16]  ( .D(n508), .CK(clk), .RN(n2203), .Q(
        \register[13][16] ) );
  DFFRX1 \register_reg[13][15]  ( .D(n507), .CK(clk), .RN(n2203), .Q(
        \register[13][15] ) );
  DFFRX1 \register_reg[13][14]  ( .D(n506), .CK(clk), .RN(n2203), .Q(
        \register[13][14] ) );
  DFFRX1 \register_reg[13][13]  ( .D(n505), .CK(clk), .RN(n2203), .Q(
        \register[13][13] ) );
  DFFRX1 \register_reg[13][12]  ( .D(n504), .CK(clk), .RN(n2203), .Q(
        \register[13][12] ) );
  DFFRX1 \register_reg[13][11]  ( .D(n503), .CK(clk), .RN(n2202), .Q(
        \register[13][11] ) );
  DFFRX1 \register_reg[13][10]  ( .D(n502), .CK(clk), .RN(n2202), .Q(
        \register[13][10] ) );
  DFFRX1 \register_reg[13][9]  ( .D(n501), .CK(clk), .RN(n2202), .Q(
        \register[13][9] ) );
  DFFRX1 \register_reg[13][8]  ( .D(n500), .CK(clk), .RN(n2202), .Q(
        \register[13][8] ) );
  DFFRX1 \register_reg[13][7]  ( .D(n499), .CK(clk), .RN(n2202), .Q(
        \register[13][7] ) );
  DFFRX1 \register_reg[13][6]  ( .D(n498), .CK(clk), .RN(n2202), .Q(
        \register[13][6] ) );
  DFFRX1 \register_reg[13][5]  ( .D(n497), .CK(clk), .RN(n2202), .Q(
        \register[13][5] ) );
  DFFRX1 \register_reg[13][4]  ( .D(n496), .CK(clk), .RN(n2202), .Q(
        \register[13][4] ) );
  DFFRX1 \register_reg[13][3]  ( .D(n495), .CK(clk), .RN(n2202), .Q(
        \register[13][3] ) );
  DFFRX1 \register_reg[13][2]  ( .D(n494), .CK(clk), .RN(n2202), .Q(
        \register[13][2] ) );
  DFFRX1 \register_reg[13][1]  ( .D(n493), .CK(clk), .RN(n2202), .Q(
        \register[13][1] ) );
  DFFRX1 \register_reg[13][0]  ( .D(n492), .CK(clk), .RN(n2202), .Q(
        \register[13][0] ) );
  DFFRX1 \register_reg[9][31]  ( .D(n395), .CK(clk), .RN(n2209), .Q(
        \register[9][31] ) );
  DFFRX1 \register_reg[9][30]  ( .D(n394), .CK(clk), .RN(n2209), .Q(
        \register[9][30] ) );
  DFFRX1 \register_reg[9][29]  ( .D(n393), .CK(clk), .RN(n2209), .Q(
        \register[9][29] ) );
  DFFRX1 \register_reg[9][28]  ( .D(n392), .CK(clk), .RN(n2209), .Q(
        \register[9][28] ) );
  DFFRX1 \register_reg[9][27]  ( .D(n391), .CK(clk), .RN(n2209), .Q(
        \register[9][27] ) );
  DFFRX1 \register_reg[9][26]  ( .D(n390), .CK(clk), .RN(n2209), .Q(
        \register[9][26] ) );
  DFFRX1 \register_reg[9][25]  ( .D(n389), .CK(clk), .RN(n2209), .Q(
        \register[9][25] ) );
  DFFRX1 \register_reg[9][24]  ( .D(n388), .CK(clk), .RN(n2209), .Q(
        \register[9][24] ) );
  DFFRX1 \register_reg[9][23]  ( .D(n387), .CK(clk), .RN(n2209), .Q(
        \register[9][23] ) );
  DFFRX1 \register_reg[9][22]  ( .D(n386), .CK(clk), .RN(n2209), .Q(
        \register[9][22] ) );
  DFFRX1 \register_reg[9][21]  ( .D(n385), .CK(clk), .RN(n2209), .Q(
        \register[9][21] ) );
  DFFRX1 \register_reg[9][20]  ( .D(n384), .CK(clk), .RN(n2209), .Q(
        \register[9][20] ) );
  DFFRX1 \register_reg[9][19]  ( .D(n383), .CK(clk), .RN(n2192), .Q(
        \register[9][19] ) );
  DFFRX1 \register_reg[9][18]  ( .D(n382), .CK(clk), .RN(n2192), .Q(
        \register[9][18] ) );
  DFFRX1 \register_reg[9][17]  ( .D(n381), .CK(clk), .RN(n2192), .Q(
        \register[9][17] ) );
  DFFRX1 \register_reg[9][16]  ( .D(n380), .CK(clk), .RN(n2192), .Q(
        \register[9][16] ) );
  DFFRX1 \register_reg[9][15]  ( .D(n379), .CK(clk), .RN(n2192), .Q(
        \register[9][15] ) );
  DFFRX1 \register_reg[9][14]  ( .D(n378), .CK(clk), .RN(n2192), .Q(
        \register[9][14] ) );
  DFFRX1 \register_reg[9][13]  ( .D(n377), .CK(clk), .RN(n2192), .Q(
        \register[9][13] ) );
  DFFRX1 \register_reg[9][12]  ( .D(n376), .CK(clk), .RN(n2192), .Q(
        \register[9][12] ) );
  DFFRX1 \register_reg[9][11]  ( .D(n375), .CK(clk), .RN(n2192), .Q(
        \register[9][11] ) );
  DFFRX1 \register_reg[9][10]  ( .D(n374), .CK(clk), .RN(n2192), .Q(
        \register[9][10] ) );
  DFFRX1 \register_reg[9][9]  ( .D(n373), .CK(clk), .RN(n2192), .Q(
        \register[9][9] ) );
  DFFRX1 \register_reg[9][8]  ( .D(n372), .CK(clk), .RN(n2192), .Q(
        \register[9][8] ) );
  DFFRX1 \register_reg[9][7]  ( .D(n371), .CK(clk), .RN(n2191), .Q(
        \register[9][7] ) );
  DFFRX1 \register_reg[9][6]  ( .D(n370), .CK(clk), .RN(n2191), .Q(
        \register[9][6] ) );
  DFFRX1 \register_reg[9][5]  ( .D(n369), .CK(clk), .RN(n2191), .Q(
        \register[9][5] ) );
  DFFRX1 \register_reg[9][4]  ( .D(n368), .CK(clk), .RN(n2191), .Q(
        \register[9][4] ) );
  DFFRX1 \register_reg[9][3]  ( .D(n367), .CK(clk), .RN(n2191), .Q(
        \register[9][3] ) );
  DFFRX1 \register_reg[9][2]  ( .D(n366), .CK(clk), .RN(n2191), .Q(
        \register[9][2] ) );
  DFFRX1 \register_reg[9][1]  ( .D(n365), .CK(clk), .RN(n2191), .Q(
        \register[9][1] ) );
  DFFRX1 \register_reg[9][0]  ( .D(n364), .CK(clk), .RN(n2191), .Q(
        \register[9][0] ) );
  DFFRX1 \register_reg[5][31]  ( .D(n267), .CK(clk), .RN(n2199), .Q(
        \register[5][31] ) );
  DFFRX1 \register_reg[5][30]  ( .D(n266), .CK(clk), .RN(n2199), .Q(
        \register[5][30] ) );
  DFFRX1 \register_reg[5][29]  ( .D(n265), .CK(clk), .RN(n2199), .Q(
        \register[5][29] ) );
  DFFRX1 \register_reg[5][28]  ( .D(n264), .CK(clk), .RN(n2199), .Q(
        \register[5][28] ) );
  DFFRX1 \register_reg[5][27]  ( .D(n263), .CK(clk), .RN(n2198), .Q(
        \register[5][27] ) );
  DFFRX1 \register_reg[5][26]  ( .D(n262), .CK(clk), .RN(n2198), .Q(
        \register[5][26] ) );
  DFFRX1 \register_reg[5][25]  ( .D(n261), .CK(clk), .RN(n2198), .Q(
        \register[5][25] ) );
  DFFRX1 \register_reg[5][24]  ( .D(n260), .CK(clk), .RN(n2198), .Q(
        \register[5][24] ) );
  DFFRX1 \register_reg[5][23]  ( .D(n259), .CK(clk), .RN(n2198), .Q(
        \register[5][23] ) );
  DFFRX1 \register_reg[5][22]  ( .D(n258), .CK(clk), .RN(n2198), .Q(
        \register[5][22] ) );
  DFFRX1 \register_reg[5][21]  ( .D(n257), .CK(clk), .RN(n2198), .Q(
        \register[5][21] ) );
  DFFRX1 \register_reg[5][20]  ( .D(n256), .CK(clk), .RN(n2198), .Q(
        \register[5][20] ) );
  DFFRX1 \register_reg[5][19]  ( .D(n255), .CK(clk), .RN(n2198), .Q(
        \register[5][19] ) );
  DFFRX1 \register_reg[5][18]  ( .D(n254), .CK(clk), .RN(n2198), .Q(
        \register[5][18] ) );
  DFFRX1 \register_reg[5][17]  ( .D(n253), .CK(clk), .RN(n2198), .Q(
        \register[5][17] ) );
  DFFRX1 \register_reg[5][16]  ( .D(n252), .CK(clk), .RN(n2198), .Q(
        \register[5][16] ) );
  DFFRX1 \register_reg[5][15]  ( .D(n251), .CK(clk), .RN(n2197), .Q(
        \register[5][15] ) );
  DFFRX1 \register_reg[5][14]  ( .D(n250), .CK(clk), .RN(n2197), .Q(
        \register[5][14] ) );
  DFFRX1 \register_reg[5][13]  ( .D(n249), .CK(clk), .RN(n2197), .Q(
        \register[5][13] ) );
  DFFRX1 \register_reg[5][12]  ( .D(n248), .CK(clk), .RN(n2197), .Q(
        \register[5][12] ) );
  DFFRX1 \register_reg[5][11]  ( .D(n247), .CK(clk), .RN(n2197), .Q(
        \register[5][11] ) );
  DFFRX1 \register_reg[5][10]  ( .D(n246), .CK(clk), .RN(n2197), .Q(
        \register[5][10] ) );
  DFFRX1 \register_reg[5][9]  ( .D(n245), .CK(clk), .RN(n2197), .Q(
        \register[5][9] ) );
  DFFRX1 \register_reg[5][8]  ( .D(n244), .CK(clk), .RN(n2197), .Q(
        \register[5][8] ) );
  DFFRX1 \register_reg[5][7]  ( .D(n243), .CK(clk), .RN(n2197), .Q(
        \register[5][7] ) );
  DFFRX1 \register_reg[5][6]  ( .D(n242), .CK(clk), .RN(n2197), .Q(
        \register[5][6] ) );
  DFFRX1 \register_reg[5][5]  ( .D(n241), .CK(clk), .RN(n2197), .Q(
        \register[5][5] ) );
  DFFRX1 \register_reg[5][4]  ( .D(n240), .CK(clk), .RN(n2197), .Q(
        \register[5][4] ) );
  DFFRX1 \register_reg[5][3]  ( .D(n239), .CK(clk), .RN(n2181), .Q(
        \register[5][3] ) );
  DFFRX1 \register_reg[5][2]  ( .D(n238), .CK(clk), .RN(n2181), .Q(
        \register[5][2] ) );
  DFFRX1 \register_reg[5][1]  ( .D(n237), .CK(clk), .RN(n2181), .Q(
        \register[5][1] ) );
  DFFRX1 \register_reg[5][0]  ( .D(n236), .CK(clk), .RN(n2181), .Q(
        \register[5][0] ) );
  DFFRX1 \register_reg[28][31]  ( .D(n1003), .CK(clk), .RN(n2260), .Q(
        \register[28][31] ) );
  DFFRX1 \register_reg[28][30]  ( .D(n1002), .CK(clk), .RN(n2260), .Q(
        \register[28][30] ) );
  DFFRX1 \register_reg[28][29]  ( .D(n1001), .CK(clk), .RN(n2260), .Q(
        \register[28][29] ) );
  DFFRX1 \register_reg[28][28]  ( .D(n1000), .CK(clk), .RN(n2260), .Q(
        \register[28][28] ) );
  DFFRX1 \register_reg[28][27]  ( .D(n999), .CK(clk), .RN(n2260), .Q(
        \register[28][27] ) );
  DFFRX1 \register_reg[28][26]  ( .D(n998), .CK(clk), .RN(n2260), .Q(
        \register[28][26] ) );
  DFFRX1 \register_reg[28][25]  ( .D(n997), .CK(clk), .RN(n2260), .Q(
        \register[28][25] ) );
  DFFRX1 \register_reg[28][24]  ( .D(n996), .CK(clk), .RN(n2260), .Q(
        \register[28][24] ) );
  DFFRX1 \register_reg[28][23]  ( .D(n995), .CK(clk), .RN(n2258), .Q(
        \register[28][23] ) );
  DFFRX1 \register_reg[28][22]  ( .D(n994), .CK(clk), .RN(n2258), .Q(
        \register[28][22] ) );
  DFFRX1 \register_reg[28][21]  ( .D(n993), .CK(clk), .RN(n2258), .Q(
        \register[28][21] ) );
  DFFRX1 \register_reg[28][20]  ( .D(n992), .CK(clk), .RN(n2258), .Q(
        \register[28][20] ) );
  DFFRX1 \register_reg[28][19]  ( .D(n991), .CK(clk), .RN(n2259), .Q(
        \register[28][19] ) );
  DFFRX1 \register_reg[28][18]  ( .D(n990), .CK(clk), .RN(n2259), .Q(
        \register[28][18] ) );
  DFFRX1 \register_reg[28][17]  ( .D(n989), .CK(clk), .RN(n2259), .Q(
        \register[28][17] ) );
  DFFRX1 \register_reg[28][16]  ( .D(n988), .CK(clk), .RN(n2259), .Q(
        \register[28][16] ) );
  DFFRX1 \register_reg[28][15]  ( .D(n987), .CK(clk), .RN(n2259), .Q(
        \register[28][15] ) );
  DFFRX1 \register_reg[28][14]  ( .D(n986), .CK(clk), .RN(n2259), .Q(
        \register[28][14] ) );
  DFFRX1 \register_reg[28][13]  ( .D(n985), .CK(clk), .RN(n2259), .Q(
        \register[28][13] ) );
  DFFRX1 \register_reg[28][12]  ( .D(n984), .CK(clk), .RN(n2259), .Q(
        \register[28][12] ) );
  DFFRX1 \register_reg[28][11]  ( .D(n983), .CK(clk), .RN(n2257), .Q(
        \register[28][11] ) );
  DFFRX1 \register_reg[28][10]  ( .D(n982), .CK(clk), .RN(n2257), .Q(
        \register[28][10] ) );
  DFFRX1 \register_reg[28][9]  ( .D(n981), .CK(clk), .RN(n2257), .Q(
        \register[28][9] ) );
  DFFRX1 \register_reg[28][8]  ( .D(n980), .CK(clk), .RN(n2257), .Q(
        \register[28][8] ) );
  DFFRX1 \register_reg[28][7]  ( .D(n979), .CK(clk), .RN(n2258), .Q(
        \register[28][7] ) );
  DFFRX1 \register_reg[28][6]  ( .D(n978), .CK(clk), .RN(n2258), .Q(
        \register[28][6] ) );
  DFFRX1 \register_reg[28][5]  ( .D(n977), .CK(clk), .RN(n2258), .Q(
        \register[28][5] ) );
  DFFRX1 \register_reg[28][4]  ( .D(n976), .CK(clk), .RN(n2258), .Q(
        \register[28][4] ) );
  DFFRX1 \register_reg[28][3]  ( .D(n975), .CK(clk), .RN(n2258), .Q(
        \register[28][3] ) );
  DFFRX1 \register_reg[28][2]  ( .D(n974), .CK(clk), .RN(n2258), .Q(
        \register[28][2] ) );
  DFFRX1 \register_reg[28][1]  ( .D(n973), .CK(clk), .RN(n2258), .Q(
        \register[28][1] ) );
  DFFRX1 \register_reg[28][0]  ( .D(n972), .CK(clk), .RN(n2258), .Q(
        \register[28][0] ) );
  DFFRX1 \register_reg[24][31]  ( .D(n875), .CK(clk), .RN(n2241), .Q(
        \register[24][31] ) );
  DFFRX1 \register_reg[24][30]  ( .D(n874), .CK(clk), .RN(n2241), .Q(
        \register[24][30] ) );
  DFFRX1 \register_reg[24][29]  ( .D(n873), .CK(clk), .RN(n2241), .Q(
        \register[24][29] ) );
  DFFRX1 \register_reg[24][28]  ( .D(n872), .CK(clk), .RN(n2241), .Q(
        \register[24][28] ) );
  DFFRX1 \register_reg[24][27]  ( .D(n871), .CK(clk), .RN(n2241), .Q(
        \register[24][27] ) );
  DFFRX1 \register_reg[24][26]  ( .D(n870), .CK(clk), .RN(n2241), .Q(
        \register[24][26] ) );
  DFFRX1 \register_reg[24][25]  ( .D(n869), .CK(clk), .RN(n2241), .Q(
        \register[24][25] ) );
  DFFRX1 \register_reg[24][24]  ( .D(n868), .CK(clk), .RN(n2241), .Q(
        \register[24][24] ) );
  DFFRX1 \register_reg[24][23]  ( .D(n867), .CK(clk), .RN(n2241), .Q(
        \register[24][23] ) );
  DFFRX1 \register_reg[24][22]  ( .D(n866), .CK(clk), .RN(n2241), .Q(
        \register[24][22] ) );
  DFFRX1 \register_reg[24][21]  ( .D(n865), .CK(clk), .RN(n2241), .Q(
        \register[24][21] ) );
  DFFRX1 \register_reg[24][20]  ( .D(n864), .CK(clk), .RN(n2241), .Q(
        \register[24][20] ) );
  DFFRX1 \register_reg[24][19]  ( .D(n863), .CK(clk), .RN(n2248), .Q(
        \register[24][19] ) );
  DFFRX1 \register_reg[24][18]  ( .D(n862), .CK(clk), .RN(n2248), .Q(
        \register[24][18] ) );
  DFFRX1 \register_reg[24][17]  ( .D(n861), .CK(clk), .RN(n2248), .Q(
        \register[24][17] ) );
  DFFRX1 \register_reg[24][16]  ( .D(n860), .CK(clk), .RN(n2248), .Q(
        \register[24][16] ) );
  DFFRX1 \register_reg[24][15]  ( .D(n859), .CK(clk), .RN(n2248), .Q(
        \register[24][15] ) );
  DFFRX1 \register_reg[24][14]  ( .D(n858), .CK(clk), .RN(n2248), .Q(
        \register[24][14] ) );
  DFFRX1 \register_reg[24][13]  ( .D(n857), .CK(clk), .RN(n2248), .Q(
        \register[24][13] ) );
  DFFRX1 \register_reg[24][12]  ( .D(n856), .CK(clk), .RN(n2248), .Q(
        \register[24][12] ) );
  DFFRX1 \register_reg[24][11]  ( .D(n855), .CK(clk), .RN(n2248), .Q(
        \register[24][11] ) );
  DFFRX1 \register_reg[24][10]  ( .D(n854), .CK(clk), .RN(n2248), .Q(
        \register[24][10] ) );
  DFFRX1 \register_reg[24][9]  ( .D(n853), .CK(clk), .RN(n2248), .Q(
        \register[24][9] ) );
  DFFRX1 \register_reg[24][8]  ( .D(n852), .CK(clk), .RN(n2248), .Q(
        \register[24][8] ) );
  DFFRX1 \register_reg[24][7]  ( .D(n851), .CK(clk), .RN(n2247), .Q(
        \register[24][7] ) );
  DFFRX1 \register_reg[24][6]  ( .D(n850), .CK(clk), .RN(n2247), .Q(
        \register[24][6] ) );
  DFFRX1 \register_reg[24][5]  ( .D(n849), .CK(clk), .RN(n2247), .Q(
        \register[24][5] ) );
  DFFRX1 \register_reg[24][4]  ( .D(n848), .CK(clk), .RN(n2247), .Q(
        \register[24][4] ) );
  DFFRX1 \register_reg[24][3]  ( .D(n847), .CK(clk), .RN(n2247), .Q(
        \register[24][3] ) );
  DFFRX1 \register_reg[24][2]  ( .D(n846), .CK(clk), .RN(n2247), .Q(
        \register[24][2] ) );
  DFFRX1 \register_reg[24][1]  ( .D(n845), .CK(clk), .RN(n2247), .Q(
        \register[24][1] ) );
  DFFRX1 \register_reg[24][0]  ( .D(n844), .CK(clk), .RN(n2247), .Q(
        \register[24][0] ) );
  DFFRX1 \register_reg[20][31]  ( .D(n747), .CK(clk), .RN(n2231), .Q(
        \register[20][31] ) );
  DFFRX1 \register_reg[20][30]  ( .D(n746), .CK(clk), .RN(n2231), .Q(
        \register[20][30] ) );
  DFFRX1 \register_reg[20][29]  ( .D(n745), .CK(clk), .RN(n2231), .Q(
        \register[20][29] ) );
  DFFRX1 \register_reg[20][28]  ( .D(n744), .CK(clk), .RN(n2231), .Q(
        \register[20][28] ) );
  DFFRX1 \register_reg[20][27]  ( .D(n743), .CK(clk), .RN(n2230), .Q(
        \register[20][27] ) );
  DFFRX1 \register_reg[20][26]  ( .D(n742), .CK(clk), .RN(n2230), .Q(
        \register[20][26] ) );
  DFFRX1 \register_reg[20][25]  ( .D(n741), .CK(clk), .RN(n2230), .Q(
        \register[20][25] ) );
  DFFRX1 \register_reg[20][24]  ( .D(n740), .CK(clk), .RN(n2230), .Q(
        \register[20][24] ) );
  DFFRX1 \register_reg[20][23]  ( .D(n739), .CK(clk), .RN(n2230), .Q(
        \register[20][23] ) );
  DFFRX1 \register_reg[20][22]  ( .D(n738), .CK(clk), .RN(n2230), .Q(
        \register[20][22] ) );
  DFFRX1 \register_reg[20][21]  ( .D(n737), .CK(clk), .RN(n2230), .Q(
        \register[20][21] ) );
  DFFRX1 \register_reg[20][20]  ( .D(n736), .CK(clk), .RN(n2230), .Q(
        \register[20][20] ) );
  DFFRX1 \register_reg[20][19]  ( .D(n735), .CK(clk), .RN(n2230), .Q(
        \register[20][19] ) );
  DFFRX1 \register_reg[20][18]  ( .D(n734), .CK(clk), .RN(n2230), .Q(
        \register[20][18] ) );
  DFFRX1 \register_reg[20][17]  ( .D(n733), .CK(clk), .RN(n2230), .Q(
        \register[20][17] ) );
  DFFRX1 \register_reg[20][16]  ( .D(n732), .CK(clk), .RN(n2230), .Q(
        \register[20][16] ) );
  DFFRX1 \register_reg[20][15]  ( .D(n731), .CK(clk), .RN(n2229), .Q(
        \register[20][15] ) );
  DFFRX1 \register_reg[20][14]  ( .D(n730), .CK(clk), .RN(n2229), .Q(
        \register[20][14] ) );
  DFFRX1 \register_reg[20][13]  ( .D(n729), .CK(clk), .RN(n2229), .Q(
        \register[20][13] ) );
  DFFRX1 \register_reg[20][12]  ( .D(n728), .CK(clk), .RN(n2229), .Q(
        \register[20][12] ) );
  DFFRX1 \register_reg[20][11]  ( .D(n727), .CK(clk), .RN(n2229), .Q(
        \register[20][11] ) );
  DFFRX1 \register_reg[20][10]  ( .D(n726), .CK(clk), .RN(n2229), .Q(
        \register[20][10] ) );
  DFFRX1 \register_reg[20][9]  ( .D(n725), .CK(clk), .RN(n2229), .Q(
        \register[20][9] ) );
  DFFRX1 \register_reg[20][8]  ( .D(n724), .CK(clk), .RN(n2229), .Q(
        \register[20][8] ) );
  DFFRX1 \register_reg[20][7]  ( .D(n723), .CK(clk), .RN(n2229), .Q(
        \register[20][7] ) );
  DFFRX1 \register_reg[20][6]  ( .D(n722), .CK(clk), .RN(n2229), .Q(
        \register[20][6] ) );
  DFFRX1 \register_reg[20][5]  ( .D(n721), .CK(clk), .RN(n2229), .Q(
        \register[20][5] ) );
  DFFRX1 \register_reg[20][4]  ( .D(n720), .CK(clk), .RN(n2229), .Q(
        \register[20][4] ) );
  DFFRX1 \register_reg[20][3]  ( .D(n719), .CK(clk), .RN(n2236), .Q(
        \register[20][3] ) );
  DFFRX1 \register_reg[20][2]  ( .D(n718), .CK(clk), .RN(n2236), .Q(
        \register[20][2] ) );
  DFFRX1 \register_reg[20][1]  ( .D(n717), .CK(clk), .RN(n2236), .Q(
        \register[20][1] ) );
  DFFRX1 \register_reg[20][0]  ( .D(n716), .CK(clk), .RN(n2236), .Q(
        \register[20][0] ) );
  DFFRX1 \register_reg[16][31]  ( .D(n619), .CK(clk), .RN(n2220), .Q(
        \register[16][31] ) );
  DFFRX1 \register_reg[16][30]  ( .D(n618), .CK(clk), .RN(n2220), .Q(
        \register[16][30] ) );
  DFFRX1 \register_reg[16][29]  ( .D(n617), .CK(clk), .RN(n2220), .Q(
        \register[16][29] ) );
  DFFRX1 \register_reg[16][28]  ( .D(n616), .CK(clk), .RN(n2220), .Q(
        \register[16][28] ) );
  DFFRX1 \register_reg[16][27]  ( .D(n615), .CK(clk), .RN(n2220), .Q(
        \register[16][27] ) );
  DFFRX1 \register_reg[16][26]  ( .D(n614), .CK(clk), .RN(n2220), .Q(
        \register[16][26] ) );
  DFFRX1 \register_reg[16][25]  ( .D(n613), .CK(clk), .RN(n2220), .Q(
        \register[16][25] ) );
  DFFRX1 \register_reg[16][24]  ( .D(n612), .CK(clk), .RN(n2220), .Q(
        \register[16][24] ) );
  DFFRX1 \register_reg[16][23]  ( .D(n611), .CK(clk), .RN(n2219), .Q(
        \register[16][23] ) );
  DFFRX1 \register_reg[16][22]  ( .D(n610), .CK(clk), .RN(n2219), .Q(
        \register[16][22] ) );
  DFFRX1 \register_reg[16][21]  ( .D(n609), .CK(clk), .RN(n2219), .Q(
        \register[16][21] ) );
  DFFRX1 \register_reg[16][20]  ( .D(n608), .CK(clk), .RN(n2219), .Q(
        \register[16][20] ) );
  DFFRX1 \register_reg[16][19]  ( .D(n607), .CK(clk), .RN(n2219), .Q(
        \register[16][19] ) );
  DFFRX1 \register_reg[16][18]  ( .D(n606), .CK(clk), .RN(n2219), .Q(
        \register[16][18] ) );
  DFFRX1 \register_reg[16][17]  ( .D(n605), .CK(clk), .RN(n2219), .Q(
        \register[16][17] ) );
  DFFRX1 \register_reg[16][16]  ( .D(n604), .CK(clk), .RN(n2219), .Q(
        \register[16][16] ) );
  DFFRX1 \register_reg[16][15]  ( .D(n603), .CK(clk), .RN(n2219), .Q(
        \register[16][15] ) );
  DFFRX1 \register_reg[16][14]  ( .D(n602), .CK(clk), .RN(n2219), .Q(
        \register[16][14] ) );
  DFFRX1 \register_reg[16][13]  ( .D(n601), .CK(clk), .RN(n2219), .Q(
        \register[16][13] ) );
  DFFRX1 \register_reg[16][12]  ( .D(n600), .CK(clk), .RN(n2219), .Q(
        \register[16][12] ) );
  DFFRX1 \register_reg[16][11]  ( .D(n599), .CK(clk), .RN(n2218), .Q(
        \register[16][11] ) );
  DFFRX1 \register_reg[16][10]  ( .D(n598), .CK(clk), .RN(n2218), .Q(
        \register[16][10] ) );
  DFFRX1 \register_reg[16][9]  ( .D(n597), .CK(clk), .RN(n2218), .Q(
        \register[16][9] ) );
  DFFRX1 \register_reg[16][8]  ( .D(n596), .CK(clk), .RN(n2218), .Q(
        \register[16][8] ) );
  DFFRX1 \register_reg[16][7]  ( .D(n595), .CK(clk), .RN(n2218), .Q(
        \register[16][7] ) );
  DFFRX1 \register_reg[16][6]  ( .D(n594), .CK(clk), .RN(n2218), .Q(
        \register[16][6] ) );
  DFFRX1 \register_reg[16][5]  ( .D(n593), .CK(clk), .RN(n2218), .Q(
        \register[16][5] ) );
  DFFRX1 \register_reg[16][4]  ( .D(n592), .CK(clk), .RN(n2218), .Q(
        \register[16][4] ) );
  DFFRX1 \register_reg[16][3]  ( .D(n591), .CK(clk), .RN(n2218), .Q(
        \register[16][3] ) );
  DFFRX1 \register_reg[16][2]  ( .D(n590), .CK(clk), .RN(n2218), .Q(
        \register[16][2] ) );
  DFFRX1 \register_reg[16][1]  ( .D(n589), .CK(clk), .RN(n2218), .Q(
        \register[16][1] ) );
  DFFRX1 \register_reg[16][0]  ( .D(n588), .CK(clk), .RN(n2218), .Q(
        \register[16][0] ) );
  DFFRX1 \register_reg[12][31]  ( .D(n491), .CK(clk), .RN(n2201), .Q(
        \register[12][31] ) );
  DFFRX1 \register_reg[12][30]  ( .D(n490), .CK(clk), .RN(n2201), .Q(
        \register[12][30] ) );
  DFFRX1 \register_reg[12][29]  ( .D(n489), .CK(clk), .RN(n2201), .Q(
        \register[12][29] ) );
  DFFRX1 \register_reg[12][28]  ( .D(n488), .CK(clk), .RN(n2201), .Q(
        \register[12][28] ) );
  DFFRX1 \register_reg[12][27]  ( .D(n487), .CK(clk), .RN(n2201), .Q(
        \register[12][27] ) );
  DFFRX1 \register_reg[12][26]  ( .D(n486), .CK(clk), .RN(n2201), .Q(
        \register[12][26] ) );
  DFFRX1 \register_reg[12][25]  ( .D(n485), .CK(clk), .RN(n2201), .Q(
        \register[12][25] ) );
  DFFRX1 \register_reg[12][24]  ( .D(n484), .CK(clk), .RN(n2201), .Q(
        \register[12][24] ) );
  DFFRX1 \register_reg[12][23]  ( .D(n483), .CK(clk), .RN(n2201), .Q(
        \register[12][23] ) );
  DFFRX1 \register_reg[12][22]  ( .D(n482), .CK(clk), .RN(n2201), .Q(
        \register[12][22] ) );
  DFFRX1 \register_reg[12][21]  ( .D(n481), .CK(clk), .RN(n2201), .Q(
        \register[12][21] ) );
  DFFRX1 \register_reg[12][20]  ( .D(n480), .CK(clk), .RN(n2201), .Q(
        \register[12][20] ) );
  DFFRX1 \register_reg[12][19]  ( .D(n479), .CK(clk), .RN(n2208), .Q(
        \register[12][19] ) );
  DFFRX1 \register_reg[12][18]  ( .D(n478), .CK(clk), .RN(n2208), .Q(
        \register[12][18] ) );
  DFFRX1 \register_reg[12][17]  ( .D(n477), .CK(clk), .RN(n2208), .Q(
        \register[12][17] ) );
  DFFRX1 \register_reg[12][16]  ( .D(n476), .CK(clk), .RN(n2208), .Q(
        \register[12][16] ) );
  DFFRX1 \register_reg[12][15]  ( .D(n475), .CK(clk), .RN(n2208), .Q(
        \register[12][15] ) );
  DFFRX1 \register_reg[12][14]  ( .D(n474), .CK(clk), .RN(n2208), .Q(
        \register[12][14] ) );
  DFFRX1 \register_reg[12][13]  ( .D(n473), .CK(clk), .RN(n2208), .Q(
        \register[12][13] ) );
  DFFRX1 \register_reg[12][12]  ( .D(n472), .CK(clk), .RN(n2208), .Q(
        \register[12][12] ) );
  DFFRX1 \register_reg[12][11]  ( .D(n471), .CK(clk), .RN(n2208), .Q(
        \register[12][11] ) );
  DFFRX1 \register_reg[12][10]  ( .D(n470), .CK(clk), .RN(n2208), .Q(
        \register[12][10] ) );
  DFFRX1 \register_reg[12][9]  ( .D(n469), .CK(clk), .RN(n2208), .Q(
        \register[12][9] ) );
  DFFRX1 \register_reg[12][8]  ( .D(n468), .CK(clk), .RN(n2208), .Q(
        \register[12][8] ) );
  DFFRX1 \register_reg[12][7]  ( .D(n467), .CK(clk), .RN(n2207), .Q(
        \register[12][7] ) );
  DFFRX1 \register_reg[12][6]  ( .D(n466), .CK(clk), .RN(n2207), .Q(
        \register[12][6] ) );
  DFFRX1 \register_reg[12][5]  ( .D(n465), .CK(clk), .RN(n2207), .Q(
        \register[12][5] ) );
  DFFRX1 \register_reg[12][4]  ( .D(n464), .CK(clk), .RN(n2207), .Q(
        \register[12][4] ) );
  DFFRX1 \register_reg[12][3]  ( .D(n463), .CK(clk), .RN(n2207), .Q(
        \register[12][3] ) );
  DFFRX1 \register_reg[12][2]  ( .D(n462), .CK(clk), .RN(n2207), .Q(
        \register[12][2] ) );
  DFFRX1 \register_reg[12][1]  ( .D(n461), .CK(clk), .RN(n2207), .Q(
        \register[12][1] ) );
  DFFRX1 \register_reg[12][0]  ( .D(n460), .CK(clk), .RN(n2207), .Q(
        \register[12][0] ) );
  DFFRX1 \register_reg[8][31]  ( .D(n363), .CK(clk), .RN(n2191), .Q(
        \register[8][31] ) );
  DFFRX1 \register_reg[8][30]  ( .D(n362), .CK(clk), .RN(n2191), .Q(
        \register[8][30] ) );
  DFFRX1 \register_reg[8][29]  ( .D(n361), .CK(clk), .RN(n2191), .Q(
        \register[8][29] ) );
  DFFRX1 \register_reg[8][28]  ( .D(n360), .CK(clk), .RN(n2191), .Q(
        \register[8][28] ) );
  DFFRX1 \register_reg[8][27]  ( .D(n359), .CK(clk), .RN(n2190), .Q(
        \register[8][27] ) );
  DFFRX1 \register_reg[8][26]  ( .D(n358), .CK(clk), .RN(n2190), .Q(
        \register[8][26] ) );
  DFFRX1 \register_reg[8][25]  ( .D(n357), .CK(clk), .RN(n2190), .Q(
        \register[8][25] ) );
  DFFRX1 \register_reg[8][24]  ( .D(n356), .CK(clk), .RN(n2190), .Q(
        \register[8][24] ) );
  DFFRX1 \register_reg[8][23]  ( .D(n355), .CK(clk), .RN(n2190), .Q(
        \register[8][23] ) );
  DFFRX1 \register_reg[8][22]  ( .D(n354), .CK(clk), .RN(n2190), .Q(
        \register[8][22] ) );
  DFFRX1 \register_reg[8][21]  ( .D(n353), .CK(clk), .RN(n2190), .Q(
        \register[8][21] ) );
  DFFRX1 \register_reg[8][20]  ( .D(n352), .CK(clk), .RN(n2190), .Q(
        \register[8][20] ) );
  DFFRX1 \register_reg[8][19]  ( .D(n351), .CK(clk), .RN(n2190), .Q(
        \register[8][19] ) );
  DFFRX1 \register_reg[8][18]  ( .D(n350), .CK(clk), .RN(n2190), .Q(
        \register[8][18] ) );
  DFFRX1 \register_reg[8][17]  ( .D(n349), .CK(clk), .RN(n2190), .Q(
        \register[8][17] ) );
  DFFRX1 \register_reg[8][16]  ( .D(n348), .CK(clk), .RN(n2190), .Q(
        \register[8][16] ) );
  DFFRX1 \register_reg[8][15]  ( .D(n347), .CK(clk), .RN(n2189), .Q(
        \register[8][15] ) );
  DFFRX1 \register_reg[8][14]  ( .D(n346), .CK(clk), .RN(n2189), .Q(
        \register[8][14] ) );
  DFFRX1 \register_reg[8][13]  ( .D(n345), .CK(clk), .RN(n2189), .Q(
        \register[8][13] ) );
  DFFRX1 \register_reg[8][12]  ( .D(n344), .CK(clk), .RN(n2189), .Q(
        \register[8][12] ) );
  DFFRX1 \register_reg[8][11]  ( .D(n343), .CK(clk), .RN(n2189), .Q(
        \register[8][11] ) );
  DFFRX1 \register_reg[8][10]  ( .D(n342), .CK(clk), .RN(n2189), .Q(
        \register[8][10] ) );
  DFFRX1 \register_reg[8][9]  ( .D(n341), .CK(clk), .RN(n2189), .Q(
        \register[8][9] ) );
  DFFRX1 \register_reg[8][8]  ( .D(n340), .CK(clk), .RN(n2189), .Q(
        \register[8][8] ) );
  DFFRX1 \register_reg[8][7]  ( .D(n339), .CK(clk), .RN(n2189), .Q(
        \register[8][7] ) );
  DFFRX1 \register_reg[8][6]  ( .D(n338), .CK(clk), .RN(n2189), .Q(
        \register[8][6] ) );
  DFFRX1 \register_reg[8][5]  ( .D(n337), .CK(clk), .RN(n2189), .Q(
        \register[8][5] ) );
  DFFRX1 \register_reg[8][4]  ( .D(n336), .CK(clk), .RN(n2189), .Q(
        \register[8][4] ) );
  DFFRX1 \register_reg[8][3]  ( .D(n335), .CK(clk), .RN(n2196), .Q(
        \register[8][3] ) );
  DFFRX1 \register_reg[8][2]  ( .D(n334), .CK(clk), .RN(n2196), .Q(
        \register[8][2] ) );
  DFFRX1 \register_reg[8][1]  ( .D(n333), .CK(clk), .RN(n2196), .Q(
        \register[8][1] ) );
  DFFRX1 \register_reg[8][0]  ( .D(n332), .CK(clk), .RN(n2196), .Q(
        \register[8][0] ) );
  DFFRX1 \register_reg[4][31]  ( .D(n235), .CK(clk), .RN(n2181), .Q(
        \register[4][31] ) );
  DFFRX1 \register_reg[4][30]  ( .D(n234), .CK(clk), .RN(n2181), .Q(
        \register[4][30] ) );
  DFFRX1 \register_reg[4][29]  ( .D(n233), .CK(clk), .RN(n2181), .Q(
        \register[4][29] ) );
  DFFRX1 \register_reg[4][28]  ( .D(n232), .CK(clk), .RN(n2181), .Q(
        \register[4][28] ) );
  DFFRX1 \register_reg[4][27]  ( .D(n231), .CK(clk), .RN(n2181), .Q(
        \register[4][27] ) );
  DFFRX1 \register_reg[4][26]  ( .D(n230), .CK(clk), .RN(n2181), .Q(
        \register[4][26] ) );
  DFFRX1 \register_reg[4][25]  ( .D(n229), .CK(clk), .RN(n2181), .Q(
        \register[4][25] ) );
  DFFRX1 \register_reg[4][24]  ( .D(n228), .CK(clk), .RN(n2181), .Q(
        \register[4][24] ) );
  DFFRX1 \register_reg[4][23]  ( .D(n227), .CK(clk), .RN(n2180), .Q(
        \register[4][23] ) );
  DFFRX1 \register_reg[4][22]  ( .D(n226), .CK(clk), .RN(n2180), .Q(
        \register[4][22] ) );
  DFFRX1 \register_reg[4][21]  ( .D(n225), .CK(clk), .RN(n2180), .Q(
        \register[4][21] ) );
  DFFRX1 \register_reg[4][20]  ( .D(n224), .CK(clk), .RN(n2180), .Q(
        \register[4][20] ) );
  DFFRX1 \register_reg[4][19]  ( .D(n223), .CK(clk), .RN(n2180), .Q(
        \register[4][19] ) );
  DFFRX1 \register_reg[4][18]  ( .D(n222), .CK(clk), .RN(n2180), .Q(
        \register[4][18] ) );
  DFFRX1 \register_reg[4][17]  ( .D(n221), .CK(clk), .RN(n2180), .Q(
        \register[4][17] ) );
  DFFRX1 \register_reg[4][16]  ( .D(n220), .CK(clk), .RN(n2180), .Q(
        \register[4][16] ) );
  DFFRX1 \register_reg[4][15]  ( .D(n219), .CK(clk), .RN(n2180), .Q(
        \register[4][15] ) );
  DFFRX1 \register_reg[4][14]  ( .D(n218), .CK(clk), .RN(n2180), .Q(
        \register[4][14] ) );
  DFFRX1 \register_reg[4][13]  ( .D(n217), .CK(clk), .RN(n2180), .Q(
        \register[4][13] ) );
  DFFRX1 \register_reg[4][12]  ( .D(n216), .CK(clk), .RN(n2180), .Q(
        \register[4][12] ) );
  DFFRX1 \register_reg[4][11]  ( .D(n215), .CK(clk), .RN(n2179), .Q(
        \register[4][11] ) );
  DFFRX1 \register_reg[4][10]  ( .D(n214), .CK(clk), .RN(n2179), .Q(
        \register[4][10] ) );
  DFFRX1 \register_reg[4][9]  ( .D(n213), .CK(clk), .RN(n2179), .Q(
        \register[4][9] ) );
  DFFRX1 \register_reg[4][8]  ( .D(n212), .CK(clk), .RN(n2179), .Q(
        \register[4][8] ) );
  DFFRX1 \register_reg[4][7]  ( .D(n211), .CK(clk), .RN(n2179), .Q(
        \register[4][7] ) );
  DFFRX1 \register_reg[4][6]  ( .D(n210), .CK(clk), .RN(n2179), .Q(
        \register[4][6] ) );
  DFFRX1 \register_reg[4][5]  ( .D(n209), .CK(clk), .RN(n2179), .Q(
        \register[4][5] ) );
  DFFRX1 \register_reg[4][4]  ( .D(n208), .CK(clk), .RN(n2179), .Q(
        \register[4][4] ) );
  DFFRX1 \register_reg[4][3]  ( .D(n207), .CK(clk), .RN(n2179), .Q(
        \register[4][3] ) );
  DFFRX1 \register_reg[4][2]  ( .D(n206), .CK(clk), .RN(n2179), .Q(
        \register[4][2] ) );
  DFFRX1 \register_reg[4][1]  ( .D(n205), .CK(clk), .RN(n2179), .Q(
        \register[4][1] ) );
  DFFRX1 \register_reg[4][0]  ( .D(n204), .CK(clk), .RN(n2179), .Q(
        \register[4][0] ) );
  DFFRX1 \register_reg[30][31]  ( .D(n1067), .CK(clk), .RN(n2249), .Q(
        \register[30][31] ) );
  DFFRX1 \register_reg[30][30]  ( .D(n1066), .CK(clk), .RN(n2249), .Q(
        \register[30][30] ) );
  DFFRX1 \register_reg[30][29]  ( .D(n1065), .CK(clk), .RN(n2249), .Q(
        \register[30][29] ) );
  DFFRX1 \register_reg[30][28]  ( .D(n1064), .CK(clk), .RN(n2249), .Q(
        \register[30][28] ) );
  DFFRX1 \register_reg[30][27]  ( .D(n1063), .CK(clk), .RN(n2249), .Q(
        \register[30][27] ) );
  DFFRX1 \register_reg[30][26]  ( .D(n1062), .CK(clk), .RN(n2249), .Q(
        \register[30][26] ) );
  DFFRX1 \register_reg[30][25]  ( .D(n1061), .CK(clk), .RN(n2249), .Q(
        \register[30][25] ) );
  DFFRX1 \register_reg[30][24]  ( .D(n1060), .CK(clk), .RN(n2249), .Q(
        \register[30][24] ) );
  DFFRX1 \register_reg[30][23]  ( .D(n1059), .CK(clk), .RN(n2249), .Q(
        \register[30][23] ) );
  DFFRX1 \register_reg[30][22]  ( .D(n1058), .CK(clk), .RN(n2249), .Q(
        \register[30][22] ) );
  DFFRX1 \register_reg[30][21]  ( .D(n1057), .CK(clk), .RN(n2249), .Q(
        \register[30][21] ) );
  DFFRX1 \register_reg[30][20]  ( .D(n1056), .CK(clk), .RN(n2249), .Q(
        \register[30][20] ) );
  DFFRX1 \register_reg[30][19]  ( .D(n1055), .CK(clk), .RN(n2255), .Q(
        \register[30][19] ) );
  DFFRX1 \register_reg[30][18]  ( .D(n1054), .CK(clk), .RN(n2255), .Q(
        \register[30][18] ) );
  DFFRX1 \register_reg[30][17]  ( .D(n1053), .CK(clk), .RN(n2255), .Q(
        \register[30][17] ) );
  DFFRX1 \register_reg[30][16]  ( .D(n1052), .CK(clk), .RN(n2255), .Q(
        \register[30][16] ) );
  DFFRX1 \register_reg[30][15]  ( .D(n1051), .CK(clk), .RN(n2256), .Q(
        \register[30][15] ) );
  DFFRX1 \register_reg[30][14]  ( .D(n1050), .CK(clk), .RN(n2256), .Q(
        \register[30][14] ) );
  DFFRX1 \register_reg[30][13]  ( .D(n1049), .CK(clk), .RN(n2256), .Q(
        \register[30][13] ) );
  DFFRX1 \register_reg[30][12]  ( .D(n1048), .CK(clk), .RN(n2256), .Q(
        \register[30][12] ) );
  DFFRX1 \register_reg[30][11]  ( .D(n1047), .CK(clk), .RN(n2256), .Q(
        \register[30][11] ) );
  DFFRX1 \register_reg[30][10]  ( .D(n1046), .CK(clk), .RN(n2256), .Q(
        \register[30][10] ) );
  DFFRX1 \register_reg[30][9]  ( .D(n1045), .CK(clk), .RN(n2256), .Q(
        \register[30][9] ) );
  DFFRX1 \register_reg[30][8]  ( .D(n1044), .CK(clk), .RN(n2256), .Q(
        \register[30][8] ) );
  DFFRX1 \register_reg[30][7]  ( .D(n1043), .CK(clk), .RN(n2254), .Q(
        \register[30][7] ) );
  DFFRX1 \register_reg[30][6]  ( .D(n1042), .CK(clk), .RN(n2254), .Q(
        \register[30][6] ) );
  DFFRX1 \register_reg[30][5]  ( .D(n1041), .CK(clk), .RN(n2254), .Q(
        \register[30][5] ) );
  DFFRX1 \register_reg[30][4]  ( .D(n1040), .CK(clk), .RN(n2254), .Q(
        \register[30][4] ) );
  DFFRX1 \register_reg[30][3]  ( .D(n1039), .CK(clk), .RN(n2255), .Q(
        \register[30][3] ) );
  DFFRX1 \register_reg[30][2]  ( .D(n1038), .CK(clk), .RN(n2255), .Q(
        \register[30][2] ) );
  DFFRX1 \register_reg[30][1]  ( .D(n1037), .CK(clk), .RN(n2255), .Q(
        \register[30][1] ) );
  DFFRX1 \register_reg[30][0]  ( .D(n1036), .CK(clk), .RN(n2255), .Q(
        \register[30][0] ) );
  DFFRX1 \register_reg[26][31]  ( .D(n939), .CK(clk), .RN(n2239), .Q(
        \register[26][31] ) );
  DFFRX1 \register_reg[26][30]  ( .D(n938), .CK(clk), .RN(n2239), .Q(
        \register[26][30] ) );
  DFFRX1 \register_reg[26][29]  ( .D(n937), .CK(clk), .RN(n2239), .Q(
        \register[26][29] ) );
  DFFRX1 \register_reg[26][28]  ( .D(n936), .CK(clk), .RN(n2239), .Q(
        \register[26][28] ) );
  DFFRX1 \register_reg[26][27]  ( .D(n935), .CK(clk), .RN(n2238), .Q(
        \register[26][27] ) );
  DFFRX1 \register_reg[26][26]  ( .D(n934), .CK(clk), .RN(n2238), .Q(
        \register[26][26] ) );
  DFFRX1 \register_reg[26][25]  ( .D(n933), .CK(clk), .RN(n2238), .Q(
        \register[26][25] ) );
  DFFRX1 \register_reg[26][24]  ( .D(n932), .CK(clk), .RN(n2238), .Q(
        \register[26][24] ) );
  DFFRX1 \register_reg[26][23]  ( .D(n931), .CK(clk), .RN(n2238), .Q(
        \register[26][23] ) );
  DFFRX1 \register_reg[26][22]  ( .D(n930), .CK(clk), .RN(n2238), .Q(
        \register[26][22] ) );
  DFFRX1 \register_reg[26][21]  ( .D(n929), .CK(clk), .RN(n2238), .Q(
        \register[26][21] ) );
  DFFRX1 \register_reg[26][20]  ( .D(n928), .CK(clk), .RN(n2238), .Q(
        \register[26][20] ) );
  DFFRX1 \register_reg[26][19]  ( .D(n927), .CK(clk), .RN(n2238), .Q(
        \register[26][19] ) );
  DFFRX1 \register_reg[26][18]  ( .D(n926), .CK(clk), .RN(n2238), .Q(
        \register[26][18] ) );
  DFFRX1 \register_reg[26][17]  ( .D(n925), .CK(clk), .RN(n2238), .Q(
        \register[26][17] ) );
  DFFRX1 \register_reg[26][16]  ( .D(n924), .CK(clk), .RN(n2238), .Q(
        \register[26][16] ) );
  DFFRX1 \register_reg[26][15]  ( .D(n923), .CK(clk), .RN(n2237), .Q(
        \register[26][15] ) );
  DFFRX1 \register_reg[26][14]  ( .D(n922), .CK(clk), .RN(n2237), .Q(
        \register[26][14] ) );
  DFFRX1 \register_reg[26][13]  ( .D(n921), .CK(clk), .RN(n2237), .Q(
        \register[26][13] ) );
  DFFRX1 \register_reg[26][12]  ( .D(n920), .CK(clk), .RN(n2237), .Q(
        \register[26][12] ) );
  DFFRX1 \register_reg[26][11]  ( .D(n919), .CK(clk), .RN(n2237), .Q(
        \register[26][11] ) );
  DFFRX1 \register_reg[26][10]  ( .D(n918), .CK(clk), .RN(n2237), .Q(
        \register[26][10] ) );
  DFFRX1 \register_reg[26][9]  ( .D(n917), .CK(clk), .RN(n2237), .Q(
        \register[26][9] ) );
  DFFRX1 \register_reg[26][8]  ( .D(n916), .CK(clk), .RN(n2237), .Q(
        \register[26][8] ) );
  DFFRX1 \register_reg[26][7]  ( .D(n915), .CK(clk), .RN(n2237), .Q(
        \register[26][7] ) );
  DFFRX1 \register_reg[26][6]  ( .D(n914), .CK(clk), .RN(n2237), .Q(
        \register[26][6] ) );
  DFFRX1 \register_reg[26][5]  ( .D(n913), .CK(clk), .RN(n2237), .Q(
        \register[26][5] ) );
  DFFRX1 \register_reg[26][4]  ( .D(n912), .CK(clk), .RN(n2237), .Q(
        \register[26][4] ) );
  DFFRX1 \register_reg[26][3]  ( .D(n911), .CK(clk), .RN(n2244), .Q(
        \register[26][3] ) );
  DFFRX1 \register_reg[26][2]  ( .D(n910), .CK(clk), .RN(n2244), .Q(
        \register[26][2] ) );
  DFFRX1 \register_reg[26][1]  ( .D(n909), .CK(clk), .RN(n2244), .Q(
        \register[26][1] ) );
  DFFRX1 \register_reg[26][0]  ( .D(n908), .CK(clk), .RN(n2244), .Q(
        \register[26][0] ) );
  DFFRX1 \register_reg[22][31]  ( .D(n811), .CK(clk), .RN(n2228), .Q(
        \register[22][31] ) );
  DFFRX1 \register_reg[22][30]  ( .D(n810), .CK(clk), .RN(n2228), .Q(
        \register[22][30] ) );
  DFFRX1 \register_reg[22][29]  ( .D(n809), .CK(clk), .RN(n2228), .Q(
        \register[22][29] ) );
  DFFRX1 \register_reg[22][28]  ( .D(n808), .CK(clk), .RN(n2228), .Q(
        \register[22][28] ) );
  DFFRX1 \register_reg[22][27]  ( .D(n807), .CK(clk), .RN(n2228), .Q(
        \register[22][27] ) );
  DFFRX1 \register_reg[22][26]  ( .D(n806), .CK(clk), .RN(n2228), .Q(
        \register[22][26] ) );
  DFFRX1 \register_reg[22][25]  ( .D(n805), .CK(clk), .RN(n2228), .Q(
        \register[22][25] ) );
  DFFRX1 \register_reg[22][24]  ( .D(n804), .CK(clk), .RN(n2228), .Q(
        \register[22][24] ) );
  DFFRX1 \register_reg[22][23]  ( .D(n803), .CK(clk), .RN(n2227), .Q(
        \register[22][23] ) );
  DFFRX1 \register_reg[22][22]  ( .D(n802), .CK(clk), .RN(n2227), .Q(
        \register[22][22] ) );
  DFFRX1 \register_reg[22][21]  ( .D(n801), .CK(clk), .RN(n2227), .Q(
        \register[22][21] ) );
  DFFRX1 \register_reg[22][20]  ( .D(n800), .CK(clk), .RN(n2227), .Q(
        \register[22][20] ) );
  DFFRX1 \register_reg[22][19]  ( .D(n799), .CK(clk), .RN(n2227), .Q(
        \register[22][19] ) );
  DFFRX1 \register_reg[22][18]  ( .D(n798), .CK(clk), .RN(n2227), .Q(
        \register[22][18] ) );
  DFFRX1 \register_reg[22][17]  ( .D(n797), .CK(clk), .RN(n2227), .Q(
        \register[22][17] ) );
  DFFRX1 \register_reg[22][16]  ( .D(n796), .CK(clk), .RN(n2227), .Q(
        \register[22][16] ) );
  DFFRX1 \register_reg[22][15]  ( .D(n795), .CK(clk), .RN(n2227), .Q(
        \register[22][15] ) );
  DFFRX1 \register_reg[22][14]  ( .D(n794), .CK(clk), .RN(n2227), .Q(
        \register[22][14] ) );
  DFFRX1 \register_reg[22][13]  ( .D(n793), .CK(clk), .RN(n2227), .Q(
        \register[22][13] ) );
  DFFRX1 \register_reg[22][12]  ( .D(n792), .CK(clk), .RN(n2227), .Q(
        \register[22][12] ) );
  DFFRX1 \register_reg[22][11]  ( .D(n791), .CK(clk), .RN(n2226), .Q(
        \register[22][11] ) );
  DFFRX1 \register_reg[22][10]  ( .D(n790), .CK(clk), .RN(n2226), .Q(
        \register[22][10] ) );
  DFFRX1 \register_reg[22][9]  ( .D(n789), .CK(clk), .RN(n2226), .Q(
        \register[22][9] ) );
  DFFRX1 \register_reg[22][8]  ( .D(n788), .CK(clk), .RN(n2226), .Q(
        \register[22][8] ) );
  DFFRX1 \register_reg[22][7]  ( .D(n787), .CK(clk), .RN(n2226), .Q(
        \register[22][7] ) );
  DFFRX1 \register_reg[22][6]  ( .D(n786), .CK(clk), .RN(n2226), .Q(
        \register[22][6] ) );
  DFFRX1 \register_reg[22][5]  ( .D(n785), .CK(clk), .RN(n2226), .Q(
        \register[22][5] ) );
  DFFRX1 \register_reg[22][4]  ( .D(n784), .CK(clk), .RN(n2226), .Q(
        \register[22][4] ) );
  DFFRX1 \register_reg[22][3]  ( .D(n783), .CK(clk), .RN(n2226), .Q(
        \register[22][3] ) );
  DFFRX1 \register_reg[22][2]  ( .D(n782), .CK(clk), .RN(n2226), .Q(
        \register[22][2] ) );
  DFFRX1 \register_reg[22][1]  ( .D(n781), .CK(clk), .RN(n2226), .Q(
        \register[22][1] ) );
  DFFRX1 \register_reg[22][0]  ( .D(n780), .CK(clk), .RN(n2226), .Q(
        \register[22][0] ) );
  DFFRX1 \register_reg[18][31]  ( .D(n683), .CK(clk), .RN(n2233), .Q(
        \register[18][31] ) );
  DFFRX1 \register_reg[18][30]  ( .D(n682), .CK(clk), .RN(n2233), .Q(
        \register[18][30] ) );
  DFFRX1 \register_reg[18][29]  ( .D(n681), .CK(clk), .RN(n2233), .Q(
        \register[18][29] ) );
  DFFRX1 \register_reg[18][28]  ( .D(n680), .CK(clk), .RN(n2233), .Q(
        \register[18][28] ) );
  DFFRX1 \register_reg[18][27]  ( .D(n679), .CK(clk), .RN(n2233), .Q(
        \register[18][27] ) );
  DFFRX1 \register_reg[18][26]  ( .D(n678), .CK(clk), .RN(n2233), .Q(
        \register[18][26] ) );
  DFFRX1 \register_reg[18][25]  ( .D(n677), .CK(clk), .RN(n2233), .Q(
        \register[18][25] ) );
  DFFRX1 \register_reg[18][24]  ( .D(n676), .CK(clk), .RN(n2233), .Q(
        \register[18][24] ) );
  DFFRX1 \register_reg[18][23]  ( .D(n675), .CK(clk), .RN(n2233), .Q(
        \register[18][23] ) );
  DFFRX1 \register_reg[18][22]  ( .D(n674), .CK(clk), .RN(n2233), .Q(
        \register[18][22] ) );
  DFFRX1 \register_reg[18][21]  ( .D(n673), .CK(clk), .RN(n2233), .Q(
        \register[18][21] ) );
  DFFRX1 \register_reg[18][20]  ( .D(n672), .CK(clk), .RN(n2233), .Q(
        \register[18][20] ) );
  DFFRX1 \register_reg[18][19]  ( .D(n671), .CK(clk), .RN(n2216), .Q(
        \register[18][19] ) );
  DFFRX1 \register_reg[18][18]  ( .D(n670), .CK(clk), .RN(n2216), .Q(
        \register[18][18] ) );
  DFFRX1 \register_reg[18][17]  ( .D(n669), .CK(clk), .RN(n2216), .Q(
        \register[18][17] ) );
  DFFRX1 \register_reg[18][16]  ( .D(n668), .CK(clk), .RN(n2216), .Q(
        \register[18][16] ) );
  DFFRX1 \register_reg[18][15]  ( .D(n667), .CK(clk), .RN(n2216), .Q(
        \register[18][15] ) );
  DFFRX1 \register_reg[18][14]  ( .D(n666), .CK(clk), .RN(n2216), .Q(
        \register[18][14] ) );
  DFFRX1 \register_reg[18][13]  ( .D(n665), .CK(clk), .RN(n2216), .Q(
        \register[18][13] ) );
  DFFRX1 \register_reg[18][12]  ( .D(n664), .CK(clk), .RN(n2216), .Q(
        \register[18][12] ) );
  DFFRX1 \register_reg[18][11]  ( .D(n663), .CK(clk), .RN(n2216), .Q(
        \register[18][11] ) );
  DFFRX1 \register_reg[18][10]  ( .D(n662), .CK(clk), .RN(n2216), .Q(
        \register[18][10] ) );
  DFFRX1 \register_reg[18][9]  ( .D(n661), .CK(clk), .RN(n2216), .Q(
        \register[18][9] ) );
  DFFRX1 \register_reg[18][8]  ( .D(n660), .CK(clk), .RN(n2216), .Q(
        \register[18][8] ) );
  DFFRX1 \register_reg[18][7]  ( .D(n659), .CK(clk), .RN(n2215), .Q(
        \register[18][7] ) );
  DFFRX1 \register_reg[18][6]  ( .D(n658), .CK(clk), .RN(n2215), .Q(
        \register[18][6] ) );
  DFFRX1 \register_reg[18][5]  ( .D(n657), .CK(clk), .RN(n2215), .Q(
        \register[18][5] ) );
  DFFRX1 \register_reg[18][4]  ( .D(n656), .CK(clk), .RN(n2215), .Q(
        \register[18][4] ) );
  DFFRX1 \register_reg[18][3]  ( .D(n655), .CK(clk), .RN(n2215), .Q(
        \register[18][3] ) );
  DFFRX1 \register_reg[18][2]  ( .D(n654), .CK(clk), .RN(n2215), .Q(
        \register[18][2] ) );
  DFFRX1 \register_reg[18][1]  ( .D(n653), .CK(clk), .RN(n2215), .Q(
        \register[18][1] ) );
  DFFRX1 \register_reg[18][0]  ( .D(n652), .CK(clk), .RN(n2215), .Q(
        \register[18][0] ) );
  DFFRX1 \register_reg[14][31]  ( .D(n555), .CK(clk), .RN(n2223), .Q(
        \register[14][31] ) );
  DFFRX1 \register_reg[14][30]  ( .D(n554), .CK(clk), .RN(n2223), .Q(
        \register[14][30] ) );
  DFFRX1 \register_reg[14][29]  ( .D(n553), .CK(clk), .RN(n2223), .Q(
        \register[14][29] ) );
  DFFRX1 \register_reg[14][28]  ( .D(n552), .CK(clk), .RN(n2223), .Q(
        \register[14][28] ) );
  DFFRX1 \register_reg[14][27]  ( .D(n551), .CK(clk), .RN(n2222), .Q(
        \register[14][27] ) );
  DFFRX1 \register_reg[14][26]  ( .D(n550), .CK(clk), .RN(n2222), .Q(
        \register[14][26] ) );
  DFFRX1 \register_reg[14][25]  ( .D(n549), .CK(clk), .RN(n2222), .Q(
        \register[14][25] ) );
  DFFRX1 \register_reg[14][24]  ( .D(n548), .CK(clk), .RN(n2222), .Q(
        \register[14][24] ) );
  DFFRX1 \register_reg[14][23]  ( .D(n547), .CK(clk), .RN(n2222), .Q(
        \register[14][23] ) );
  DFFRX1 \register_reg[14][22]  ( .D(n546), .CK(clk), .RN(n2222), .Q(
        \register[14][22] ) );
  DFFRX1 \register_reg[14][21]  ( .D(n545), .CK(clk), .RN(n2222), .Q(
        \register[14][21] ) );
  DFFRX1 \register_reg[14][20]  ( .D(n544), .CK(clk), .RN(n2222), .Q(
        \register[14][20] ) );
  DFFRX1 \register_reg[14][19]  ( .D(n543), .CK(clk), .RN(n2222), .Q(
        \register[14][19] ) );
  DFFRX1 \register_reg[14][18]  ( .D(n542), .CK(clk), .RN(n2222), .Q(
        \register[14][18] ) );
  DFFRX1 \register_reg[14][17]  ( .D(n541), .CK(clk), .RN(n2222), .Q(
        \register[14][17] ) );
  DFFRX1 \register_reg[14][16]  ( .D(n540), .CK(clk), .RN(n2222), .Q(
        \register[14][16] ) );
  DFFRX1 \register_reg[14][15]  ( .D(n539), .CK(clk), .RN(n2221), .Q(
        \register[14][15] ) );
  DFFRX1 \register_reg[14][14]  ( .D(n538), .CK(clk), .RN(n2221), .Q(
        \register[14][14] ) );
  DFFRX1 \register_reg[14][13]  ( .D(n537), .CK(clk), .RN(n2221), .Q(
        \register[14][13] ) );
  DFFRX1 \register_reg[14][12]  ( .D(n536), .CK(clk), .RN(n2221), .Q(
        \register[14][12] ) );
  DFFRX1 \register_reg[14][11]  ( .D(n535), .CK(clk), .RN(n2221), .Q(
        \register[14][11] ) );
  DFFRX1 \register_reg[14][10]  ( .D(n534), .CK(clk), .RN(n2221), .Q(
        \register[14][10] ) );
  DFFRX1 \register_reg[14][9]  ( .D(n533), .CK(clk), .RN(n2221), .Q(
        \register[14][9] ) );
  DFFRX1 \register_reg[14][8]  ( .D(n532), .CK(clk), .RN(n2221), .Q(
        \register[14][8] ) );
  DFFRX1 \register_reg[14][7]  ( .D(n531), .CK(clk), .RN(n2221), .Q(
        \register[14][7] ) );
  DFFRX1 \register_reg[14][6]  ( .D(n530), .CK(clk), .RN(n2221), .Q(
        \register[14][6] ) );
  DFFRX1 \register_reg[14][5]  ( .D(n529), .CK(clk), .RN(n2221), .Q(
        \register[14][5] ) );
  DFFRX1 \register_reg[14][4]  ( .D(n528), .CK(clk), .RN(n2221), .Q(
        \register[14][4] ) );
  DFFRX1 \register_reg[14][3]  ( .D(n527), .CK(clk), .RN(n2204), .Q(
        \register[14][3] ) );
  DFFRX1 \register_reg[14][2]  ( .D(n526), .CK(clk), .RN(n2204), .Q(
        \register[14][2] ) );
  DFFRX1 \register_reg[14][1]  ( .D(n525), .CK(clk), .RN(n2204), .Q(
        \register[14][1] ) );
  DFFRX1 \register_reg[14][0]  ( .D(n524), .CK(clk), .RN(n2204), .Q(
        \register[14][0] ) );
  DFFRX1 \register_reg[10][31]  ( .D(n427), .CK(clk), .RN(n2212), .Q(
        \register[10][31] ) );
  DFFRX1 \register_reg[10][30]  ( .D(n426), .CK(clk), .RN(n2212), .Q(
        \register[10][30] ) );
  DFFRX1 \register_reg[10][29]  ( .D(n425), .CK(clk), .RN(n2212), .Q(
        \register[10][29] ) );
  DFFRX1 \register_reg[10][28]  ( .D(n424), .CK(clk), .RN(n2212), .Q(
        \register[10][28] ) );
  DFFRX1 \register_reg[10][27]  ( .D(n423), .CK(clk), .RN(n2212), .Q(
        \register[10][27] ) );
  DFFRX1 \register_reg[10][26]  ( .D(n422), .CK(clk), .RN(n2212), .Q(
        \register[10][26] ) );
  DFFRX1 \register_reg[10][25]  ( .D(n421), .CK(clk), .RN(n2212), .Q(
        \register[10][25] ) );
  DFFRX1 \register_reg[10][24]  ( .D(n420), .CK(clk), .RN(n2212), .Q(
        \register[10][24] ) );
  DFFRX1 \register_reg[10][23]  ( .D(n419), .CK(clk), .RN(n2211), .Q(
        \register[10][23] ) );
  DFFRX1 \register_reg[10][22]  ( .D(n418), .CK(clk), .RN(n2211), .Q(
        \register[10][22] ) );
  DFFRX1 \register_reg[10][21]  ( .D(n417), .CK(clk), .RN(n2211), .Q(
        \register[10][21] ) );
  DFFRX1 \register_reg[10][20]  ( .D(n416), .CK(clk), .RN(n2211), .Q(
        \register[10][20] ) );
  DFFRX1 \register_reg[10][19]  ( .D(n415), .CK(clk), .RN(n2211), .Q(
        \register[10][19] ) );
  DFFRX1 \register_reg[10][18]  ( .D(n414), .CK(clk), .RN(n2211), .Q(
        \register[10][18] ) );
  DFFRX1 \register_reg[10][17]  ( .D(n413), .CK(clk), .RN(n2211), .Q(
        \register[10][17] ) );
  DFFRX1 \register_reg[10][16]  ( .D(n412), .CK(clk), .RN(n2211), .Q(
        \register[10][16] ) );
  DFFRX1 \register_reg[10][15]  ( .D(n411), .CK(clk), .RN(n2211), .Q(
        \register[10][15] ) );
  DFFRX1 \register_reg[10][14]  ( .D(n410), .CK(clk), .RN(n2211), .Q(
        \register[10][14] ) );
  DFFRX1 \register_reg[10][13]  ( .D(n409), .CK(clk), .RN(n2211), .Q(
        \register[10][13] ) );
  DFFRX1 \register_reg[10][12]  ( .D(n408), .CK(clk), .RN(n2211), .Q(
        \register[10][12] ) );
  DFFRX1 \register_reg[10][11]  ( .D(n407), .CK(clk), .RN(n2210), .Q(
        \register[10][11] ) );
  DFFRX1 \register_reg[10][10]  ( .D(n406), .CK(clk), .RN(n2210), .Q(
        \register[10][10] ) );
  DFFRX1 \register_reg[10][9]  ( .D(n405), .CK(clk), .RN(n2210), .Q(
        \register[10][9] ) );
  DFFRX1 \register_reg[10][8]  ( .D(n404), .CK(clk), .RN(n2210), .Q(
        \register[10][8] ) );
  DFFRX1 \register_reg[10][7]  ( .D(n403), .CK(clk), .RN(n2210), .Q(
        \register[10][7] ) );
  DFFRX1 \register_reg[10][6]  ( .D(n402), .CK(clk), .RN(n2210), .Q(
        \register[10][6] ) );
  DFFRX1 \register_reg[10][5]  ( .D(n401), .CK(clk), .RN(n2210), .Q(
        \register[10][5] ) );
  DFFRX1 \register_reg[10][4]  ( .D(n400), .CK(clk), .RN(n2210), .Q(
        \register[10][4] ) );
  DFFRX1 \register_reg[10][3]  ( .D(n399), .CK(clk), .RN(n2210), .Q(
        \register[10][3] ) );
  DFFRX1 \register_reg[10][2]  ( .D(n398), .CK(clk), .RN(n2210), .Q(
        \register[10][2] ) );
  DFFRX1 \register_reg[10][1]  ( .D(n397), .CK(clk), .RN(n2210), .Q(
        \register[10][1] ) );
  DFFRX1 \register_reg[10][0]  ( .D(n396), .CK(clk), .RN(n2210), .Q(
        \register[10][0] ) );
  DFFRX1 \register_reg[6][31]  ( .D(n299), .CK(clk), .RN(n2193), .Q(
        \register[6][31] ) );
  DFFRX1 \register_reg[6][30]  ( .D(n298), .CK(clk), .RN(n2193), .Q(
        \register[6][30] ) );
  DFFRX1 \register_reg[6][29]  ( .D(n297), .CK(clk), .RN(n2193), .Q(
        \register[6][29] ) );
  DFFRX1 \register_reg[6][28]  ( .D(n296), .CK(clk), .RN(n2193), .Q(
        \register[6][28] ) );
  DFFRX1 \register_reg[6][27]  ( .D(n295), .CK(clk), .RN(n2193), .Q(
        \register[6][27] ) );
  DFFRX1 \register_reg[6][26]  ( .D(n294), .CK(clk), .RN(n2193), .Q(
        \register[6][26] ) );
  DFFRX1 \register_reg[6][25]  ( .D(n293), .CK(clk), .RN(n2193), .Q(
        \register[6][25] ) );
  DFFRX1 \register_reg[6][24]  ( .D(n292), .CK(clk), .RN(n2193), .Q(
        \register[6][24] ) );
  DFFRX1 \register_reg[6][23]  ( .D(n291), .CK(clk), .RN(n2193), .Q(
        \register[6][23] ) );
  DFFRX1 \register_reg[6][22]  ( .D(n290), .CK(clk), .RN(n2193), .Q(
        \register[6][22] ) );
  DFFRX1 \register_reg[6][21]  ( .D(n289), .CK(clk), .RN(n2193), .Q(
        \register[6][21] ) );
  DFFRX1 \register_reg[6][20]  ( .D(n288), .CK(clk), .RN(n2193), .Q(
        \register[6][20] ) );
  DFFRX1 \register_reg[6][19]  ( .D(n287), .CK(clk), .RN(n2200), .Q(
        \register[6][19] ) );
  DFFRX1 \register_reg[6][18]  ( .D(n286), .CK(clk), .RN(n2200), .Q(
        \register[6][18] ) );
  DFFRX1 \register_reg[6][17]  ( .D(n285), .CK(clk), .RN(n2200), .Q(
        \register[6][17] ) );
  DFFRX1 \register_reg[6][16]  ( .D(n284), .CK(clk), .RN(n2200), .Q(
        \register[6][16] ) );
  DFFRX1 \register_reg[6][15]  ( .D(n283), .CK(clk), .RN(n2200), .Q(
        \register[6][15] ) );
  DFFRX1 \register_reg[6][14]  ( .D(n282), .CK(clk), .RN(n2200), .Q(
        \register[6][14] ) );
  DFFRX1 \register_reg[6][13]  ( .D(n281), .CK(clk), .RN(n2200), .Q(
        \register[6][13] ) );
  DFFRX1 \register_reg[6][12]  ( .D(n280), .CK(clk), .RN(n2200), .Q(
        \register[6][12] ) );
  DFFRX1 \register_reg[6][11]  ( .D(n279), .CK(clk), .RN(n2200), .Q(
        \register[6][11] ) );
  DFFRX1 \register_reg[6][10]  ( .D(n278), .CK(clk), .RN(n2200), .Q(
        \register[6][10] ) );
  DFFRX1 \register_reg[6][9]  ( .D(n277), .CK(clk), .RN(n2200), .Q(
        \register[6][9] ) );
  DFFRX1 \register_reg[6][8]  ( .D(n276), .CK(clk), .RN(n2200), .Q(
        \register[6][8] ) );
  DFFRX1 \register_reg[6][7]  ( .D(n275), .CK(clk), .RN(n2199), .Q(
        \register[6][7] ) );
  DFFRX1 \register_reg[6][6]  ( .D(n274), .CK(clk), .RN(n2199), .Q(
        \register[6][6] ) );
  DFFRX1 \register_reg[6][5]  ( .D(n273), .CK(clk), .RN(n2199), .Q(
        \register[6][5] ) );
  DFFRX1 \register_reg[6][4]  ( .D(n272), .CK(clk), .RN(n2199), .Q(
        \register[6][4] ) );
  DFFRX1 \register_reg[6][3]  ( .D(n271), .CK(clk), .RN(n2199), .Q(
        \register[6][3] ) );
  DFFRX1 \register_reg[6][2]  ( .D(n270), .CK(clk), .RN(n2199), .Q(
        \register[6][2] ) );
  DFFRX1 \register_reg[6][1]  ( .D(n269), .CK(clk), .RN(n2199), .Q(
        \register[6][1] ) );
  DFFRX1 \register_reg[6][0]  ( .D(n268), .CK(clk), .RN(n2199), .Q(
        \register[6][0] ) );
  DFFRX1 \register_reg[3][31]  ( .D(n203), .CK(clk), .RN(n2178), .Q(
        \register[3][31] ) );
  DFFRX1 \register_reg[3][30]  ( .D(n202), .CK(clk), .RN(n2178), .Q(
        \register[3][30] ) );
  DFFRX1 \register_reg[3][29]  ( .D(n201), .CK(clk), .RN(n2178), .Q(
        \register[3][29] ) );
  DFFRX1 \register_reg[3][28]  ( .D(n200), .CK(clk), .RN(n2178), .Q(
        \register[3][28] ) );
  DFFRX1 \register_reg[3][27]  ( .D(n199), .CK(clk), .RN(n2178), .Q(
        \register[3][27] ) );
  DFFRX1 \register_reg[3][26]  ( .D(n198), .CK(clk), .RN(n2178), .Q(
        \register[3][26] ) );
  DFFRX1 \register_reg[3][25]  ( .D(n197), .CK(clk), .RN(n2178), .Q(
        \register[3][25] ) );
  DFFRX1 \register_reg[3][24]  ( .D(n196), .CK(clk), .RN(n2178), .Q(
        \register[3][24] ) );
  DFFRX1 \register_reg[3][23]  ( .D(n195), .CK(clk), .RN(n2178), .Q(
        \register[3][23] ) );
  DFFRX1 \register_reg[3][22]  ( .D(n194), .CK(clk), .RN(n2178), .Q(
        \register[3][22] ) );
  DFFRX1 \register_reg[3][21]  ( .D(n193), .CK(clk), .RN(n2178), .Q(
        \register[3][21] ) );
  DFFRX1 \register_reg[3][20]  ( .D(n192), .CK(clk), .RN(n2178), .Q(
        \register[3][20] ) );
  DFFRX1 \register_reg[3][19]  ( .D(n191), .CK(clk), .RN(n2185), .Q(
        \register[3][19] ) );
  DFFRX1 \register_reg[3][18]  ( .D(n190), .CK(clk), .RN(n2185), .Q(
        \register[3][18] ) );
  DFFRX1 \register_reg[3][17]  ( .D(n189), .CK(clk), .RN(n2185), .Q(
        \register[3][17] ) );
  DFFRX1 \register_reg[3][16]  ( .D(n188), .CK(clk), .RN(n2185), .Q(
        \register[3][16] ) );
  DFFRX1 \register_reg[3][15]  ( .D(n187), .CK(clk), .RN(n2185), .Q(
        \register[3][15] ) );
  DFFRX1 \register_reg[3][14]  ( .D(n186), .CK(clk), .RN(n2185), .Q(
        \register[3][14] ) );
  DFFRX1 \register_reg[3][13]  ( .D(n185), .CK(clk), .RN(n2185), .Q(
        \register[3][13] ) );
  DFFRX1 \register_reg[3][12]  ( .D(n184), .CK(clk), .RN(n2185), .Q(
        \register[3][12] ) );
  DFFRX1 \register_reg[3][11]  ( .D(n183), .CK(clk), .RN(n2185), .Q(
        \register[3][11] ) );
  DFFRX1 \register_reg[3][10]  ( .D(n182), .CK(clk), .RN(n2185), .Q(
        \register[3][10] ) );
  DFFRX1 \register_reg[3][9]  ( .D(n181), .CK(clk), .RN(n2185), .Q(
        \register[3][9] ) );
  DFFRX1 \register_reg[3][8]  ( .D(n180), .CK(clk), .RN(n2185), .Q(
        \register[3][8] ) );
  DFFRX1 \register_reg[3][7]  ( .D(n179), .CK(clk), .RN(n2184), .Q(
        \register[3][7] ) );
  DFFRX1 \register_reg[3][6]  ( .D(n178), .CK(clk), .RN(n2184), .Q(
        \register[3][6] ) );
  DFFRX1 \register_reg[3][5]  ( .D(n177), .CK(clk), .RN(n2184), .Q(
        \register[3][5] ) );
  DFFRX1 \register_reg[3][4]  ( .D(n176), .CK(clk), .RN(n2184), .Q(
        \register[3][4] ) );
  DFFRX1 \register_reg[3][3]  ( .D(n175), .CK(clk), .RN(n2184), .Q(
        \register[3][3] ) );
  DFFRX1 \register_reg[3][2]  ( .D(n174), .CK(clk), .RN(n2184), .Q(
        \register[3][2] ) );
  DFFRX1 \register_reg[3][1]  ( .D(n173), .CK(clk), .RN(n2184), .Q(
        \register[3][1] ) );
  DFFRX1 \register_reg[3][0]  ( .D(n172), .CK(clk), .RN(n2184), .Q(
        \register[3][0] ) );
  DFFRX1 \register_reg[1][31]  ( .D(n139), .CK(clk), .RN(n2188), .Q(
        \register[1][31] ) );
  DFFRX1 \register_reg[1][30]  ( .D(n138), .CK(clk), .RN(n2188), .Q(
        \register[1][30] ) );
  DFFRX1 \register_reg[1][29]  ( .D(n137), .CK(clk), .RN(n2188), .Q(
        \register[1][29] ) );
  DFFRX1 \register_reg[1][28]  ( .D(n136), .CK(clk), .RN(n2188), .Q(
        \register[1][28] ) );
  DFFRX1 \register_reg[1][27]  ( .D(n135), .CK(clk), .RN(n2188), .Q(
        \register[1][27] ) );
  DFFRX1 \register_reg[1][26]  ( .D(n134), .CK(clk), .RN(n2188), .Q(
        \register[1][26] ) );
  DFFRX1 \register_reg[1][25]  ( .D(n133), .CK(clk), .RN(n2188), .Q(
        \register[1][25] ) );
  DFFRX1 \register_reg[1][24]  ( .D(n132), .CK(clk), .RN(n2188), .Q(
        \register[1][24] ) );
  DFFRX1 \register_reg[1][23]  ( .D(n131), .CK(clk), .RN(n2187), .Q(
        \register[1][23] ) );
  DFFRX1 \register_reg[1][22]  ( .D(n130), .CK(clk), .RN(n2187), .Q(
        \register[1][22] ) );
  DFFRX1 \register_reg[1][21]  ( .D(n129), .CK(clk), .RN(n2187), .Q(
        \register[1][21] ) );
  DFFRX1 \register_reg[1][20]  ( .D(n128), .CK(clk), .RN(n2187), .Q(
        \register[1][20] ) );
  DFFRX1 \register_reg[1][19]  ( .D(n127), .CK(clk), .RN(n2187), .Q(
        \register[1][19] ) );
  DFFRX1 \register_reg[1][18]  ( .D(n126), .CK(clk), .RN(n2187), .Q(
        \register[1][18] ) );
  DFFRX1 \register_reg[1][17]  ( .D(n125), .CK(clk), .RN(n2187), .Q(
        \register[1][17] ) );
  DFFRX1 \register_reg[1][16]  ( .D(n124), .CK(clk), .RN(n2187), .Q(
        \register[1][16] ) );
  DFFRX1 \register_reg[1][15]  ( .D(n123), .CK(clk), .RN(n2187), .Q(
        \register[1][15] ) );
  DFFRX1 \register_reg[1][14]  ( .D(n122), .CK(clk), .RN(n2187), .Q(
        \register[1][14] ) );
  DFFRX1 \register_reg[1][13]  ( .D(n121), .CK(clk), .RN(n2187), .Q(
        \register[1][13] ) );
  DFFRX1 \register_reg[1][12]  ( .D(n120), .CK(clk), .RN(n2187), .Q(
        \register[1][12] ) );
  DFFRX1 \register_reg[1][11]  ( .D(n119), .CK(clk), .RN(n2186), .Q(
        \register[1][11] ) );
  DFFRX1 \register_reg[1][10]  ( .D(n118), .CK(clk), .RN(n2186), .Q(
        \register[1][10] ) );
  DFFRX1 \register_reg[1][9]  ( .D(n117), .CK(clk), .RN(n2186), .Q(
        \register[1][9] ) );
  DFFRX1 \register_reg[1][8]  ( .D(n116), .CK(clk), .RN(n2186), .Q(
        \register[1][8] ) );
  DFFRX1 \register_reg[1][7]  ( .D(n115), .CK(clk), .RN(n2186), .Q(
        \register[1][7] ) );
  DFFRX1 \register_reg[1][6]  ( .D(n114), .CK(clk), .RN(n2186), .Q(
        \register[1][6] ) );
  DFFRX1 \register_reg[1][5]  ( .D(n113), .CK(clk), .RN(n2186), .Q(
        \register[1][5] ) );
  DFFRX1 \register_reg[1][4]  ( .D(n112), .CK(clk), .RN(n2186), .Q(
        \register[1][4] ) );
  DFFRX1 \register_reg[1][3]  ( .D(n111), .CK(clk), .RN(n2186), .Q(
        \register[1][3] ) );
  DFFRX1 \register_reg[1][2]  ( .D(n110), .CK(clk), .RN(n2186), .Q(
        \register[1][2] ) );
  DFFRX1 \register_reg[1][1]  ( .D(n109), .CK(clk), .RN(n2186), .Q(
        \register[1][1] ) );
  DFFRX1 \register_reg[1][0]  ( .D(n108), .CK(clk), .RN(n2186), .Q(
        \register[1][0] ) );
  DFFRX1 \register_reg[2][31]  ( .D(n171), .CK(clk), .RN(n2184), .Q(
        \register[2][31] ), .QN(n2582) );
  DFFRX1 \register_reg[2][30]  ( .D(n170), .CK(clk), .RN(n2184), .Q(
        \register[2][30] ), .QN(n2581) );
  DFFRX1 \register_reg[2][23]  ( .D(n163), .CK(clk), .RN(n2183), .Q(
        \register[2][23] ), .QN(n2574) );
  DFFRX1 \register_reg[2][24]  ( .D(n164), .CK(clk), .RN(n2183), .Q(
        \register[2][24] ), .QN(n2575) );
  DFFRX1 \register_reg[2][22]  ( .D(n162), .CK(clk), .RN(n2183), .Q(
        \register[2][22] ), .QN(n2573) );
  DFFRX1 \register_reg[2][16]  ( .D(n156), .CK(clk), .RN(n2183), .Q(
        \register[2][16] ), .QN(n2567) );
  DFFRX1 \register_reg[2][14]  ( .D(n154), .CK(clk), .RN(n2182), .Q(
        \register[2][14] ), .QN(n2565) );
  DFFRX1 \register_reg[2][13]  ( .D(n153), .CK(clk), .RN(n2182), .Q(
        \register[2][13] ), .QN(n2564) );
  DFFRX1 \register_reg[2][12]  ( .D(n152), .CK(clk), .RN(n2182), .Q(
        \register[2][12] ), .QN(n2563) );
  DFFRX1 \register_reg[2][11]  ( .D(n151), .CK(clk), .RN(n2182), .Q(
        \register[2][11] ), .QN(n2562) );
  DFFRX1 \register_reg[2][10]  ( .D(n150), .CK(clk), .RN(n2182), .Q(
        \register[2][10] ), .QN(n2561) );
  DFFRX1 \register_reg[2][9]  ( .D(n149), .CK(clk), .RN(n2182), .Q(
        \register[2][9] ), .QN(n2560) );
  DFFRX1 \register_reg[2][8]  ( .D(n148), .CK(clk), .RN(n2182), .Q(
        \register[2][8] ), .QN(n2559) );
  DFFRX1 \register_reg[2][7]  ( .D(n147), .CK(clk), .RN(n2182), .Q(
        \register[2][7] ), .QN(n2558) );
  DFFRX1 \register_reg[2][6]  ( .D(n146), .CK(clk), .RN(n2182), .Q(
        \register[2][6] ), .QN(n2557) );
  DFFRX1 \register_reg[2][5]  ( .D(n145), .CK(clk), .RN(n2182), .Q(
        \register[2][5] ), .QN(n2556) );
  DFFRX1 \register_reg[2][3]  ( .D(n143), .CK(clk), .RN(n2188), .Q(
        \register[2][3] ), .QN(n2554) );
  DFFRX1 \register_reg[2][29]  ( .D(n169), .CK(clk), .RN(n2184), .Q(
        \register[2][29] ), .QN(n2580) );
  DFFRX1 \register_reg[2][28]  ( .D(n168), .CK(clk), .RN(n2184), .Q(
        \register[2][28] ), .QN(n2579) );
  DFFRX1 \register_reg[2][27]  ( .D(n167), .CK(clk), .RN(n2183), .Q(
        \register[2][27] ), .QN(n2578) );
  DFFRX1 \register_reg[2][26]  ( .D(n166), .CK(clk), .RN(n2183), .Q(
        \register[2][26] ), .QN(n2577) );
  DFFRX1 \register_reg[2][25]  ( .D(n165), .CK(clk), .RN(n2183), .Q(
        \register[2][25] ), .QN(n2576) );
  CLKINVX4 U3 ( .A(n1), .Y(n2) );
  INVXL U4 ( .A(wdata[6]), .Y(n2608) );
  CLKBUFX3 U5 ( .A(n2608), .Y(n2350) );
  CLKBUFX2 U6 ( .A(rst_n), .Y(n2289) );
  CLKBUFX2 U7 ( .A(rst_n), .Y(n2288) );
  CLKBUFX3 U8 ( .A(N12), .Y(n2546) );
  CLKBUFX3 U9 ( .A(N17), .Y(n2544) );
  BUFX2 U10 ( .A(N18), .Y(n2545) );
  OR3XL U11 ( .A(wsel[3]), .B(wsel[4]), .C(n2620), .Y(n1) );
  CLKBUFX2 U12 ( .A(n2128), .Y(n2129) );
  BUFX4 U13 ( .A(n2126), .Y(n2143) );
  INVX1 U14 ( .A(wdata[0]), .Y(n2614) );
  INVX2 U15 ( .A(wdata[1]), .Y(n2613) );
  INVX2 U16 ( .A(wdata[2]), .Y(n2612) );
  INVX2 U17 ( .A(wdata[4]), .Y(n2610) );
  BUFX2 U18 ( .A(n2548), .Y(n1574) );
  BUFX2 U19 ( .A(n88), .Y(n2458) );
  BUFX2 U20 ( .A(n97), .Y(n2413) );
  BUFX2 U21 ( .A(n106), .Y(n2371) );
  BUFX2 U22 ( .A(n103), .Y(n2386) );
  BUFX2 U23 ( .A(n70), .Y(n2517) );
  BUFX2 U24 ( .A(n95), .Y(n2424) );
  BUFX2 U25 ( .A(n72), .Y(n2513) );
  BUFX2 U26 ( .A(N13), .Y(n1576) );
  BUFX2 U27 ( .A(N21), .Y(n2109) );
  BUFX2 U28 ( .A(N18), .Y(n2127) );
  BUFX2 U29 ( .A(n10), .Y(n2406) );
  BUFX2 U30 ( .A(n8), .Y(n2418) );
  BUFX2 U31 ( .A(n2550), .Y(n1559) );
  BUFX2 U32 ( .A(n2125), .Y(n2118) );
  BUFX2 U33 ( .A(n2125), .Y(n2117) );
  BUFX4 U34 ( .A(N20), .Y(n2116) );
  BUFX2 U35 ( .A(n5), .Y(n2496) );
  BUFX2 U36 ( .A(n6), .Y(n2508) );
  BUFX2 U37 ( .A(n7), .Y(n2463) );
  BUFX2 U38 ( .A(n4), .Y(n2376) );
  BUFX2 U39 ( .A(n9), .Y(n2451) );
  BUFX2 U40 ( .A(n3), .Y(n2364) );
  BUFX4 U41 ( .A(n2539), .Y(n2543) );
  BUFX2 U42 ( .A(n2533), .Y(n2536) );
  CLKBUFX2 U43 ( .A(n101), .Y(n2397) );
  CLKBUFX2 U44 ( .A(n84), .Y(n2481) );
  CLKBUFX2 U45 ( .A(n102), .Y(n2391) );
  NOR3X4 U46 ( .A(wsel[1]), .B(wsel[2]), .C(wsel[0]), .Y(n82) );
  NOR3X4 U47 ( .A(wsel[0]), .B(wsel[2]), .C(n2618), .Y(n69) );
  INVX3 U48 ( .A(wsel[1]), .Y(n2618) );
  AND2X2 U49 ( .A(n71), .B(n2), .Y(n14) );
  AND2X1 U50 ( .A(n91), .B(n71), .Y(n16) );
  CLKAND2X2 U51 ( .A(n100), .B(n71), .Y(n12) );
  NOR3X1 U52 ( .A(n2619), .B(wsel[2]), .C(n2618), .Y(n71) );
  NOR3X4 U53 ( .A(wsel[1]), .B(wsel[2]), .C(n2619), .Y(n66) );
  INVX6 U54 ( .A(wsel[0]), .Y(n2619) );
  NOR3X6 U55 ( .A(n2616), .B(n2615), .C(n2620), .Y(n100) );
  XNOR2X2 U56 ( .A(n2616), .B(n2549), .Y(n63) );
  INVX6 U57 ( .A(wsel[3]), .Y(n2616) );
  NOR3X2 U58 ( .A(n2615), .B(wsel[3]), .C(n2620), .Y(n91) );
  INVXL U59 ( .A(wdata[3]), .Y(n2611) );
  INVX4 U60 ( .A(wsel[2]), .Y(n2617) );
  CLKINVX6 U61 ( .A(wsel[4]), .Y(n2615) );
  NOR3X6 U62 ( .A(n2616), .B(wsel[4]), .C(n2620), .Y(n81) );
  AND2X2 U63 ( .A(n91), .B(n82), .Y(n30) );
  AND2X2 U64 ( .A(n100), .B(n82), .Y(n31) );
  AND2X2 U65 ( .A(n81), .B(n82), .Y(n29) );
  AND2X2 U66 ( .A(n91), .B(n73), .Y(n24) );
  AND2X2 U67 ( .A(n81), .B(n73), .Y(n23) );
  AND2X2 U68 ( .A(n73), .B(n2), .Y(n20) );
  AND2X2 U69 ( .A(n100), .B(n73), .Y(n25) );
  NOR3X1 U70 ( .A(wsel[0]), .B(wsel[1]), .C(n2617), .Y(n73) );
  NOR3X1 U71 ( .A(n2618), .B(wsel[0]), .C(n2617), .Y(n77) );
  NOR2XL U72 ( .A(n1596), .B(n1625), .Y(n1552) );
  CLKBUFX4 U73 ( .A(n2156), .Y(n2172) );
  BUFX2 U74 ( .A(n2130), .Y(n2150) );
  BUFX8 U75 ( .A(n1605), .Y(n1624) );
  BUFX2 U76 ( .A(n1579), .Y(n1599) );
  CLKBUFX6 U77 ( .A(n1560), .Y(n1562) );
  BUFX8 U78 ( .A(n2110), .Y(n2112) );
  CLKBUFX2 U79 ( .A(n2110), .Y(n2111) );
  CLKBUFX2 U80 ( .A(n1560), .Y(n1561) );
  CLKBUFX2 U81 ( .A(n2118), .Y(n2119) );
  CLKBUFX2 U82 ( .A(n1574), .Y(n1568) );
  BUFX2 U83 ( .A(n2533), .Y(n2535) );
  NOR2X1 U84 ( .A(n2150), .B(\register[1][20] ), .Y(n2003) );
  MXI2XL U85 ( .A(n2565), .B(n1481), .S0(n1621), .Y(n1484) );
  MXI2XL U86 ( .A(n2558), .B(n1516), .S0(n1621), .Y(n1519) );
  MXI2XL U87 ( .A(n2560), .B(n1506), .S0(n1621), .Y(n1509) );
  MXI2XL U88 ( .A(n2556), .B(n1526), .S0(n1621), .Y(n1529) );
  MXI4XL U89 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n1615), .S1(n1590), .Y(
        n1148) );
  MXI4XL U90 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n1619), .S1(n1594), 
        .Y(n1252) );
  MXI4XL U91 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n1616), .S1(n1590), .Y(
        n1150) );
  BUFX8 U92 ( .A(n1605), .Y(n1625) );
  MXI2X1 U93 ( .A(n2571), .B(n2001), .S0(n2174), .Y(n2004) );
  CLKBUFX4 U94 ( .A(n1606), .Y(n1620) );
  BUFX4 U95 ( .A(n2154), .Y(n2157) );
  BUFX4 U96 ( .A(n1602), .Y(n1607) );
  NOR4X1 U97 ( .A(n64), .B(n2548), .C(n2550), .D(n2549), .Y(n61) );
  NAND2X1 U98 ( .A(n100), .B(n79), .Y(n3) );
  NAND2X1 U99 ( .A(n100), .B(n75), .Y(n4) );
  XNOR2X1 U100 ( .A(n2615), .B(n2550), .Y(n62) );
  INVXL U101 ( .A(wdata[15]), .Y(n2599) );
  INVXL U102 ( .A(wdata[10]), .Y(n2604) );
  INVXL U103 ( .A(wdata[16]), .Y(n2598) );
  INVXL U104 ( .A(wdata[7]), .Y(n2607) );
  INVXL U105 ( .A(wdata[20]), .Y(n2594) );
  INVXL U106 ( .A(wdata[28]), .Y(n2586) );
  INVXL U107 ( .A(wdata[31]), .Y(n2583) );
  INVXL U108 ( .A(wdata[24]), .Y(n2590) );
  INVXL U109 ( .A(wdata[13]), .Y(n2601) );
  INVXL U110 ( .A(wdata[23]), .Y(n2591) );
  INVXL U111 ( .A(wdata[22]), .Y(n2592) );
  INVXL U112 ( .A(wdata[29]), .Y(n2585) );
  INVXL U113 ( .A(wdata[30]), .Y(n2584) );
  INVXL U114 ( .A(wdata[26]), .Y(n2588) );
  MXI2X1 U115 ( .A(n2558), .B(n2066), .S0(n2173), .Y(n2069) );
  NOR2BX1 U116 ( .AN(n2146), .B(\register[3][20] ), .Y(n2001) );
  NOR2BX1 U117 ( .AN(n1596), .B(\register[3][1] ), .Y(n1546) );
  NOR2XL U118 ( .A(n1596), .B(n1625), .Y(n1527) );
  NOR2XL U119 ( .A(n1597), .B(n1625), .Y(n1532) );
  NOR2XL U120 ( .A(n1598), .B(n1625), .Y(n1522) );
  NOR2XL U121 ( .A(n1597), .B(n1624), .Y(n1507) );
  NOR2XL U122 ( .A(n1597), .B(n1625), .Y(n1517) );
  NOR2XL U123 ( .A(n1597), .B(n1625), .Y(n1537) );
  CLKBUFX3 U124 ( .A(n2155), .Y(n2175) );
  CLKBUFX3 U125 ( .A(n1604), .Y(n1623) );
  CLKBUFX3 U126 ( .A(n2155), .Y(n2176) );
  CLKBUFX3 U127 ( .A(n2155), .Y(n2177) );
  BUFX4 U128 ( .A(n1604), .Y(n1605) );
  BUFX4 U129 ( .A(n2127), .Y(n2132) );
  BUFX4 U130 ( .A(n2118), .Y(n2120) );
  BUFX4 U131 ( .A(n1570), .Y(n1569) );
  CLKBUFX2 U132 ( .A(n1576), .Y(n1581) );
  CLKBUFX4 U133 ( .A(n2534), .Y(n2538) );
  NOR4XL U134 ( .A(n55), .B(N19), .C(N21), .D(N20), .Y(n52) );
  OR2XL U135 ( .A(n2544), .B(n2545), .Y(n55) );
  OR2XL U136 ( .A(n2546), .B(n2547), .Y(n64) );
  CLKBUFX2 U137 ( .A(n2487), .Y(n2486) );
  CLKBUFX2 U138 ( .A(n2475), .Y(n2474) );
  BUFX2 U139 ( .A(n2549), .Y(n1567) );
  CLKBUFX2 U140 ( .A(N19), .Y(n2125) );
  AND2XL U141 ( .A(n100), .B(n66), .Y(n11) );
  INVX3 U142 ( .A(n11), .Y(n101) );
  INVX3 U143 ( .A(n12), .Y(n103) );
  CLKBUFX2 U144 ( .A(n90), .Y(n2446) );
  NOR4X2 U145 ( .A(n52), .B(n2620), .C(n53), .D(n54), .Y(n51) );
  NAND4X2 U146 ( .A(n48), .B(n49), .C(n50), .D(n51), .Y(n47) );
  NOR4X2 U147 ( .A(n61), .B(n2620), .C(n62), .D(n63), .Y(n60) );
  NAND4X2 U148 ( .A(n57), .B(n58), .C(n59), .D(n60), .Y(n56) );
  INVX3 U149 ( .A(n18), .Y(n97) );
  INVX3 U150 ( .A(n19), .Y(n106) );
  INVX3 U151 ( .A(n23), .Y(n86) );
  INVX3 U152 ( .A(n24), .Y(n95) );
  INVX3 U153 ( .A(n13), .Y(n65) );
  INVX3 U154 ( .A(n14), .Y(n70) );
  AND2XL U155 ( .A(n91), .B(n66), .Y(n15) );
  INVX3 U156 ( .A(n15), .Y(n92) );
  INVX3 U157 ( .A(n16), .Y(n94) );
  INVX3 U158 ( .A(n26), .Y(n84) );
  INVX3 U159 ( .A(n27), .Y(n93) );
  AND2XL U160 ( .A(n100), .B(n69), .Y(n28) );
  INVX3 U161 ( .A(n28), .Y(n102) );
  INVX3 U162 ( .A(n25), .Y(n104) );
  CLKBUFX2 U163 ( .A(N16), .Y(n2550) );
  INVXL U164 ( .A(wdata[14]), .Y(n2600) );
  INVXL U165 ( .A(wdata[8]), .Y(n2606) );
  INVXL U166 ( .A(wdata[11]), .Y(n2603) );
  CLKINVX1 U167 ( .A(wdata[9]), .Y(n2605) );
  CLKINVX1 U168 ( .A(wdata[27]), .Y(n2587) );
  CLKINVX1 U169 ( .A(wdata[18]), .Y(n2596) );
  INVXL U170 ( .A(wdata[19]), .Y(n2595) );
  INVXL U171 ( .A(wdata[21]), .Y(n2593) );
  INVXL U172 ( .A(wdata[25]), .Y(n2589) );
  INVXL U173 ( .A(wdata[5]), .Y(n2609) );
  INVXL U174 ( .A(wdata[12]), .Y(n2602) );
  INVXL U175 ( .A(wdata[17]), .Y(n2597) );
  AND2XL U176 ( .A(n81), .B(n77), .Y(n17) );
  INVX3 U177 ( .A(n17), .Y(n88) );
  AND2XL U178 ( .A(n77), .B(n2), .Y(n21) );
  INVX3 U179 ( .A(n21), .Y(n76) );
  AND2XL U180 ( .A(n69), .B(n2), .Y(n22) );
  INVX3 U181 ( .A(n22), .Y(n68) );
  NAND2X1 U182 ( .A(n79), .B(n2), .Y(n5) );
  NAND2X1 U183 ( .A(n75), .B(n2), .Y(n6) );
  NAND2X1 U184 ( .A(n81), .B(n75), .Y(n7) );
  NAND2X1 U185 ( .A(n91), .B(n75), .Y(n8) );
  NAND2X1 U186 ( .A(n81), .B(n79), .Y(n9) );
  NAND2X1 U187 ( .A(n91), .B(n79), .Y(n10) );
  INVX3 U188 ( .A(n20), .Y(n72) );
  MXI2XL U189 ( .A(n2552), .B(n1546), .S0(n1620), .Y(n1549) );
  NOR2XL U190 ( .A(n1597), .B(\register[1][9] ), .Y(n1508) );
  NOR2XL U191 ( .A(n1597), .B(\register[1][5] ), .Y(n1528) );
  NOR2XL U192 ( .A(n1597), .B(\register[1][7] ), .Y(n1518) );
  NOR2XL U193 ( .A(n1596), .B(\register[1][4] ), .Y(n1533) );
  NOR2XL U194 ( .A(n1596), .B(\register[1][6] ), .Y(n1523) );
  MXI2XL U195 ( .A(n2554), .B(n1536), .S0(n1621), .Y(n1539) );
  NOR2XL U196 ( .A(n1597), .B(\register[1][3] ), .Y(n1538) );
  MXI4XL U197 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n2172), .S1(n2146), 
        .Y(n1815) );
  MXI4XL U198 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n2160), .S1(n2137), 
        .Y(n1853) );
  MXI4XL U199 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n2168), .S1(n2143), .Y(
        n1749) );
  MXI4XL U200 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n1616), .S1(n1590), .Y(
        n1153) );
  NOR2BXL U201 ( .AN(n2146), .B(\register[3][7] ), .Y(n2066) );
  NOR2BXL U202 ( .AN(n1595), .B(\register[3][14] ), .Y(n1481) );
  NOR2BXL U203 ( .AN(n1595), .B(\register[3][9] ), .Y(n1506) );
  NOR2BXL U204 ( .AN(n1595), .B(\register[3][5] ), .Y(n1526) );
  NOR2BXL U205 ( .AN(n1595), .B(\register[3][7] ), .Y(n1516) );
  NOR2BXL U206 ( .AN(n1596), .B(\register[3][4] ), .Y(n1531) );
  NOR2BXL U207 ( .AN(n1596), .B(\register[3][6] ), .Y(n1521) );
  NOR2BXL U208 ( .AN(n1596), .B(\register[3][3] ), .Y(n1536) );
  MXI4XL U209 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n2172), .S1(n2146), .Y(
        n1754) );
  MXI4XL U210 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n2172), .S1(n2146), 
        .Y(n1814) );
  MXI4XL U211 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n2172), .S1(n2146), .Y(
        n1944) );
  MXI4XL U212 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n2168), .S1(n2143), .Y(
        n1746) );
  MXI4XL U213 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n2168), .S1(n2143), .Y(
        n1750) );
  MXI4XL U214 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n1616), .S1(n1590), .Y(
        n1152) );
  MXI4XL U215 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n1620), .S1(n1594), 
        .Y(n1256) );
  MXI4XL U216 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n1605), .S1(n1592), .Y(
        n1212) );
  MXI4XL U217 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n1616), .S1(n1591), .Y(
        n1164) );
  MXI4XL U218 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n2159), .S1(n2137), 
        .Y(n1850) );
  MXI4XL U219 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n1605), .S1(n1593), .Y(
        n1216) );
  MXI4XL U220 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n2160), .S1(n2137), 
        .Y(n1854) );
  MXI4XL U221 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n1620), .S1(n1594), 
        .Y(n1257) );
  MXI4XL U222 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n1605), .S1(n1593), .Y(
        n1215) );
  MXI4XL U223 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n1616), .S1(n1590), .Y(
        n1151) );
  MXI4XL U224 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n1620), .S1(n1594), 
        .Y(n1255) );
  MXI4XL U225 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n2168), .S1(n2143), .Y(
        n1748) );
  MXI4XL U226 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n1620), .S1(n1594), 
        .Y(n1254) );
  MXI4XL U227 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n2169), .S1(n2143), .Y(
        n1752) );
  MXI4XL U228 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n1616), .S1(n1590), .Y(
        n1154) );
  MXI4XL U229 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n1620), .S1(n1594), .Y(
        n1258) );
  MXI4XL U230 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n1605), .S1(n1593), .Y(
        n1214) );
  MXI4XL U231 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n1616), .S1(n1591), .Y(
        n1166) );
  MXI4XL U232 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n2160), .S1(n2137), 
        .Y(n1852) );
  MXI4XL U233 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n1618), .S1(n1593), .Y(
        n1218) );
  MXI4XL U234 ( .A(\register[4][7] ), .B(\register[5][7] ), .C(
        \register[6][7] ), .D(\register[7][7] ), .S0(n1605), .S1(n1592), .Y(
        n1202) );
  MXI4XL U235 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n2160), .S1(n2137), .Y(
        n1856) );
  MXI4XL U236 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n2168), .S1(n2143), .Y(
        n1747) );
  MXI4XL U237 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n1620), .S1(n1594), 
        .Y(n1253) );
  MXI4XL U238 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n2169), .S1(n2143), .Y(
        n1751) );
  MXI4XL U239 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n1605), .S1(n1593), .Y(
        n1213) );
  MXI4XL U240 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n1616), .S1(n1591), .Y(
        n1165) );
  MXI4XL U241 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n2159), .S1(n2137), 
        .Y(n1851) );
  MXI4XL U242 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n1615), .S1(n1590), .Y(
        n1149) );
  MXI4XL U243 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n1618), .S1(n1593), .Y(
        n1217) );
  MXI4XL U244 ( .A(\register[8][7] ), .B(\register[9][7] ), .C(
        \register[10][7] ), .D(\register[11][7] ), .S0(n1605), .S1(n1592), .Y(
        n1201) );
  MXI4XL U245 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n2160), .S1(n2137), 
        .Y(n1855) );
  NOR2X1 U246 ( .A(n2150), .B(n2175), .Y(n2022) );
  NOR2X1 U247 ( .A(n2150), .B(n2175), .Y(n2017) );
  NOR2X1 U248 ( .A(n2150), .B(n2175), .Y(n2007) );
  NOR2X1 U249 ( .A(n2151), .B(n2175), .Y(n2002) );
  NOR2X1 U250 ( .A(n2151), .B(n2175), .Y(n1997) );
  NOR2X1 U251 ( .A(n2151), .B(n2175), .Y(n1992) );
  NOR2X1 U252 ( .A(n2151), .B(n2175), .Y(n1987) );
  NOR2X1 U253 ( .A(n2151), .B(n2175), .Y(n1982) );
  NOR2X1 U254 ( .A(n1599), .B(n1623), .Y(n1472) );
  NOR2X1 U255 ( .A(n1599), .B(n1623), .Y(n1467) );
  NOR2X1 U256 ( .A(n1599), .B(n1623), .Y(n1457) );
  NOR2X1 U257 ( .A(n1600), .B(n1623), .Y(n1452) );
  NOR2X1 U258 ( .A(n1600), .B(n1623), .Y(n1447) );
  NOR2X1 U259 ( .A(n1600), .B(n1623), .Y(n1442) );
  NOR2X1 U260 ( .A(n1600), .B(n1623), .Y(n1437) );
  NOR2X1 U261 ( .A(n1600), .B(n1623), .Y(n1432) );
  NOR2X1 U262 ( .A(n2147), .B(n2177), .Y(n2102) );
  NOR2X1 U263 ( .A(n2147), .B(n2177), .Y(n2077) );
  NOR2X1 U264 ( .A(n2149), .B(n2177), .Y(n2097) );
  NOR2X1 U265 ( .A(n2148), .B(n2177), .Y(n2092) );
  NOR2X1 U266 ( .A(n2148), .B(n2177), .Y(n2087) );
  NOR2X1 U267 ( .A(n2148), .B(n2177), .Y(n2082) );
  NOR2X1 U268 ( .A(n2149), .B(n2177), .Y(n2072) );
  NOR2X1 U269 ( .A(n2148), .B(n2177), .Y(n2067) );
  NOR2X1 U270 ( .A(n2148), .B(n2176), .Y(n2062) );
  NOR2X1 U271 ( .A(n2148), .B(n2176), .Y(n2057) );
  NOR2X1 U272 ( .A(n2148), .B(n2176), .Y(n2052) );
  NOR2X1 U273 ( .A(n2149), .B(n2176), .Y(n2047) );
  NOR2X1 U274 ( .A(n2149), .B(n2176), .Y(n2042) );
  NOR2X1 U275 ( .A(n2149), .B(n2176), .Y(n2037) );
  NOR2X1 U276 ( .A(n2150), .B(n2176), .Y(n2032) );
  NOR2X1 U277 ( .A(n2150), .B(n2176), .Y(n2027) );
  NOR2X1 U278 ( .A(n2150), .B(n2176), .Y(n2012) );
  NOR2X1 U279 ( .A(n2151), .B(n2176), .Y(n1977) );
  NOR2X1 U280 ( .A(n1598), .B(n1625), .Y(n1547) );
  NOR2X1 U281 ( .A(n1597), .B(n1625), .Y(n1542) );
  NOR2X1 U282 ( .A(n1597), .B(n1624), .Y(n1512) );
  NOR2X1 U283 ( .A(n1597), .B(n1624), .Y(n1502) );
  NOR2X1 U284 ( .A(n1598), .B(n1624), .Y(n1497) );
  NOR2X1 U285 ( .A(n1598), .B(n1624), .Y(n1492) );
  NOR2X1 U286 ( .A(n1598), .B(n1624), .Y(n1487) );
  NOR2X1 U287 ( .A(n1599), .B(n1624), .Y(n1482) );
  NOR2X1 U288 ( .A(n1599), .B(n1624), .Y(n1477) );
  NOR2X1 U289 ( .A(n1599), .B(n1624), .Y(n1462) );
  NOR2X1 U290 ( .A(n1600), .B(n1624), .Y(n1427) );
  CLKBUFX3 U291 ( .A(n2276), .Y(n2197) );
  CLKBUFX3 U292 ( .A(n2276), .Y(n2198) );
  CLKBUFX3 U293 ( .A(n2276), .Y(n2199) );
  CLKBUFX3 U294 ( .A(n2276), .Y(n2200) );
  CLKBUFX3 U295 ( .A(n2277), .Y(n2193) );
  CLKBUFX3 U296 ( .A(n2277), .Y(n2194) );
  CLKBUFX3 U297 ( .A(n2277), .Y(n2195) );
  CLKBUFX3 U298 ( .A(n2277), .Y(n2196) );
  CLKBUFX3 U299 ( .A(n2278), .Y(n2189) );
  CLKBUFX3 U300 ( .A(n2278), .Y(n2190) );
  CLKBUFX3 U301 ( .A(n2278), .Y(n2191) );
  CLKBUFX3 U302 ( .A(n2278), .Y(n2192) );
  CLKBUFX3 U303 ( .A(n2273), .Y(n2209) );
  CLKBUFX3 U304 ( .A(n2273), .Y(n2210) );
  CLKBUFX3 U305 ( .A(n2273), .Y(n2211) );
  CLKBUFX3 U306 ( .A(n2273), .Y(n2212) );
  CLKBUFX3 U307 ( .A(n2274), .Y(n2205) );
  CLKBUFX3 U308 ( .A(n2274), .Y(n2206) );
  CLKBUFX3 U309 ( .A(n2274), .Y(n2207) );
  CLKBUFX3 U310 ( .A(n2274), .Y(n2208) );
  CLKBUFX3 U311 ( .A(n2275), .Y(n2201) );
  CLKBUFX3 U312 ( .A(n2275), .Y(n2202) );
  CLKBUFX3 U313 ( .A(n2275), .Y(n2203) );
  CLKBUFX3 U314 ( .A(n2275), .Y(n2204) );
  CLKBUFX3 U315 ( .A(n2270), .Y(n2221) );
  CLKBUFX3 U316 ( .A(n2270), .Y(n2222) );
  CLKBUFX3 U317 ( .A(n2270), .Y(n2223) );
  CLKBUFX3 U318 ( .A(n2270), .Y(n2224) );
  CLKBUFX3 U319 ( .A(n2271), .Y(n2217) );
  CLKBUFX3 U320 ( .A(n2271), .Y(n2218) );
  CLKBUFX3 U321 ( .A(n2271), .Y(n2219) );
  CLKBUFX3 U322 ( .A(n2271), .Y(n2220) );
  CLKBUFX3 U323 ( .A(n2272), .Y(n2213) );
  CLKBUFX3 U324 ( .A(n2272), .Y(n2214) );
  CLKBUFX3 U325 ( .A(n2272), .Y(n2215) );
  CLKBUFX3 U326 ( .A(n2272), .Y(n2216) );
  CLKBUFX3 U327 ( .A(n2267), .Y(n2233) );
  CLKBUFX3 U328 ( .A(n2267), .Y(n2234) );
  CLKBUFX3 U329 ( .A(n2267), .Y(n2235) );
  CLKBUFX3 U330 ( .A(n2267), .Y(n2236) );
  CLKBUFX3 U331 ( .A(n2268), .Y(n2229) );
  CLKBUFX3 U332 ( .A(n2268), .Y(n2230) );
  CLKBUFX3 U333 ( .A(n2268), .Y(n2231) );
  CLKBUFX3 U334 ( .A(n2268), .Y(n2232) );
  CLKBUFX3 U335 ( .A(n2269), .Y(n2225) );
  CLKBUFX3 U336 ( .A(n2269), .Y(n2226) );
  CLKBUFX3 U337 ( .A(n2269), .Y(n2227) );
  CLKBUFX3 U338 ( .A(n2269), .Y(n2228) );
  CLKBUFX3 U339 ( .A(n2264), .Y(n2245) );
  CLKBUFX3 U340 ( .A(n2264), .Y(n2246) );
  CLKBUFX3 U341 ( .A(n2264), .Y(n2247) );
  CLKBUFX3 U342 ( .A(n2264), .Y(n2248) );
  CLKBUFX3 U343 ( .A(n2265), .Y(n2241) );
  CLKBUFX3 U344 ( .A(n2265), .Y(n2242) );
  CLKBUFX3 U345 ( .A(n2265), .Y(n2243) );
  CLKBUFX3 U346 ( .A(n2265), .Y(n2244) );
  CLKBUFX3 U347 ( .A(n2266), .Y(n2237) );
  CLKBUFX3 U348 ( .A(n2266), .Y(n2238) );
  CLKBUFX3 U349 ( .A(n2266), .Y(n2239) );
  CLKBUFX3 U350 ( .A(n2266), .Y(n2240) );
  CLKBUFX3 U351 ( .A(n2261), .Y(n2257) );
  CLKBUFX3 U352 ( .A(n2261), .Y(n2258) );
  CLKBUFX3 U353 ( .A(n2261), .Y(n2259) );
  CLKBUFX3 U354 ( .A(n2262), .Y(n2253) );
  CLKBUFX3 U355 ( .A(n2262), .Y(n2254) );
  CLKBUFX3 U356 ( .A(n2262), .Y(n2256) );
  CLKBUFX3 U357 ( .A(n2262), .Y(n2255) );
  CLKBUFX3 U358 ( .A(n2263), .Y(n2249) );
  CLKBUFX3 U359 ( .A(n2263), .Y(n2250) );
  CLKBUFX3 U360 ( .A(n2263), .Y(n2251) );
  CLKBUFX3 U361 ( .A(n2263), .Y(n2252) );
  CLKBUFX3 U362 ( .A(n2261), .Y(n2260) );
  CLKBUFX3 U363 ( .A(n2132), .Y(n2146) );
  CLKBUFX3 U364 ( .A(n1576), .Y(n1595) );
  CLKBUFX3 U365 ( .A(n2156), .Y(n2173) );
  CLKBUFX3 U366 ( .A(n2155), .Y(n2174) );
  CLKBUFX3 U367 ( .A(n1606), .Y(n1621) );
  CLKBUFX3 U368 ( .A(n1604), .Y(n1622) );
  NOR2X1 U369 ( .A(n2129), .B(n2176), .Y(n1972) );
  NOR2X1 U370 ( .A(n2129), .B(n2176), .Y(n1967) );
  NOR2X1 U371 ( .A(n2129), .B(n2177), .Y(n1962) );
  NOR2X1 U372 ( .A(n2129), .B(n2177), .Y(n1957) );
  NOR2X1 U373 ( .A(n2129), .B(n2177), .Y(n1952) );
  NOR2X1 U374 ( .A(n2137), .B(n2177), .Y(n1947) );
  NOR2X1 U375 ( .A(n1578), .B(n1624), .Y(n1417) );
  NOR2X1 U376 ( .A(n1578), .B(n1625), .Y(n1412) );
  NOR2X1 U377 ( .A(n1578), .B(n1625), .Y(n1407) );
  NOR2X1 U378 ( .A(n1594), .B(n1625), .Y(n1402) );
  NOR2X1 U379 ( .A(n1578), .B(n1625), .Y(n1397) );
  CLKBUFX3 U380 ( .A(n2153), .Y(n2166) );
  CLKBUFX3 U381 ( .A(n2153), .Y(n2167) );
  CLKBUFX3 U382 ( .A(n2153), .Y(n2168) );
  CLKBUFX3 U383 ( .A(n2157), .Y(n2170) );
  CLKBUFX3 U384 ( .A(n2157), .Y(n2171) );
  CLKBUFX3 U385 ( .A(n2153), .Y(n2169) );
  CLKBUFX3 U386 ( .A(n2152), .Y(n2158) );
  CLKBUFX3 U387 ( .A(n2152), .Y(n2159) );
  CLKBUFX3 U388 ( .A(n2152), .Y(n2160) );
  CLKBUFX3 U389 ( .A(n2154), .Y(n2162) );
  CLKBUFX3 U390 ( .A(n2154), .Y(n2163) );
  CLKBUFX3 U391 ( .A(n2155), .Y(n2164) );
  CLKBUFX3 U392 ( .A(n2544), .Y(n2161) );
  CLKBUFX3 U393 ( .A(n2155), .Y(n2165) );
  CLKBUFX3 U394 ( .A(n1607), .Y(n1616) );
  CLKBUFX3 U395 ( .A(n1607), .Y(n1617) );
  CLKBUFX3 U396 ( .A(n1603), .Y(n1618) );
  CLKBUFX3 U397 ( .A(n1603), .Y(n1619) );
  CLKBUFX3 U398 ( .A(n1601), .Y(n1608) );
  CLKBUFX3 U399 ( .A(n1601), .Y(n1609) );
  CLKBUFX3 U400 ( .A(n2546), .Y(n1610) );
  CLKBUFX3 U401 ( .A(n1602), .Y(n1612) );
  CLKBUFX3 U402 ( .A(n1603), .Y(n1613) );
  CLKBUFX3 U403 ( .A(n1604), .Y(n1614) );
  CLKBUFX3 U404 ( .A(n2546), .Y(n1611) );
  CLKBUFX3 U405 ( .A(n1603), .Y(n1615) );
  BUFX4 U406 ( .A(n2133), .Y(n2142) );
  BUFX4 U407 ( .A(n2133), .Y(n2144) );
  BUFX4 U408 ( .A(n2133), .Y(n2145) );
  BUFX4 U409 ( .A(n2133), .Y(n2136) );
  BUFX4 U410 ( .A(n2126), .Y(n2137) );
  BUFX4 U411 ( .A(n2135), .Y(n2139) );
  BUFX4 U412 ( .A(n2134), .Y(n2141) );
  BUFX4 U413 ( .A(n2135), .Y(n2138) );
  BUFX4 U414 ( .A(n2134), .Y(n2140) );
  BUFX4 U415 ( .A(n1581), .Y(n1591) );
  BUFX4 U416 ( .A(n1581), .Y(n1593) );
  BUFX4 U417 ( .A(n1575), .Y(n1594) );
  BUFX4 U418 ( .A(n1581), .Y(n1592) );
  BUFX4 U419 ( .A(n1584), .Y(n1585) );
  BUFX4 U420 ( .A(n1584), .Y(n1586) );
  BUFX4 U421 ( .A(n1583), .Y(n1588) );
  BUFX4 U422 ( .A(n1582), .Y(n1590) );
  BUFX4 U423 ( .A(n1583), .Y(n1587) );
  BUFX4 U424 ( .A(n1582), .Y(n1589) );
  CLKBUFX3 U425 ( .A(n2132), .Y(n2147) );
  CLKBUFX3 U426 ( .A(n1576), .Y(n1596) );
  CLKBUFX3 U427 ( .A(n2131), .Y(n2148) );
  CLKBUFX3 U428 ( .A(n2131), .Y(n2149) );
  CLKBUFX3 U429 ( .A(n2130), .Y(n2151) );
  CLKBUFX3 U430 ( .A(n1580), .Y(n1597) );
  CLKBUFX3 U431 ( .A(n1580), .Y(n1598) );
  CLKBUFX3 U432 ( .A(n1579), .Y(n1600) );
  CLKBUFX3 U433 ( .A(n2279), .Y(n2186) );
  CLKBUFX3 U434 ( .A(n2279), .Y(n2187) );
  CLKBUFX3 U435 ( .A(n2279), .Y(n2188) );
  CLKBUFX3 U436 ( .A(n2280), .Y(n2182) );
  CLKBUFX3 U437 ( .A(n2280), .Y(n2183) );
  CLKBUFX3 U438 ( .A(n2280), .Y(n2184) );
  CLKBUFX3 U439 ( .A(n2279), .Y(n2185) );
  CLKBUFX3 U440 ( .A(n2280), .Y(n2181) );
  CLKBUFX3 U441 ( .A(n2281), .Y(n2178) );
  CLKBUFX3 U442 ( .A(n2281), .Y(n2179) );
  CLKBUFX3 U443 ( .A(n2289), .Y(n2180) );
  CLKBUFX3 U444 ( .A(n2282), .Y(n2276) );
  CLKBUFX3 U445 ( .A(n2282), .Y(n2277) );
  CLKBUFX3 U446 ( .A(n2282), .Y(n2278) );
  CLKBUFX3 U447 ( .A(n2283), .Y(n2273) );
  CLKBUFX3 U448 ( .A(n2283), .Y(n2274) );
  CLKBUFX3 U449 ( .A(n2283), .Y(n2275) );
  CLKBUFX3 U450 ( .A(n2284), .Y(n2270) );
  CLKBUFX3 U451 ( .A(n2284), .Y(n2271) );
  CLKBUFX3 U452 ( .A(n2284), .Y(n2272) );
  CLKBUFX3 U453 ( .A(n2285), .Y(n2267) );
  CLKBUFX3 U454 ( .A(n2285), .Y(n2268) );
  CLKBUFX3 U455 ( .A(n2285), .Y(n2269) );
  CLKBUFX3 U456 ( .A(n2286), .Y(n2264) );
  CLKBUFX3 U457 ( .A(n2286), .Y(n2265) );
  CLKBUFX3 U458 ( .A(n2286), .Y(n2266) );
  CLKBUFX3 U459 ( .A(n2287), .Y(n2261) );
  CLKBUFX3 U460 ( .A(n2287), .Y(n2262) );
  CLKBUFX3 U461 ( .A(n2287), .Y(n2263) );
  CLKBUFX3 U462 ( .A(n101), .Y(n2400) );
  CLKBUFX3 U463 ( .A(n103), .Y(n2388) );
  CLKBUFX3 U464 ( .A(n2396), .Y(n2398) );
  CLKBUFX3 U465 ( .A(n2396), .Y(n2399) );
  CLKBUFX3 U466 ( .A(n103), .Y(n2387) );
  CLKBUFX3 U467 ( .A(n2116), .Y(n2113) );
  CLKBUFX3 U468 ( .A(n2116), .Y(n2114) );
  CLKBUFX3 U469 ( .A(n2116), .Y(n2115) );
  CLKBUFX3 U470 ( .A(n1567), .Y(n1563) );
  CLKBUFX3 U471 ( .A(n1567), .Y(n1564) );
  CLKBUFX3 U472 ( .A(n1567), .Y(n1565) );
  CLKBUFX3 U473 ( .A(n2549), .Y(n1566) );
  CLKBUFX3 U474 ( .A(n1577), .Y(n1578) );
  CLKBUFX3 U475 ( .A(n2365), .Y(n2368) );
  CLKBUFX3 U476 ( .A(n2376), .Y(n2379) );
  CLKBUFX3 U477 ( .A(n101), .Y(n2401) );
  CLKBUFX3 U478 ( .A(n103), .Y(n2389) );
  CLKBUFX3 U479 ( .A(n2365), .Y(n2369) );
  CLKBUFX3 U480 ( .A(n2376), .Y(n2380) );
  CLKBUFX3 U481 ( .A(n2364), .Y(n2366) );
  CLKBUFX3 U482 ( .A(n2364), .Y(n2367) );
  CLKBUFX3 U483 ( .A(n2376), .Y(n2377) );
  CLKBUFX3 U484 ( .A(n2376), .Y(n2378) );
  CLKBUFX3 U485 ( .A(n2117), .Y(n2121) );
  CLKBUFX3 U486 ( .A(n2117), .Y(n2122) );
  CLKBUFX3 U487 ( .A(n2118), .Y(n2123) );
  CLKBUFX3 U488 ( .A(n2117), .Y(n2124) );
  CLKBUFX3 U489 ( .A(n2548), .Y(n1570) );
  CLKBUFX3 U490 ( .A(n1574), .Y(n1571) );
  CLKBUFX3 U491 ( .A(n1574), .Y(n1572) );
  CLKBUFX3 U492 ( .A(n2548), .Y(n1573) );
  CLKBUFX3 U493 ( .A(n2128), .Y(n2131) );
  CLKBUFX3 U494 ( .A(n2128), .Y(n2130) );
  CLKBUFX3 U495 ( .A(n1577), .Y(n1580) );
  CLKBUFX3 U496 ( .A(n1577), .Y(n1579) );
  CLKBUFX3 U497 ( .A(n2127), .Y(n2133) );
  CLKBUFX3 U498 ( .A(n2126), .Y(n2135) );
  CLKBUFX3 U499 ( .A(n2126), .Y(n2134) );
  CLKBUFX3 U500 ( .A(n1575), .Y(n1584) );
  CLKBUFX3 U501 ( .A(n1575), .Y(n1583) );
  CLKBUFX3 U502 ( .A(n1575), .Y(n1582) );
  CLKBUFX3 U503 ( .A(n2154), .Y(n2156) );
  CLKBUFX3 U504 ( .A(n1603), .Y(n1606) );
  CLKBUFX3 U505 ( .A(n2288), .Y(n2282) );
  CLKBUFX3 U506 ( .A(n2288), .Y(n2283) );
  CLKBUFX3 U507 ( .A(n2289), .Y(n2284) );
  CLKBUFX3 U508 ( .A(n2288), .Y(n2285) );
  CLKBUFX3 U509 ( .A(n2289), .Y(n2286) );
  CLKBUFX3 U510 ( .A(n2288), .Y(n2287) );
  CLKBUFX3 U511 ( .A(n2281), .Y(n2279) );
  CLKBUFX3 U512 ( .A(n2281), .Y(n2280) );
  CLKBUFX3 U513 ( .A(n65), .Y(n2531) );
  CLKBUFX3 U514 ( .A(n70), .Y(n2519) );
  CLKBUFX3 U515 ( .A(n2487), .Y(n2490) );
  CLKBUFX3 U516 ( .A(n92), .Y(n2444) );
  CLKBUFX3 U517 ( .A(n2475), .Y(n2478) );
  CLKBUFX3 U518 ( .A(n94), .Y(n2432) );
  CLKBUFX3 U519 ( .A(n2527), .Y(n2529) );
  CLKBUFX3 U520 ( .A(n2527), .Y(n2530) );
  CLKBUFX3 U521 ( .A(n70), .Y(n2518) );
  CLKBUFX3 U522 ( .A(n2487), .Y(n2488) );
  CLKBUFX3 U523 ( .A(n2487), .Y(n2489) );
  CLKBUFX3 U524 ( .A(n2440), .Y(n2442) );
  CLKBUFX3 U525 ( .A(n2440), .Y(n2443) );
  CLKBUFX3 U526 ( .A(n2475), .Y(n2476) );
  CLKBUFX3 U527 ( .A(n2475), .Y(n2477) );
  CLKBUFX3 U528 ( .A(n2428), .Y(n2430) );
  CLKBUFX3 U529 ( .A(n2428), .Y(n2431) );
  CLKBUFX3 U530 ( .A(n101), .Y(n2396) );
  CLKBUFX3 U531 ( .A(n2539), .Y(n2542) );
  CLKBUFX3 U532 ( .A(n2109), .Y(n2107) );
  CLKBUFX3 U533 ( .A(n2109), .Y(n2108) );
  CLKBUFX3 U534 ( .A(n1559), .Y(n1557) );
  CLKBUFX3 U535 ( .A(n1559), .Y(n1558) );
  CLKBUFX3 U536 ( .A(n72), .Y(n2515) );
  CLKBUFX3 U537 ( .A(n76), .Y(n2506) );
  CLKBUFX3 U538 ( .A(n86), .Y(n2471) );
  CLKBUFX3 U539 ( .A(n2457), .Y(n2461) );
  CLKBUFX3 U540 ( .A(n95), .Y(n2426) );
  CLKBUFX3 U541 ( .A(n2412), .Y(n2416) );
  CLKBUFX3 U542 ( .A(n104), .Y(n2383) );
  CLKBUFX3 U543 ( .A(n2370), .Y(n2374) );
  CLKBUFX3 U544 ( .A(n68), .Y(n2525) );
  CLKBUFX3 U545 ( .A(n84), .Y(n2484) );
  CLKBUFX3 U546 ( .A(n93), .Y(n2438) );
  CLKBUFX3 U547 ( .A(n102), .Y(n2394) );
  CLKBUFX3 U548 ( .A(n2497), .Y(n2500) );
  CLKBUFX3 U549 ( .A(n2452), .Y(n2455) );
  CLKBUFX3 U550 ( .A(n10), .Y(n2409) );
  CLKBUFX3 U551 ( .A(n2508), .Y(n2511) );
  CLKBUFX3 U552 ( .A(n80), .Y(n2494) );
  CLKBUFX3 U553 ( .A(n90), .Y(n2449) );
  CLKBUFX3 U554 ( .A(n99), .Y(n2404) );
  CLKBUFX3 U555 ( .A(n2464), .Y(n2467) );
  CLKBUFX3 U556 ( .A(n8), .Y(n2421) );
  CLKBUFX3 U557 ( .A(n2534), .Y(n2537) );
  CLKBUFX3 U558 ( .A(n2539), .Y(n2541) );
  CLKBUFX3 U559 ( .A(n47), .Y(n2540) );
  CLKBUFX3 U560 ( .A(n65), .Y(n2532) );
  CLKBUFX3 U561 ( .A(n70), .Y(n2520) );
  CLKBUFX3 U562 ( .A(n2487), .Y(n2491) );
  CLKBUFX3 U563 ( .A(n92), .Y(n2445) );
  CLKBUFX3 U564 ( .A(n2475), .Y(n2479) );
  CLKBUFX3 U565 ( .A(n94), .Y(n2433) );
  CLKBUFX3 U566 ( .A(n72), .Y(n2516) );
  CLKBUFX3 U567 ( .A(n76), .Y(n2507) );
  CLKBUFX3 U568 ( .A(n86), .Y(n2472) );
  CLKBUFX3 U569 ( .A(n2457), .Y(n2462) );
  CLKBUFX3 U570 ( .A(n95), .Y(n2427) );
  CLKBUFX3 U571 ( .A(n2412), .Y(n2417) );
  CLKBUFX3 U572 ( .A(n104), .Y(n2384) );
  CLKBUFX3 U573 ( .A(n2370), .Y(n2375) );
  CLKBUFX3 U574 ( .A(n68), .Y(n2526) );
  CLKBUFX3 U575 ( .A(n84), .Y(n2485) );
  CLKBUFX3 U576 ( .A(n93), .Y(n2439) );
  CLKBUFX3 U577 ( .A(n102), .Y(n2395) );
  CLKBUFX3 U578 ( .A(n2497), .Y(n2501) );
  CLKBUFX3 U579 ( .A(n2452), .Y(n2456) );
  CLKBUFX3 U580 ( .A(n10), .Y(n2410) );
  CLKBUFX3 U581 ( .A(n2464), .Y(n2468) );
  CLKBUFX3 U582 ( .A(n8), .Y(n2422) );
  CLKBUFX3 U583 ( .A(n2508), .Y(n2512) );
  CLKBUFX3 U584 ( .A(n80), .Y(n2495) );
  CLKBUFX3 U585 ( .A(n90), .Y(n2450) );
  CLKBUFX3 U586 ( .A(n99), .Y(n2405) );
  CLKBUFX3 U587 ( .A(n72), .Y(n2514) );
  CLKBUFX3 U588 ( .A(n2502), .Y(n2504) );
  CLKBUFX3 U589 ( .A(n2502), .Y(n2505) );
  CLKBUFX3 U590 ( .A(n86), .Y(n2469) );
  CLKBUFX3 U591 ( .A(n86), .Y(n2470) );
  CLKBUFX3 U592 ( .A(n2458), .Y(n2459) );
  CLKBUFX3 U593 ( .A(n88), .Y(n2460) );
  CLKBUFX3 U594 ( .A(n95), .Y(n2425) );
  CLKBUFX3 U595 ( .A(n2413), .Y(n2414) );
  CLKBUFX3 U596 ( .A(n97), .Y(n2415) );
  CLKBUFX3 U597 ( .A(n104), .Y(n2381) );
  CLKBUFX3 U598 ( .A(n104), .Y(n2382) );
  CLKBUFX3 U599 ( .A(n2371), .Y(n2372) );
  CLKBUFX3 U600 ( .A(n106), .Y(n2373) );
  CLKBUFX3 U601 ( .A(n2521), .Y(n2523) );
  CLKBUFX3 U602 ( .A(n2521), .Y(n2524) );
  CLKBUFX3 U603 ( .A(n2480), .Y(n2482) );
  CLKBUFX3 U604 ( .A(n2480), .Y(n2483) );
  CLKBUFX3 U605 ( .A(n2434), .Y(n2436) );
  CLKBUFX3 U606 ( .A(n2434), .Y(n2437) );
  CLKBUFX3 U607 ( .A(n2390), .Y(n2392) );
  CLKBUFX3 U608 ( .A(n2390), .Y(n2393) );
  CLKBUFX3 U609 ( .A(n2496), .Y(n2498) );
  CLKBUFX3 U610 ( .A(n2496), .Y(n2499) );
  CLKBUFX3 U611 ( .A(n2451), .Y(n2453) );
  CLKBUFX3 U612 ( .A(n2451), .Y(n2454) );
  CLKBUFX3 U613 ( .A(n2406), .Y(n2407) );
  CLKBUFX3 U614 ( .A(n2406), .Y(n2408) );
  CLKBUFX3 U615 ( .A(n2508), .Y(n2509) );
  CLKBUFX3 U616 ( .A(n2508), .Y(n2510) );
  CLKBUFX3 U617 ( .A(n80), .Y(n2492) );
  CLKBUFX3 U618 ( .A(n80), .Y(n2493) );
  CLKBUFX3 U619 ( .A(n90), .Y(n2447) );
  CLKBUFX3 U620 ( .A(n90), .Y(n2448) );
  CLKBUFX3 U621 ( .A(n99), .Y(n2402) );
  CLKBUFX3 U622 ( .A(n99), .Y(n2403) );
  CLKBUFX3 U623 ( .A(n2463), .Y(n2465) );
  CLKBUFX3 U624 ( .A(n2463), .Y(n2466) );
  CLKBUFX3 U625 ( .A(n2418), .Y(n2419) );
  CLKBUFX3 U626 ( .A(n2418), .Y(n2420) );
  CLKBUFX3 U627 ( .A(N17), .Y(n2152) );
  CLKBUFX3 U628 ( .A(N12), .Y(n1601) );
  CLKBUFX3 U629 ( .A(N17), .Y(n2153) );
  CLKBUFX3 U630 ( .A(N12), .Y(n1602) );
  CLKBUFX3 U631 ( .A(N17), .Y(n2154) );
  CLKBUFX3 U632 ( .A(N12), .Y(n1603) );
  CLKBUFX3 U633 ( .A(N17), .Y(n2155) );
  CLKBUFX3 U634 ( .A(N12), .Y(n1604) );
  CLKBUFX3 U635 ( .A(n2545), .Y(n2128) );
  CLKBUFX3 U636 ( .A(n2547), .Y(n1577) );
  CLKBUFX3 U637 ( .A(n2545), .Y(n2126) );
  CLKBUFX3 U638 ( .A(n2547), .Y(n1575) );
  CLKBUFX3 U639 ( .A(n2116), .Y(n2110) );
  CLKBUFX3 U640 ( .A(n1567), .Y(n1560) );
  CLKBUFX3 U641 ( .A(n3), .Y(n2365) );
  CLKBUFX3 U642 ( .A(n2289), .Y(n2281) );
  CLKBUFX3 U643 ( .A(n65), .Y(n2527) );
  CLKBUFX3 U644 ( .A(n92), .Y(n2440) );
  CLKBUFX3 U645 ( .A(n94), .Y(n2428) );
  CLKBUFX3 U646 ( .A(n2610), .Y(n2354) );
  CLKBUFX3 U647 ( .A(n2609), .Y(n2351) );
  CLKBUFX3 U648 ( .A(n2589), .Y(n2303) );
  CLKBUFX3 U649 ( .A(n2610), .Y(n2353) );
  CLKBUFX3 U650 ( .A(n2613), .Y(n2361) );
  CLKBUFX3 U651 ( .A(n2612), .Y(n2359) );
  CLKBUFX3 U652 ( .A(n2608), .Y(n2349) );
  CLKBUFX3 U653 ( .A(n2593), .Y(n2312) );
  CLKBUFX3 U654 ( .A(n2588), .Y(n2301) );
  CLKBUFX3 U655 ( .A(n2586), .Y(n2296) );
  CLKBUFX3 U656 ( .A(n2613), .Y(n2360) );
  CLKBUFX3 U657 ( .A(n2612), .Y(n2358) );
  CLKBUFX3 U658 ( .A(n2608), .Y(n2348) );
  CLKBUFX3 U659 ( .A(n2607), .Y(n2346) );
  CLKBUFX3 U660 ( .A(n2606), .Y(n2344) );
  CLKBUFX3 U661 ( .A(n2602), .Y(n2335) );
  CLKBUFX3 U662 ( .A(n2601), .Y(n2332) );
  CLKBUFX3 U663 ( .A(n2600), .Y(n2330) );
  CLKBUFX3 U664 ( .A(n2599), .Y(n2327) );
  CLKBUFX3 U665 ( .A(n2598), .Y(n2324) );
  CLKBUFX3 U666 ( .A(n2591), .Y(n2307) );
  CLKBUFX3 U667 ( .A(n2590), .Y(n2305) );
  CLKBUFX3 U668 ( .A(n2595), .Y(n2316) );
  CLKBUFX3 U669 ( .A(n2587), .Y(n2299) );
  CLKBUFX3 U670 ( .A(n2602), .Y(n2334) );
  CLKBUFX3 U671 ( .A(n2600), .Y(n2329) );
  CLKBUFX3 U672 ( .A(n2599), .Y(n2326) );
  CLKBUFX3 U673 ( .A(n2611), .Y(n2356) );
  CLKBUFX3 U674 ( .A(n2605), .Y(n2342) );
  CLKBUFX3 U675 ( .A(n2604), .Y(n2339) );
  CLKBUFX3 U676 ( .A(n2603), .Y(n2337) );
  CLKBUFX3 U677 ( .A(n2597), .Y(n2322) );
  CLKBUFX3 U678 ( .A(n2596), .Y(n2319) );
  CLKBUFX3 U679 ( .A(n2594), .Y(n2314) );
  CLKBUFX3 U680 ( .A(n2592), .Y(n2310) );
  CLKBUFX3 U681 ( .A(n2585), .Y(n2294) );
  CLKBUFX3 U682 ( .A(n2584), .Y(n2292) );
  CLKBUFX3 U683 ( .A(n2597), .Y(n2321) );
  CLKBUFX3 U684 ( .A(n2596), .Y(n2318) );
  CLKBUFX3 U685 ( .A(n2592), .Y(n2309) );
  CLKBUFX3 U686 ( .A(n2587), .Y(n2298) );
  CLKBUFX3 U687 ( .A(n2583), .Y(n2290) );
  CLKBUFX3 U688 ( .A(n2611), .Y(n2355) );
  CLKBUFX3 U689 ( .A(n2605), .Y(n2341) );
  CLKBUFX3 U690 ( .A(n2614), .Y(n2362) );
  CLKBUFX3 U691 ( .A(n2609), .Y(n2352) );
  CLKBUFX3 U692 ( .A(n2589), .Y(n2304) );
  CLKBUFX3 U693 ( .A(n2593), .Y(n2313) );
  CLKBUFX3 U694 ( .A(n2588), .Y(n2302) );
  CLKBUFX3 U695 ( .A(n2586), .Y(n2297) );
  CLKBUFX3 U696 ( .A(n2598), .Y(n2325) );
  CLKBUFX3 U697 ( .A(n2591), .Y(n2308) );
  CLKBUFX3 U698 ( .A(n2590), .Y(n2306) );
  CLKBUFX3 U699 ( .A(n2607), .Y(n2347) );
  CLKBUFX3 U700 ( .A(n2606), .Y(n2345) );
  CLKBUFX3 U701 ( .A(n2602), .Y(n2336) );
  CLKBUFX3 U702 ( .A(n2601), .Y(n2333) );
  CLKBUFX3 U703 ( .A(n2600), .Y(n2331) );
  CLKBUFX3 U704 ( .A(n2599), .Y(n2328) );
  CLKBUFX3 U705 ( .A(n2596), .Y(n2320) );
  CLKBUFX3 U706 ( .A(n2595), .Y(n2317) );
  CLKBUFX3 U707 ( .A(n2592), .Y(n2311) );
  CLKBUFX3 U708 ( .A(n2587), .Y(n2300) );
  CLKBUFX3 U709 ( .A(n2611), .Y(n2357) );
  CLKBUFX3 U710 ( .A(n2603), .Y(n2338) );
  CLKBUFX3 U711 ( .A(n2597), .Y(n2323) );
  CLKBUFX3 U712 ( .A(n2594), .Y(n2315) );
  CLKBUFX3 U713 ( .A(n2585), .Y(n2295) );
  CLKBUFX3 U714 ( .A(n2584), .Y(n2293) );
  CLKBUFX3 U715 ( .A(n2605), .Y(n2343) );
  CLKBUFX3 U716 ( .A(n2604), .Y(n2340) );
  CLKBUFX3 U717 ( .A(n2583), .Y(n2291) );
  CLKBUFX3 U718 ( .A(n2614), .Y(n2363) );
  CLKBUFX3 U719 ( .A(n2109), .Y(n2106) );
  CLKBUFX3 U720 ( .A(n1559), .Y(n1556) );
  CLKBUFX3 U721 ( .A(n47), .Y(n2539) );
  CLKBUFX3 U722 ( .A(n56), .Y(n2533) );
  CLKBUFX3 U723 ( .A(n56), .Y(n2534) );
  CLKBUFX3 U724 ( .A(n5), .Y(n2497) );
  CLKBUFX3 U725 ( .A(n9), .Y(n2452) );
  CLKBUFX3 U726 ( .A(n7), .Y(n2464) );
  CLKBUFX3 U727 ( .A(n68), .Y(n2521) );
  CLKBUFX3 U728 ( .A(n84), .Y(n2480) );
  CLKBUFX3 U729 ( .A(n93), .Y(n2434) );
  CLKBUFX3 U730 ( .A(n102), .Y(n2390) );
  CLKBUFX3 U731 ( .A(n76), .Y(n2502) );
  CLKBUFX3 U732 ( .A(n88), .Y(n2457) );
  CLKBUFX3 U733 ( .A(n97), .Y(n2412) );
  CLKBUFX3 U734 ( .A(n106), .Y(n2370) );
  CLKBUFX3 U735 ( .A(n2406), .Y(n2411) );
  CLKBUFX3 U736 ( .A(n2418), .Y(n2423) );
  CLKBUFX3 U737 ( .A(n68), .Y(n2522) );
  CLKBUFX3 U738 ( .A(n93), .Y(n2435) );
  CLKBUFX3 U739 ( .A(n65), .Y(n2528) );
  CLKBUFX3 U740 ( .A(n76), .Y(n2503) );
  CLKBUFX3 U741 ( .A(n92), .Y(n2441) );
  CLKBUFX3 U742 ( .A(n94), .Y(n2429) );
  CLKBUFX3 U743 ( .A(n86), .Y(n2473) );
  CLKBUFX3 U744 ( .A(n104), .Y(n2385) );
  AND2XL U745 ( .A(n66), .B(n2), .Y(n13) );
  BUFX4 U746 ( .A(n83), .Y(n2487) );
  NAND2XL U747 ( .A(n81), .B(n66), .Y(n83) );
  BUFX4 U748 ( .A(n85), .Y(n2475) );
  NAND2XL U749 ( .A(n81), .B(n71), .Y(n85) );
  AND2XL U750 ( .A(n91), .B(n77), .Y(n18) );
  AND2XL U751 ( .A(n100), .B(n77), .Y(n19) );
  NOR3X1 U752 ( .A(n2618), .B(n2619), .C(n2617), .Y(n79) );
  XNOR2X1 U753 ( .A(n2616), .B(N20), .Y(n54) );
  XNOR2X1 U754 ( .A(n2615), .B(N21), .Y(n53) );
  AND2XL U755 ( .A(n81), .B(n69), .Y(n26) );
  AND2XL U756 ( .A(n91), .B(n69), .Y(n27) );
  INVX3 U757 ( .A(n29), .Y(n80) );
  INVX3 U758 ( .A(n30), .Y(n90) );
  INVX3 U759 ( .A(n31), .Y(n99) );
  CLKBUFX3 U760 ( .A(N15), .Y(n2549) );
  CLKBUFX3 U761 ( .A(N14), .Y(n2548) );
  CLKBUFX3 U762 ( .A(N13), .Y(n2547) );
  OAI2BB2XL U763 ( .B0(n2308), .B1(n2531), .A0N(\register[1][23] ), .A1N(n2531), .Y(n131) );
  OAI2BB2XL U764 ( .B0(n2304), .B1(n2531), .A0N(\register[1][25] ), .A1N(n2532), .Y(n133) );
  OAI2BB2XL U765 ( .B0(n2302), .B1(n2531), .A0N(\register[1][26] ), .A1N(n2532), .Y(n134) );
  OAI2BB2XL U766 ( .B0(n2300), .B1(n2531), .A0N(\register[1][27] ), .A1N(n2532), .Y(n135) );
  OAI2BB2XL U767 ( .B0(n2297), .B1(n2531), .A0N(\register[1][28] ), .A1N(n2532), .Y(n136) );
  OAI2BB2XL U768 ( .B0(n2295), .B1(n2531), .A0N(\register[1][29] ), .A1N(n2532), .Y(n137) );
  OAI2BB2XL U769 ( .B0(n2293), .B1(n2531), .A0N(\register[1][30] ), .A1N(n2528), .Y(n138) );
  OAI2BB2XL U770 ( .B0(n2291), .B1(n2531), .A0N(\register[1][31] ), .A1N(n2528), .Y(n139) );
  OAI2BB2XL U771 ( .B0(n2308), .B1(n2519), .A0N(\register[3][23] ), .A1N(n2519), .Y(n195) );
  OAI2BB2XL U772 ( .B0(n2304), .B1(n2519), .A0N(\register[3][25] ), .A1N(n2520), .Y(n197) );
  OAI2BB2XL U773 ( .B0(n2302), .B1(n2519), .A0N(\register[3][26] ), .A1N(n2520), .Y(n198) );
  OAI2BB2XL U774 ( .B0(n2300), .B1(n2519), .A0N(\register[3][27] ), .A1N(n2520), .Y(n199) );
  OAI2BB2XL U775 ( .B0(n2297), .B1(n2519), .A0N(\register[3][28] ), .A1N(n2520), .Y(n200) );
  OAI2BB2XL U776 ( .B0(n2295), .B1(n2519), .A0N(\register[3][29] ), .A1N(n2520), .Y(n201) );
  OAI2BB2XL U777 ( .B0(n2293), .B1(n2519), .A0N(\register[3][30] ), .A1N(n2517), .Y(n202) );
  OAI2BB2XL U778 ( .B0(n2291), .B1(n2519), .A0N(\register[3][31] ), .A1N(n2517), .Y(n203) );
  OAI2BB2XL U779 ( .B0(n2307), .B1(n2490), .A0N(\register[9][23] ), .A1N(n2490), .Y(n387) );
  OAI2BB2XL U780 ( .B0(n2303), .B1(n2490), .A0N(\register[9][25] ), .A1N(n2491), .Y(n389) );
  OAI2BB2XL U781 ( .B0(n2301), .B1(n2490), .A0N(\register[9][26] ), .A1N(n2491), .Y(n390) );
  OAI2BB2XL U782 ( .B0(n2299), .B1(n2490), .A0N(\register[9][27] ), .A1N(n2491), .Y(n391) );
  OAI2BB2XL U783 ( .B0(n2296), .B1(n2490), .A0N(\register[9][28] ), .A1N(n2491), .Y(n392) );
  OAI2BB2XL U784 ( .B0(n2294), .B1(n2490), .A0N(\register[9][29] ), .A1N(n2491), .Y(n393) );
  OAI2BB2XL U785 ( .B0(n2292), .B1(n2490), .A0N(\register[9][30] ), .A1N(n2486), .Y(n394) );
  OAI2BB2XL U786 ( .B0(n2290), .B1(n2490), .A0N(\register[9][31] ), .A1N(n2486), .Y(n395) );
  OAI2BB2XL U787 ( .B0(n2307), .B1(n2444), .A0N(\register[17][23] ), .A1N(
        n2444), .Y(n643) );
  OAI2BB2XL U788 ( .B0(n2303), .B1(n2444), .A0N(\register[17][25] ), .A1N(
        n2445), .Y(n645) );
  OAI2BB2XL U789 ( .B0(n2301), .B1(n2444), .A0N(\register[17][26] ), .A1N(
        n2445), .Y(n646) );
  OAI2BB2XL U790 ( .B0(n2299), .B1(n2444), .A0N(\register[17][27] ), .A1N(
        n2445), .Y(n647) );
  OAI2BB2XL U791 ( .B0(n2296), .B1(n2444), .A0N(\register[17][28] ), .A1N(
        n2445), .Y(n648) );
  OAI2BB2XL U792 ( .B0(n2294), .B1(n2444), .A0N(\register[17][29] ), .A1N(
        n2445), .Y(n649) );
  OAI2BB2XL U793 ( .B0(n2292), .B1(n2444), .A0N(\register[17][30] ), .A1N(
        n2441), .Y(n650) );
  OAI2BB2XL U794 ( .B0(n2290), .B1(n2444), .A0N(\register[17][31] ), .A1N(
        n2441), .Y(n651) );
  OAI2BB2XL U795 ( .B0(n2307), .B1(n2400), .A0N(\register[25][23] ), .A1N(
        n2400), .Y(n899) );
  OAI2BB2XL U796 ( .B0(n2303), .B1(n2400), .A0N(\register[25][25] ), .A1N(
        n2401), .Y(n901) );
  OAI2BB2XL U797 ( .B0(n2301), .B1(n2400), .A0N(\register[25][26] ), .A1N(
        n2401), .Y(n902) );
  OAI2BB2XL U798 ( .B0(n2298), .B1(n2400), .A0N(\register[25][27] ), .A1N(
        n2401), .Y(n903) );
  OAI2BB2XL U799 ( .B0(n2296), .B1(n2400), .A0N(\register[25][28] ), .A1N(
        n2401), .Y(n904) );
  OAI2BB2XL U800 ( .B0(n2294), .B1(n2400), .A0N(\register[25][29] ), .A1N(
        n2401), .Y(n905) );
  OAI2BB2XL U801 ( .B0(n2292), .B1(n2400), .A0N(\register[25][30] ), .A1N(
        n2397), .Y(n906) );
  OAI2BB2XL U802 ( .B0(n2290), .B1(n2400), .A0N(\register[25][31] ), .A1N(
        n2397), .Y(n907) );
  OAI2BB2XL U803 ( .B0(n2307), .B1(n2478), .A0N(\register[11][23] ), .A1N(
        n2478), .Y(n451) );
  OAI2BB2XL U804 ( .B0(n2303), .B1(n2478), .A0N(\register[11][25] ), .A1N(
        n2479), .Y(n453) );
  OAI2BB2XL U805 ( .B0(n2301), .B1(n2478), .A0N(\register[11][26] ), .A1N(
        n2479), .Y(n454) );
  OAI2BB2XL U806 ( .B0(n2299), .B1(n2478), .A0N(\register[11][27] ), .A1N(
        n2479), .Y(n455) );
  OAI2BB2XL U807 ( .B0(n2296), .B1(n2478), .A0N(\register[11][28] ), .A1N(
        n2479), .Y(n456) );
  OAI2BB2XL U808 ( .B0(n2294), .B1(n2478), .A0N(\register[11][29] ), .A1N(
        n2479), .Y(n457) );
  OAI2BB2XL U809 ( .B0(n2292), .B1(n2478), .A0N(\register[11][30] ), .A1N(
        n2474), .Y(n458) );
  OAI2BB2XL U810 ( .B0(n2290), .B1(n2478), .A0N(\register[11][31] ), .A1N(
        n2474), .Y(n459) );
  OAI2BB2XL U811 ( .B0(n2307), .B1(n2432), .A0N(\register[19][23] ), .A1N(
        n2432), .Y(n707) );
  OAI2BB2XL U812 ( .B0(n2303), .B1(n2432), .A0N(\register[19][25] ), .A1N(
        n2433), .Y(n709) );
  OAI2BB2XL U813 ( .B0(n2301), .B1(n2432), .A0N(\register[19][26] ), .A1N(
        n2433), .Y(n710) );
  OAI2BB2XL U814 ( .B0(n2299), .B1(n2432), .A0N(\register[19][27] ), .A1N(
        n2433), .Y(n711) );
  OAI2BB2XL U815 ( .B0(n2296), .B1(n2432), .A0N(\register[19][28] ), .A1N(
        n2433), .Y(n712) );
  OAI2BB2XL U816 ( .B0(n2294), .B1(n2432), .A0N(\register[19][29] ), .A1N(
        n2433), .Y(n713) );
  OAI2BB2XL U817 ( .B0(n2292), .B1(n2432), .A0N(\register[19][30] ), .A1N(
        n2429), .Y(n714) );
  OAI2BB2XL U818 ( .B0(n2290), .B1(n2432), .A0N(\register[19][31] ), .A1N(
        n2429), .Y(n715) );
  OAI2BB2XL U819 ( .B0(n2307), .B1(n2388), .A0N(\register[27][23] ), .A1N(
        n2388), .Y(n963) );
  OAI2BB2XL U820 ( .B0(n2303), .B1(n2388), .A0N(\register[27][25] ), .A1N(
        n2389), .Y(n965) );
  OAI2BB2XL U821 ( .B0(n2301), .B1(n2388), .A0N(\register[27][26] ), .A1N(
        n2389), .Y(n966) );
  OAI2BB2XL U822 ( .B0(n2298), .B1(n2388), .A0N(\register[27][27] ), .A1N(
        n2389), .Y(n967) );
  OAI2BB2XL U823 ( .B0(n2296), .B1(n2388), .A0N(\register[27][28] ), .A1N(
        n2389), .Y(n968) );
  OAI2BB2XL U824 ( .B0(n2294), .B1(n2388), .A0N(\register[27][29] ), .A1N(
        n2389), .Y(n969) );
  OAI2BB2XL U825 ( .B0(n2292), .B1(n2388), .A0N(\register[27][30] ), .A1N(
        n2386), .Y(n970) );
  OAI2BB2XL U826 ( .B0(n2290), .B1(n2388), .A0N(\register[27][31] ), .A1N(
        n2386), .Y(n971) );
  OAI2BB2XL U827 ( .B0(n2362), .B1(n2489), .A0N(\register[9][0] ), .A1N(n2486), 
        .Y(n364) );
  OAI2BB2XL U828 ( .B0(n2361), .B1(n2488), .A0N(\register[9][1] ), .A1N(n2486), 
        .Y(n365) );
  OAI2BB2XL U829 ( .B0(n2359), .B1(n2488), .A0N(\register[9][2] ), .A1N(n2486), 
        .Y(n366) );
  OAI2BB2XL U830 ( .B0(n2356), .B1(n2488), .A0N(\register[9][3] ), .A1N(n2491), 
        .Y(n367) );
  OAI2BB2XL U831 ( .B0(n2354), .B1(n2488), .A0N(\register[9][4] ), .A1N(n2486), 
        .Y(n368) );
  OAI2BB2XL U832 ( .B0(n2351), .B1(n2488), .A0N(\register[9][5] ), .A1N(n2491), 
        .Y(n369) );
  OAI2BB2XL U833 ( .B0(n2349), .B1(n2488), .A0N(\register[9][6] ), .A1N(n2491), 
        .Y(n370) );
  OAI2BB2XL U834 ( .B0(n2346), .B1(n2488), .A0N(\register[9][7] ), .A1N(n2491), 
        .Y(n371) );
  OAI2BB2XL U835 ( .B0(n2344), .B1(n2488), .A0N(\register[9][8] ), .A1N(n2491), 
        .Y(n372) );
  OAI2BB2XL U836 ( .B0(n2342), .B1(n2488), .A0N(\register[9][9] ), .A1N(n2491), 
        .Y(n373) );
  OAI2BB2XL U837 ( .B0(n2339), .B1(n2488), .A0N(\register[9][10] ), .A1N(n2491), .Y(n374) );
  OAI2BB2XL U838 ( .B0(n2337), .B1(n2488), .A0N(\register[9][11] ), .A1N(n2491), .Y(n375) );
  OAI2BB2XL U839 ( .B0(n2335), .B1(n2488), .A0N(\register[9][12] ), .A1N(n2491), .Y(n376) );
  OAI2BB2XL U840 ( .B0(n2332), .B1(n2489), .A0N(\register[9][13] ), .A1N(n2491), .Y(n377) );
  OAI2BB2XL U841 ( .B0(n2330), .B1(n2489), .A0N(\register[9][14] ), .A1N(n2491), .Y(n378) );
  OAI2BB2XL U842 ( .B0(n2327), .B1(n2489), .A0N(\register[9][15] ), .A1N(n2490), .Y(n379) );
  OAI2BB2XL U843 ( .B0(n2324), .B1(n2489), .A0N(\register[9][16] ), .A1N(n2491), .Y(n380) );
  OAI2BB2XL U844 ( .B0(n2322), .B1(n2489), .A0N(\register[9][17] ), .A1N(n2490), .Y(n381) );
  OAI2BB2XL U845 ( .B0(n2319), .B1(n2489), .A0N(\register[9][18] ), .A1N(n2490), .Y(n382) );
  OAI2BB2XL U846 ( .B0(n2316), .B1(n2489), .A0N(\register[9][19] ), .A1N(n2490), .Y(n383) );
  OAI2BB2XL U847 ( .B0(n2314), .B1(n2489), .A0N(\register[9][20] ), .A1N(n2490), .Y(n384) );
  OAI2BB2XL U848 ( .B0(n2312), .B1(n2489), .A0N(\register[9][21] ), .A1N(n2490), .Y(n385) );
  OAI2BB2XL U849 ( .B0(n2310), .B1(n2489), .A0N(\register[9][22] ), .A1N(n2491), .Y(n386) );
  OAI2BB2XL U850 ( .B0(n2305), .B1(n2489), .A0N(\register[9][24] ), .A1N(n2491), .Y(n388) );
  OAI2BB2XL U851 ( .B0(n2362), .B1(n2443), .A0N(\register[17][0] ), .A1N(n2441), .Y(n620) );
  OAI2BB2XL U852 ( .B0(n2361), .B1(n2442), .A0N(\register[17][1] ), .A1N(n2441), .Y(n621) );
  OAI2BB2XL U853 ( .B0(n2359), .B1(n2442), .A0N(\register[17][2] ), .A1N(n2441), .Y(n622) );
  OAI2BB2XL U854 ( .B0(n2356), .B1(n2442), .A0N(\register[17][3] ), .A1N(n2445), .Y(n623) );
  OAI2BB2XL U855 ( .B0(n2354), .B1(n2442), .A0N(\register[17][4] ), .A1N(n2441), .Y(n624) );
  OAI2BB2XL U856 ( .B0(n2351), .B1(n2442), .A0N(\register[17][5] ), .A1N(n2445), .Y(n625) );
  OAI2BB2XL U857 ( .B0(n2349), .B1(n2442), .A0N(\register[17][6] ), .A1N(n2445), .Y(n626) );
  OAI2BB2XL U858 ( .B0(n2346), .B1(n2442), .A0N(\register[17][7] ), .A1N(n2445), .Y(n627) );
  OAI2BB2XL U859 ( .B0(n2344), .B1(n2442), .A0N(\register[17][8] ), .A1N(n2445), .Y(n628) );
  OAI2BB2XL U860 ( .B0(n2342), .B1(n2442), .A0N(\register[17][9] ), .A1N(n2445), .Y(n629) );
  OAI2BB2XL U861 ( .B0(n2339), .B1(n2442), .A0N(\register[17][10] ), .A1N(
        n2445), .Y(n630) );
  OAI2BB2XL U862 ( .B0(n2337), .B1(n2442), .A0N(\register[17][11] ), .A1N(
        n2445), .Y(n631) );
  OAI2BB2XL U863 ( .B0(n2335), .B1(n2442), .A0N(\register[17][12] ), .A1N(
        n2445), .Y(n632) );
  OAI2BB2XL U864 ( .B0(n2332), .B1(n2443), .A0N(\register[17][13] ), .A1N(
        n2445), .Y(n633) );
  OAI2BB2XL U865 ( .B0(n2330), .B1(n2443), .A0N(\register[17][14] ), .A1N(
        n2445), .Y(n634) );
  OAI2BB2XL U866 ( .B0(n2327), .B1(n2443), .A0N(\register[17][15] ), .A1N(
        n2444), .Y(n635) );
  OAI2BB2XL U867 ( .B0(n2324), .B1(n2443), .A0N(\register[17][16] ), .A1N(
        n2445), .Y(n636) );
  OAI2BB2XL U868 ( .B0(n2322), .B1(n2443), .A0N(\register[17][17] ), .A1N(
        n2444), .Y(n637) );
  OAI2BB2XL U869 ( .B0(n2319), .B1(n2443), .A0N(\register[17][18] ), .A1N(
        n2444), .Y(n638) );
  OAI2BB2XL U870 ( .B0(n2316), .B1(n2443), .A0N(\register[17][19] ), .A1N(
        n2444), .Y(n639) );
  OAI2BB2XL U871 ( .B0(n2314), .B1(n2443), .A0N(\register[17][20] ), .A1N(
        n2444), .Y(n640) );
  OAI2BB2XL U872 ( .B0(n2312), .B1(n2443), .A0N(\register[17][21] ), .A1N(
        n2444), .Y(n641) );
  OAI2BB2XL U873 ( .B0(n2310), .B1(n2443), .A0N(\register[17][22] ), .A1N(
        n2445), .Y(n642) );
  OAI2BB2XL U874 ( .B0(n2305), .B1(n2443), .A0N(\register[17][24] ), .A1N(
        n2445), .Y(n644) );
  OAI2BB2XL U875 ( .B0(n2362), .B1(n2399), .A0N(\register[25][0] ), .A1N(n2397), .Y(n876) );
  OAI2BB2XL U876 ( .B0(n2360), .B1(n2398), .A0N(\register[25][1] ), .A1N(n2397), .Y(n877) );
  OAI2BB2XL U877 ( .B0(n2358), .B1(n2398), .A0N(\register[25][2] ), .A1N(n2397), .Y(n878) );
  OAI2BB2XL U878 ( .B0(n2355), .B1(n2398), .A0N(\register[25][3] ), .A1N(n2401), .Y(n879) );
  OAI2BB2XL U879 ( .B0(n2353), .B1(n2398), .A0N(\register[25][4] ), .A1N(n2397), .Y(n880) );
  OAI2BB2XL U880 ( .B0(n2351), .B1(n2398), .A0N(\register[25][5] ), .A1N(n2401), .Y(n881) );
  OAI2BB2XL U881 ( .B0(n2348), .B1(n2398), .A0N(\register[25][6] ), .A1N(n2401), .Y(n882) );
  OAI2BB2XL U882 ( .B0(n2346), .B1(n2398), .A0N(\register[25][7] ), .A1N(n2401), .Y(n883) );
  OAI2BB2XL U883 ( .B0(n2344), .B1(n2398), .A0N(\register[25][8] ), .A1N(n2401), .Y(n884) );
  OAI2BB2XL U884 ( .B0(n2341), .B1(n2398), .A0N(\register[25][9] ), .A1N(n2401), .Y(n885) );
  OAI2BB2XL U885 ( .B0(n2339), .B1(n2398), .A0N(\register[25][10] ), .A1N(
        n2401), .Y(n886) );
  OAI2BB2XL U886 ( .B0(n2337), .B1(n2398), .A0N(\register[25][11] ), .A1N(
        n2401), .Y(n887) );
  OAI2BB2XL U887 ( .B0(n2334), .B1(n2398), .A0N(\register[25][12] ), .A1N(
        n2401), .Y(n888) );
  OAI2BB2XL U888 ( .B0(n2332), .B1(n2399), .A0N(\register[25][13] ), .A1N(
        n2401), .Y(n889) );
  OAI2BB2XL U889 ( .B0(n2329), .B1(n2399), .A0N(\register[25][14] ), .A1N(
        n2401), .Y(n890) );
  OAI2BB2XL U890 ( .B0(n2326), .B1(n2399), .A0N(\register[25][15] ), .A1N(
        n2400), .Y(n891) );
  OAI2BB2XL U891 ( .B0(n2324), .B1(n2399), .A0N(\register[25][16] ), .A1N(
        n2401), .Y(n892) );
  OAI2BB2XL U892 ( .B0(n2321), .B1(n2399), .A0N(\register[25][17] ), .A1N(
        n2400), .Y(n893) );
  OAI2BB2XL U893 ( .B0(n2318), .B1(n2399), .A0N(\register[25][18] ), .A1N(
        n2400), .Y(n894) );
  OAI2BB2XL U894 ( .B0(n2316), .B1(n2399), .A0N(\register[25][19] ), .A1N(
        n2400), .Y(n895) );
  OAI2BB2XL U895 ( .B0(n2314), .B1(n2399), .A0N(\register[25][20] ), .A1N(
        n2400), .Y(n896) );
  OAI2BB2XL U896 ( .B0(n2312), .B1(n2399), .A0N(\register[25][21] ), .A1N(
        n2400), .Y(n897) );
  OAI2BB2XL U897 ( .B0(n2309), .B1(n2399), .A0N(\register[25][22] ), .A1N(
        n2401), .Y(n898) );
  OAI2BB2XL U898 ( .B0(n2305), .B1(n2399), .A0N(\register[25][24] ), .A1N(
        n2401), .Y(n900) );
  OAI2BB2XL U899 ( .B0(n2362), .B1(n2477), .A0N(\register[11][0] ), .A1N(n2474), .Y(n428) );
  OAI2BB2XL U900 ( .B0(n2361), .B1(n2476), .A0N(\register[11][1] ), .A1N(n2474), .Y(n429) );
  OAI2BB2XL U901 ( .B0(n2359), .B1(n2476), .A0N(\register[11][2] ), .A1N(n2474), .Y(n430) );
  OAI2BB2XL U902 ( .B0(n2356), .B1(n2476), .A0N(\register[11][3] ), .A1N(n2479), .Y(n431) );
  OAI2BB2XL U903 ( .B0(n2354), .B1(n2476), .A0N(\register[11][4] ), .A1N(n2474), .Y(n432) );
  OAI2BB2XL U904 ( .B0(n2351), .B1(n2476), .A0N(\register[11][5] ), .A1N(n2479), .Y(n433) );
  OAI2BB2XL U905 ( .B0(n2349), .B1(n2476), .A0N(\register[11][6] ), .A1N(n2479), .Y(n434) );
  OAI2BB2XL U906 ( .B0(n2346), .B1(n2476), .A0N(\register[11][7] ), .A1N(n2479), .Y(n435) );
  OAI2BB2XL U907 ( .B0(n2344), .B1(n2476), .A0N(\register[11][8] ), .A1N(n2479), .Y(n436) );
  OAI2BB2XL U908 ( .B0(n2342), .B1(n2476), .A0N(\register[11][9] ), .A1N(n2479), .Y(n437) );
  OAI2BB2XL U909 ( .B0(n2339), .B1(n2476), .A0N(\register[11][10] ), .A1N(
        n2479), .Y(n438) );
  OAI2BB2XL U910 ( .B0(n2337), .B1(n2476), .A0N(\register[11][11] ), .A1N(
        n2479), .Y(n439) );
  OAI2BB2XL U911 ( .B0(n2335), .B1(n2476), .A0N(\register[11][12] ), .A1N(
        n2479), .Y(n440) );
  OAI2BB2XL U912 ( .B0(n2332), .B1(n2477), .A0N(\register[11][13] ), .A1N(
        n2479), .Y(n441) );
  OAI2BB2XL U913 ( .B0(n2330), .B1(n2477), .A0N(\register[11][14] ), .A1N(
        n2479), .Y(n442) );
  OAI2BB2XL U914 ( .B0(n2327), .B1(n2477), .A0N(\register[11][15] ), .A1N(
        n2478), .Y(n443) );
  OAI2BB2XL U915 ( .B0(n2324), .B1(n2477), .A0N(\register[11][16] ), .A1N(
        n2479), .Y(n444) );
  OAI2BB2XL U916 ( .B0(n2322), .B1(n2477), .A0N(\register[11][17] ), .A1N(
        n2478), .Y(n445) );
  OAI2BB2XL U917 ( .B0(n2319), .B1(n2477), .A0N(\register[11][18] ), .A1N(
        n2478), .Y(n446) );
  OAI2BB2XL U918 ( .B0(n2316), .B1(n2477), .A0N(\register[11][19] ), .A1N(
        n2478), .Y(n447) );
  OAI2BB2XL U919 ( .B0(n2314), .B1(n2477), .A0N(\register[11][20] ), .A1N(
        n2478), .Y(n448) );
  OAI2BB2XL U920 ( .B0(n2312), .B1(n2477), .A0N(\register[11][21] ), .A1N(
        n2478), .Y(n449) );
  OAI2BB2XL U921 ( .B0(n2310), .B1(n2477), .A0N(\register[11][22] ), .A1N(
        n2479), .Y(n450) );
  OAI2BB2XL U922 ( .B0(n2305), .B1(n2477), .A0N(\register[11][24] ), .A1N(
        n2479), .Y(n452) );
  OAI2BB2XL U923 ( .B0(n2362), .B1(n2431), .A0N(\register[19][0] ), .A1N(n2429), .Y(n684) );
  OAI2BB2XL U924 ( .B0(n2361), .B1(n2430), .A0N(\register[19][1] ), .A1N(n2429), .Y(n685) );
  OAI2BB2XL U925 ( .B0(n2359), .B1(n2430), .A0N(\register[19][2] ), .A1N(n2429), .Y(n686) );
  OAI2BB2XL U926 ( .B0(n2356), .B1(n2430), .A0N(\register[19][3] ), .A1N(n2433), .Y(n687) );
  OAI2BB2XL U927 ( .B0(n2354), .B1(n2430), .A0N(\register[19][4] ), .A1N(n2429), .Y(n688) );
  OAI2BB2XL U928 ( .B0(n2351), .B1(n2430), .A0N(\register[19][5] ), .A1N(n2433), .Y(n689) );
  OAI2BB2XL U929 ( .B0(n2349), .B1(n2430), .A0N(\register[19][6] ), .A1N(n2433), .Y(n690) );
  OAI2BB2XL U930 ( .B0(n2346), .B1(n2430), .A0N(\register[19][7] ), .A1N(n2433), .Y(n691) );
  OAI2BB2XL U931 ( .B0(n2344), .B1(n2430), .A0N(\register[19][8] ), .A1N(n2433), .Y(n692) );
  OAI2BB2XL U932 ( .B0(n2342), .B1(n2430), .A0N(\register[19][9] ), .A1N(n2433), .Y(n693) );
  OAI2BB2XL U933 ( .B0(n2339), .B1(n2430), .A0N(\register[19][10] ), .A1N(
        n2433), .Y(n694) );
  OAI2BB2XL U934 ( .B0(n2337), .B1(n2430), .A0N(\register[19][11] ), .A1N(
        n2433), .Y(n695) );
  OAI2BB2XL U935 ( .B0(n2335), .B1(n2430), .A0N(\register[19][12] ), .A1N(
        n2433), .Y(n696) );
  OAI2BB2XL U936 ( .B0(n2332), .B1(n2431), .A0N(\register[19][13] ), .A1N(
        n2433), .Y(n697) );
  OAI2BB2XL U937 ( .B0(n2330), .B1(n2431), .A0N(\register[19][14] ), .A1N(
        n2433), .Y(n698) );
  OAI2BB2XL U938 ( .B0(n2327), .B1(n2431), .A0N(\register[19][15] ), .A1N(
        n2432), .Y(n699) );
  OAI2BB2XL U939 ( .B0(n2324), .B1(n2431), .A0N(\register[19][16] ), .A1N(
        n2433), .Y(n700) );
  OAI2BB2XL U940 ( .B0(n2322), .B1(n2431), .A0N(\register[19][17] ), .A1N(
        n2432), .Y(n701) );
  OAI2BB2XL U941 ( .B0(n2319), .B1(n2431), .A0N(\register[19][18] ), .A1N(
        n2432), .Y(n702) );
  OAI2BB2XL U942 ( .B0(n2316), .B1(n2431), .A0N(\register[19][19] ), .A1N(
        n2432), .Y(n703) );
  OAI2BB2XL U943 ( .B0(n2314), .B1(n2431), .A0N(\register[19][20] ), .A1N(
        n2432), .Y(n704) );
  OAI2BB2XL U944 ( .B0(n2312), .B1(n2431), .A0N(\register[19][21] ), .A1N(
        n2432), .Y(n705) );
  OAI2BB2XL U945 ( .B0(n2310), .B1(n2431), .A0N(\register[19][22] ), .A1N(
        n2433), .Y(n706) );
  OAI2BB2XL U946 ( .B0(n2305), .B1(n2431), .A0N(\register[19][24] ), .A1N(
        n2433), .Y(n708) );
  OAI2BB2XL U947 ( .B0(n2362), .B1(n2387), .A0N(\register[27][0] ), .A1N(n2386), .Y(n940) );
  OAI2BB2XL U948 ( .B0(n2360), .B1(n2386), .A0N(\register[27][1] ), .A1N(n2386), .Y(n941) );
  OAI2BB2XL U949 ( .B0(n2358), .B1(n2386), .A0N(\register[27][2] ), .A1N(n2386), .Y(n942) );
  OAI2BB2XL U950 ( .B0(n2355), .B1(n2386), .A0N(\register[27][3] ), .A1N(n2389), .Y(n943) );
  OAI2BB2XL U951 ( .B0(n2353), .B1(n2387), .A0N(\register[27][4] ), .A1N(n2386), .Y(n944) );
  OAI2BB2XL U952 ( .B0(n2351), .B1(n2386), .A0N(\register[27][5] ), .A1N(n2389), .Y(n945) );
  OAI2BB2XL U953 ( .B0(n2348), .B1(n2387), .A0N(\register[27][6] ), .A1N(n2389), .Y(n946) );
  OAI2BB2XL U954 ( .B0(n2346), .B1(n2386), .A0N(\register[27][7] ), .A1N(n2389), .Y(n947) );
  OAI2BB2XL U955 ( .B0(n2344), .B1(n2386), .A0N(\register[27][8] ), .A1N(n2389), .Y(n948) );
  OAI2BB2XL U956 ( .B0(n2341), .B1(n2387), .A0N(\register[27][9] ), .A1N(n2389), .Y(n949) );
  OAI2BB2XL U957 ( .B0(n2339), .B1(n2386), .A0N(\register[27][10] ), .A1N(
        n2389), .Y(n950) );
  OAI2BB2XL U958 ( .B0(n2337), .B1(n2386), .A0N(\register[27][11] ), .A1N(
        n2389), .Y(n951) );
  OAI2BB2XL U959 ( .B0(n2334), .B1(n2387), .A0N(\register[27][12] ), .A1N(
        n2389), .Y(n952) );
  OAI2BB2XL U960 ( .B0(n2332), .B1(n2387), .A0N(\register[27][13] ), .A1N(
        n2389), .Y(n953) );
  OAI2BB2XL U961 ( .B0(n2329), .B1(n2387), .A0N(\register[27][14] ), .A1N(
        n2389), .Y(n954) );
  OAI2BB2XL U962 ( .B0(n2326), .B1(n2387), .A0N(\register[27][15] ), .A1N(
        n2388), .Y(n955) );
  OAI2BB2XL U963 ( .B0(n2324), .B1(n2387), .A0N(\register[27][16] ), .A1N(
        n2389), .Y(n956) );
  OAI2BB2XL U964 ( .B0(n2321), .B1(n2387), .A0N(\register[27][17] ), .A1N(
        n2388), .Y(n957) );
  OAI2BB2XL U965 ( .B0(n2318), .B1(n2387), .A0N(\register[27][18] ), .A1N(
        n2388), .Y(n958) );
  OAI2BB2XL U966 ( .B0(n2316), .B1(n2387), .A0N(\register[27][19] ), .A1N(
        n2388), .Y(n959) );
  OAI2BB2XL U967 ( .B0(n2314), .B1(n2387), .A0N(\register[27][20] ), .A1N(
        n2388), .Y(n960) );
  OAI2BB2XL U968 ( .B0(n2312), .B1(n2387), .A0N(\register[27][21] ), .A1N(
        n2388), .Y(n961) );
  OAI2BB2XL U969 ( .B0(n2309), .B1(n2387), .A0N(\register[27][22] ), .A1N(
        n2389), .Y(n962) );
  OAI2BB2XL U970 ( .B0(n2305), .B1(n2387), .A0N(\register[27][24] ), .A1N(
        n2389), .Y(n964) );
  OAI2BB2XL U971 ( .B0(n2363), .B1(n2530), .A0N(\register[1][0] ), .A1N(n2528), 
        .Y(n108) );
  OAI2BB2XL U972 ( .B0(n2613), .B1(n2529), .A0N(\register[1][1] ), .A1N(n2528), 
        .Y(n109) );
  OAI2BB2XL U973 ( .B0(n2612), .B1(n2529), .A0N(\register[1][2] ), .A1N(n2528), 
        .Y(n110) );
  OAI2BB2XL U974 ( .B0(n2357), .B1(n2529), .A0N(\register[1][3] ), .A1N(n2532), 
        .Y(n111) );
  OAI2BB2XL U975 ( .B0(n2610), .B1(n2529), .A0N(\register[1][4] ), .A1N(n2528), 
        .Y(n112) );
  OAI2BB2XL U976 ( .B0(n2352), .B1(n2529), .A0N(\register[1][5] ), .A1N(n2532), 
        .Y(n113) );
  OAI2BB2XL U977 ( .B0(n2350), .B1(n2529), .A0N(\register[1][6] ), .A1N(n2532), 
        .Y(n114) );
  OAI2BB2XL U978 ( .B0(n2347), .B1(n2529), .A0N(\register[1][7] ), .A1N(n2532), 
        .Y(n115) );
  OAI2BB2XL U979 ( .B0(n2345), .B1(n2529), .A0N(\register[1][8] ), .A1N(n2532), 
        .Y(n116) );
  OAI2BB2XL U980 ( .B0(n2343), .B1(n2529), .A0N(\register[1][9] ), .A1N(n2532), 
        .Y(n117) );
  OAI2BB2XL U981 ( .B0(n2340), .B1(n2529), .A0N(\register[1][10] ), .A1N(n2532), .Y(n118) );
  OAI2BB2XL U982 ( .B0(n2338), .B1(n2529), .A0N(\register[1][11] ), .A1N(n2532), .Y(n119) );
  OAI2BB2XL U983 ( .B0(n2336), .B1(n2529), .A0N(\register[1][12] ), .A1N(n2532), .Y(n120) );
  OAI2BB2XL U984 ( .B0(n2333), .B1(n2530), .A0N(\register[1][13] ), .A1N(n2532), .Y(n121) );
  OAI2BB2XL U985 ( .B0(n2331), .B1(n2530), .A0N(\register[1][14] ), .A1N(n2532), .Y(n122) );
  OAI2BB2XL U986 ( .B0(n2328), .B1(n2530), .A0N(\register[1][15] ), .A1N(n2531), .Y(n123) );
  OAI2BB2XL U987 ( .B0(n2325), .B1(n2530), .A0N(\register[1][16] ), .A1N(n2532), .Y(n124) );
  OAI2BB2XL U988 ( .B0(n2323), .B1(n2530), .A0N(\register[1][17] ), .A1N(n2531), .Y(n125) );
  OAI2BB2XL U989 ( .B0(n2320), .B1(n2530), .A0N(\register[1][18] ), .A1N(n2531), .Y(n126) );
  OAI2BB2XL U990 ( .B0(n2317), .B1(n2530), .A0N(\register[1][19] ), .A1N(n2531), .Y(n127) );
  OAI2BB2XL U991 ( .B0(n2315), .B1(n2530), .A0N(\register[1][20] ), .A1N(n2531), .Y(n128) );
  OAI2BB2XL U992 ( .B0(n2313), .B1(n2530), .A0N(\register[1][21] ), .A1N(n2531), .Y(n129) );
  OAI2BB2XL U993 ( .B0(n2311), .B1(n2530), .A0N(\register[1][22] ), .A1N(n2532), .Y(n130) );
  OAI2BB2XL U994 ( .B0(n2306), .B1(n2530), .A0N(\register[1][24] ), .A1N(n2532), .Y(n132) );
  OAI2BB2XL U995 ( .B0(n2363), .B1(n2518), .A0N(\register[3][0] ), .A1N(n2517), 
        .Y(n172) );
  OAI2BB2XL U996 ( .B0(n2613), .B1(n2517), .A0N(\register[3][1] ), .A1N(n2517), 
        .Y(n173) );
  OAI2BB2XL U997 ( .B0(n2612), .B1(n2517), .A0N(\register[3][2] ), .A1N(n2517), 
        .Y(n174) );
  OAI2BB2XL U998 ( .B0(n2357), .B1(n2517), .A0N(\register[3][3] ), .A1N(n2520), 
        .Y(n175) );
  OAI2BB2XL U999 ( .B0(n2610), .B1(n2517), .A0N(\register[3][4] ), .A1N(n2517), 
        .Y(n176) );
  OAI2BB2XL U1000 ( .B0(n2352), .B1(n2517), .A0N(\register[3][5] ), .A1N(n2520), .Y(n177) );
  OAI2BB2XL U1001 ( .B0(n2350), .B1(n2517), .A0N(\register[3][6] ), .A1N(n2520), .Y(n178) );
  OAI2BB2XL U1002 ( .B0(n2347), .B1(n2517), .A0N(\register[3][7] ), .A1N(n2520), .Y(n179) );
  OAI2BB2XL U1003 ( .B0(n2345), .B1(n2517), .A0N(\register[3][8] ), .A1N(n2520), .Y(n180) );
  OAI2BB2XL U1004 ( .B0(n2343), .B1(n2518), .A0N(\register[3][9] ), .A1N(n2520), .Y(n181) );
  OAI2BB2XL U1005 ( .B0(n2340), .B1(n2518), .A0N(\register[3][10] ), .A1N(
        n2520), .Y(n182) );
  OAI2BB2XL U1006 ( .B0(n2338), .B1(n2518), .A0N(\register[3][11] ), .A1N(
        n2520), .Y(n183) );
  OAI2BB2XL U1007 ( .B0(n2336), .B1(n2518), .A0N(\register[3][12] ), .A1N(
        n2520), .Y(n184) );
  OAI2BB2XL U1008 ( .B0(n2333), .B1(n2518), .A0N(\register[3][13] ), .A1N(
        n2520), .Y(n185) );
  OAI2BB2XL U1009 ( .B0(n2331), .B1(n2518), .A0N(\register[3][14] ), .A1N(
        n2520), .Y(n186) );
  OAI2BB2XL U1010 ( .B0(n2328), .B1(n2518), .A0N(\register[3][15] ), .A1N(
        n2519), .Y(n187) );
  OAI2BB2XL U1011 ( .B0(n2325), .B1(n2518), .A0N(\register[3][16] ), .A1N(
        n2520), .Y(n188) );
  OAI2BB2XL U1012 ( .B0(n2323), .B1(n2518), .A0N(\register[3][17] ), .A1N(
        n2519), .Y(n189) );
  OAI2BB2XL U1013 ( .B0(n2320), .B1(n2518), .A0N(\register[3][18] ), .A1N(
        n2519), .Y(n190) );
  OAI2BB2XL U1014 ( .B0(n2317), .B1(n2518), .A0N(\register[3][19] ), .A1N(
        n2519), .Y(n191) );
  OAI2BB2XL U1015 ( .B0(n2315), .B1(n2518), .A0N(\register[3][20] ), .A1N(
        n2519), .Y(n192) );
  OAI2BB2XL U1016 ( .B0(n2313), .B1(n2518), .A0N(\register[3][21] ), .A1N(
        n2519), .Y(n193) );
  OAI2BB2XL U1017 ( .B0(n2311), .B1(n2518), .A0N(\register[3][22] ), .A1N(
        n2520), .Y(n194) );
  OAI2BB2XL U1018 ( .B0(n2306), .B1(n2518), .A0N(\register[3][24] ), .A1N(
        n2520), .Y(n196) );
  OAI2BB2XL U1019 ( .B0(n2542), .B1(n2363), .A0N(N91), .A1N(n2543), .Y(
        rdata2[0]) );
  OAI2BB2XL U1020 ( .B0(n2541), .B1(n2613), .A0N(N90), .A1N(n2542), .Y(
        rdata2[1]) );
  OAI2BB2XL U1021 ( .B0(n2540), .B1(n2612), .A0N(N89), .A1N(n2543), .Y(
        rdata2[2]) );
  OAI2BB2XL U1022 ( .B0(n2540), .B1(n2357), .A0N(N88), .A1N(n2543), .Y(
        rdata2[3]) );
  OAI2BB2XL U1023 ( .B0(n2540), .B1(n2610), .A0N(N87), .A1N(n2543), .Y(
        rdata2[4]) );
  OAI2BB2XL U1024 ( .B0(n2540), .B1(n2352), .A0N(N86), .A1N(n2543), .Y(
        rdata2[5]) );
  OAI2BB2XL U1025 ( .B0(n2540), .B1(n2350), .A0N(N85), .A1N(n2543), .Y(
        rdata2[6]) );
  OAI2BB2XL U1026 ( .B0(n2540), .B1(n2347), .A0N(N84), .A1N(n2543), .Y(
        rdata2[7]) );
  OAI2BB2XL U1027 ( .B0(n2540), .B1(n2345), .A0N(N83), .A1N(n2543), .Y(
        rdata2[8]) );
  OAI2BB2XL U1028 ( .B0(n2541), .B1(n2343), .A0N(N82), .A1N(n2543), .Y(
        rdata2[9]) );
  OAI2BB2XL U1029 ( .B0(n2542), .B1(n2340), .A0N(N81), .A1N(n2543), .Y(
        rdata2[10]) );
  OAI2BB2XL U1030 ( .B0(n2542), .B1(n2338), .A0N(N80), .A1N(n2543), .Y(
        rdata2[11]) );
  OAI2BB2XL U1031 ( .B0(n2542), .B1(n2336), .A0N(N79), .A1N(n2543), .Y(
        rdata2[12]) );
  OAI2BB2XL U1032 ( .B0(n2542), .B1(n2333), .A0N(N78), .A1N(n2543), .Y(
        rdata2[13]) );
  OAI2BB2XL U1033 ( .B0(n2542), .B1(n2331), .A0N(N77), .A1N(n2543), .Y(
        rdata2[14]) );
  OAI2BB2XL U1034 ( .B0(n2542), .B1(n2328), .A0N(N76), .A1N(n2543), .Y(
        rdata2[15]) );
  OAI2BB2XL U1035 ( .B0(n2541), .B1(n2325), .A0N(N75), .A1N(n2543), .Y(
        rdata2[16]) );
  OAI2BB2XL U1036 ( .B0(n2542), .B1(n2323), .A0N(N74), .A1N(n2542), .Y(
        rdata2[17]) );
  OAI2BB2XL U1037 ( .B0(n2541), .B1(n2320), .A0N(N73), .A1N(n2543), .Y(
        rdata2[18]) );
  OAI2BB2XL U1038 ( .B0(n2541), .B1(n2317), .A0N(N72), .A1N(n2542), .Y(
        rdata2[19]) );
  OAI2BB2XL U1039 ( .B0(n2541), .B1(n2315), .A0N(N71), .A1N(n2542), .Y(
        rdata2[20]) );
  OAI2BB2XL U1040 ( .B0(n2541), .B1(n2313), .A0N(N70), .A1N(n2542), .Y(
        rdata2[21]) );
  OAI2BB2XL U1041 ( .B0(n2541), .B1(n2311), .A0N(N69), .A1N(n2542), .Y(
        rdata2[22]) );
  OAI2BB2XL U1042 ( .B0(n2541), .B1(n2308), .A0N(N68), .A1N(n2543), .Y(
        rdata2[23]) );
  OAI2BB2XL U1043 ( .B0(n2541), .B1(n2306), .A0N(N67), .A1N(n2542), .Y(
        rdata2[24]) );
  OAI2BB2XL U1044 ( .B0(n2541), .B1(n2304), .A0N(N66), .A1N(n2543), .Y(
        rdata2[25]) );
  OAI2BB2XL U1045 ( .B0(n2541), .B1(n2302), .A0N(N65), .A1N(n2543), .Y(
        rdata2[26]) );
  OAI2BB2XL U1046 ( .B0(n2540), .B1(n2300), .A0N(N64), .A1N(n2543), .Y(
        rdata2[27]) );
  OAI2BB2XL U1047 ( .B0(n2540), .B1(n2297), .A0N(N63), .A1N(n2543), .Y(
        rdata2[28]) );
  OAI2BB2XL U1048 ( .B0(n2540), .B1(n2295), .A0N(N62), .A1N(n2543), .Y(
        rdata2[29]) );
  OAI2BB2XL U1049 ( .B0(n2540), .B1(n2293), .A0N(N61), .A1N(n2543), .Y(
        rdata2[30]) );
  OAI2BB2XL U1050 ( .B0(n2540), .B1(n2291), .A0N(N60), .A1N(n2543), .Y(
        rdata2[31]) );
  OAI2BB2XL U1051 ( .B0(n2363), .B1(n2537), .A0N(N56), .A1N(n2538), .Y(
        rdata1[0]) );
  OAI2BB2XL U1052 ( .B0(n2613), .B1(n2536), .A0N(N55), .A1N(n2537), .Y(
        rdata1[1]) );
  OAI2BB2XL U1053 ( .B0(n2612), .B1(n2535), .A0N(N54), .A1N(n2538), .Y(
        rdata1[2]) );
  OAI2BB2XL U1054 ( .B0(n2357), .B1(n2535), .A0N(N53), .A1N(n2538), .Y(
        rdata1[3]) );
  OAI2BB2XL U1055 ( .B0(n2610), .B1(n2535), .A0N(N52), .A1N(n2538), .Y(
        rdata1[4]) );
  OAI2BB2XL U1056 ( .B0(n2352), .B1(n2535), .A0N(N51), .A1N(n2538), .Y(
        rdata1[5]) );
  OAI2BB2XL U1057 ( .B0(n2350), .B1(n2535), .A0N(N50), .A1N(n2538), .Y(
        rdata1[6]) );
  OAI2BB2XL U1058 ( .B0(n2347), .B1(n2535), .A0N(N49), .A1N(n2536), .Y(
        rdata1[7]) );
  OAI2BB2XL U1059 ( .B0(n2345), .B1(n2535), .A0N(N48), .A1N(n2538), .Y(
        rdata1[8]) );
  OAI2BB2XL U1060 ( .B0(n2343), .B1(n2536), .A0N(N47), .A1N(n2538), .Y(
        rdata1[9]) );
  OAI2BB2XL U1061 ( .B0(n2340), .B1(n2537), .A0N(N46), .A1N(n2538), .Y(
        rdata1[10]) );
  OAI2BB2XL U1062 ( .B0(n2338), .B1(n2537), .A0N(N45), .A1N(n2538), .Y(
        rdata1[11]) );
  OAI2BB2XL U1063 ( .B0(n2336), .B1(n2537), .A0N(N44), .A1N(n2538), .Y(
        rdata1[12]) );
  OAI2BB2XL U1064 ( .B0(n2333), .B1(n2537), .A0N(N43), .A1N(n2538), .Y(
        rdata1[13]) );
  OAI2BB2XL U1065 ( .B0(n2331), .B1(n2537), .A0N(N42), .A1N(n2538), .Y(
        rdata1[14]) );
  OAI2BB2XL U1066 ( .B0(n2328), .B1(n2537), .A0N(N41), .A1N(n2538), .Y(
        rdata1[15]) );
  OAI2BB2XL U1067 ( .B0(n2325), .B1(n2536), .A0N(N40), .A1N(n2538), .Y(
        rdata1[16]) );
  OAI2BB2XL U1068 ( .B0(n2323), .B1(n2537), .A0N(N39), .A1N(n2537), .Y(
        rdata1[17]) );
  OAI2BB2XL U1069 ( .B0(n2320), .B1(n2536), .A0N(N38), .A1N(n2538), .Y(
        rdata1[18]) );
  OAI2BB2XL U1070 ( .B0(n2317), .B1(n2536), .A0N(N37), .A1N(n2537), .Y(
        rdata1[19]) );
  OAI2BB2XL U1071 ( .B0(n2315), .B1(n2536), .A0N(N36), .A1N(n2537), .Y(
        rdata1[20]) );
  OAI2BB2XL U1072 ( .B0(n2313), .B1(n2536), .A0N(N35), .A1N(n2537), .Y(
        rdata1[21]) );
  OAI2BB2XL U1073 ( .B0(n2311), .B1(n2536), .A0N(N34), .A1N(n2537), .Y(
        rdata1[22]) );
  OAI2BB2XL U1074 ( .B0(n2308), .B1(n2536), .A0N(N33), .A1N(n2538), .Y(
        rdata1[23]) );
  OAI2BB2XL U1075 ( .B0(n2306), .B1(n2536), .A0N(N32), .A1N(n2537), .Y(
        rdata1[24]) );
  OAI2BB2XL U1076 ( .B0(n2304), .B1(n2536), .A0N(N31), .A1N(n2538), .Y(
        rdata1[25]) );
  OAI2BB2XL U1077 ( .B0(n2302), .B1(n2536), .A0N(N30), .A1N(n2538), .Y(
        rdata1[26]) );
  OAI2BB2XL U1078 ( .B0(n2300), .B1(n2535), .A0N(N29), .A1N(n2538), .Y(
        rdata1[27]) );
  OAI2BB2XL U1079 ( .B0(n2297), .B1(n2535), .A0N(N28), .A1N(n2538), .Y(
        rdata1[28]) );
  OAI2BB2XL U1080 ( .B0(n2295), .B1(n2535), .A0N(N27), .A1N(n2538), .Y(
        rdata1[29]) );
  OAI2BB2XL U1081 ( .B0(n2293), .B1(n2535), .A0N(N26), .A1N(n2538), .Y(
        rdata1[30]) );
  OAI2BB2XL U1082 ( .B0(n2291), .B1(n2535), .A0N(N25), .A1N(n2538), .Y(
        rdata1[31]) );
  CLKINVX2 U1083 ( .A(wen), .Y(n2620) );
  MXI2X1 U1084 ( .A(n1626), .B(n1627), .S0(n2106), .Y(N91) );
  MX4X1 U1085 ( .A(n1693), .B(n1691), .C(n1692), .D(n1690), .S0(n2111), .S1(
        n2119), .Y(n1627) );
  MX4X1 U1086 ( .A(n1697), .B(n1695), .C(n1696), .D(n1694), .S0(n2111), .S1(
        n2119), .Y(n1626) );
  MXI4X1 U1087 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n2165), .S1(n2141), .Y(
        n1693) );
  MXI2X1 U1088 ( .A(n1628), .B(n1629), .S0(n2106), .Y(N90) );
  MX4X1 U1089 ( .A(n1705), .B(n1703), .C(n1704), .D(n1702), .S0(n2111), .S1(
        n2119), .Y(n1628) );
  MX4X1 U1090 ( .A(n1701), .B(n1699), .C(n1700), .D(n1698), .S0(n2111), .S1(
        n2119), .Y(n1629) );
  MXI4X1 U1091 ( .A(\register[8][1] ), .B(\register[9][1] ), .C(
        \register[10][1] ), .D(\register[11][1] ), .S0(n2166), .S1(n2141), .Y(
        n1703) );
  MXI2X1 U1092 ( .A(n1630), .B(n1631), .S0(n2106), .Y(N89) );
  MX4X1 U1093 ( .A(n1713), .B(n1711), .C(n1712), .D(n1710), .S0(n2112), .S1(
        n2120), .Y(n1630) );
  MX4X1 U1094 ( .A(n1709), .B(n1707), .C(n1708), .D(n1706), .S0(n2112), .S1(
        n2120), .Y(n1631) );
  MXI4X1 U1095 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n2166), .S1(n2141), .Y(
        n1711) );
  MXI2X1 U1096 ( .A(n1632), .B(n1633), .S0(n2106), .Y(N88) );
  MX4X1 U1097 ( .A(n1721), .B(n1719), .C(n1720), .D(n1718), .S0(n2112), .S1(
        n2120), .Y(n1632) );
  MX4X1 U1098 ( .A(n1717), .B(n1715), .C(n1716), .D(n1714), .S0(n2112), .S1(
        n2120), .Y(n1633) );
  MXI4X1 U1099 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n2167), .S1(n2142), .Y(
        n1719) );
  MXI2X1 U1100 ( .A(n1634), .B(n1635), .S0(n2106), .Y(N87) );
  MX4X1 U1101 ( .A(n1729), .B(n1727), .C(n1728), .D(n1726), .S0(n2112), .S1(
        n2120), .Y(n1634) );
  MX4X1 U1102 ( .A(n1725), .B(n1723), .C(n1724), .D(n1722), .S0(n2112), .S1(
        n2120), .Y(n1635) );
  MXI4X1 U1103 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n2167), .S1(n2142), .Y(
        n1727) );
  MXI2X1 U1104 ( .A(n1636), .B(n1637), .S0(n2106), .Y(N86) );
  MX4X1 U1105 ( .A(n1733), .B(n1731), .C(n1732), .D(n1730), .S0(n2112), .S1(
        n2120), .Y(n1637) );
  MX4X1 U1106 ( .A(n1737), .B(n1735), .C(n1736), .D(n1734), .S0(n2112), .S1(
        n2120), .Y(n1636) );
  MXI4X1 U1107 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n2167), .S1(n2142), .Y(
        n1733) );
  MXI2X1 U1108 ( .A(n1638), .B(n1639), .S0(n2106), .Y(N85) );
  MX4X1 U1109 ( .A(n1745), .B(n1743), .C(n1744), .D(n1742), .S0(n2112), .S1(
        n2120), .Y(n1638) );
  MX4X1 U1110 ( .A(n1741), .B(n1739), .C(n1740), .D(n1738), .S0(n2112), .S1(
        n2120), .Y(n1639) );
  MXI4X1 U1111 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n2168), .S1(n2143), .Y(
        n1743) );
  MXI2X1 U1112 ( .A(n1640), .B(n1641), .S0(n2106), .Y(N84) );
  MX4X1 U1113 ( .A(n1749), .B(n1747), .C(n1748), .D(n1746), .S0(n2112), .S1(
        n2120), .Y(n1641) );
  MX4X1 U1114 ( .A(n1753), .B(n1751), .C(n1752), .D(n1750), .S0(n2112), .S1(
        n2120), .Y(n1640) );
  MXI2X1 U1115 ( .A(n1642), .B(n1643), .S0(n2107), .Y(N83) );
  MX4X1 U1116 ( .A(n1757), .B(n1755), .C(n1756), .D(n1754), .S0(n2113), .S1(
        n2121), .Y(n1643) );
  MX4X1 U1117 ( .A(n1761), .B(n1759), .C(n1760), .D(n1758), .S0(n2113), .S1(
        n2121), .Y(n1642) );
  MXI4X1 U1118 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n2169), .S1(n2143), .Y(
        n1757) );
  MXI2X1 U1119 ( .A(n1644), .B(n1645), .S0(n2107), .Y(N82) );
  MX4X1 U1120 ( .A(n1765), .B(n1763), .C(n1764), .D(n1762), .S0(n2113), .S1(
        n2121), .Y(n1645) );
  MX4X1 U1121 ( .A(n1769), .B(n1767), .C(n1768), .D(n1766), .S0(n2113), .S1(
        n2121), .Y(n1644) );
  MXI4X1 U1122 ( .A(\register[16][9] ), .B(\register[17][9] ), .C(
        \register[18][9] ), .D(\register[19][9] ), .S0(n2169), .S1(n2144), .Y(
        n1765) );
  MXI2X1 U1123 ( .A(n1646), .B(n1647), .S0(n2107), .Y(N81) );
  MX4X1 U1124 ( .A(n1773), .B(n1771), .C(n1772), .D(n1770), .S0(n2113), .S1(
        n2121), .Y(n1647) );
  MX4X1 U1125 ( .A(n1777), .B(n1775), .C(n1776), .D(n1774), .S0(n2113), .S1(
        n2121), .Y(n1646) );
  MXI4X1 U1126 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1773) );
  MXI2X1 U1127 ( .A(n1648), .B(n1649), .S0(n2107), .Y(N80) );
  MX4X1 U1128 ( .A(n1781), .B(n1779), .C(n1780), .D(n1778), .S0(n2113), .S1(
        n2121), .Y(n1649) );
  MX4X1 U1129 ( .A(n1785), .B(n1783), .C(n1784), .D(n1782), .S0(n2113), .S1(
        n2121), .Y(n1648) );
  MXI4X1 U1130 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1781) );
  MXI2X1 U1131 ( .A(n1650), .B(n1651), .S0(n2107), .Y(N79) );
  MX4X1 U1132 ( .A(n1793), .B(n1791), .C(n1792), .D(n1790), .S0(n2113), .S1(
        n2121), .Y(n1650) );
  MX4X1 U1133 ( .A(n1789), .B(n1787), .C(n1788), .D(n1786), .S0(n2113), .S1(
        n2121), .Y(n1651) );
  MXI4X1 U1134 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n2171), .S1(n2145), 
        .Y(n1791) );
  MXI2X1 U1135 ( .A(n1652), .B(n1653), .S0(n2107), .Y(N78) );
  MX4X1 U1136 ( .A(n1797), .B(n1795), .C(n1796), .D(n1794), .S0(n2113), .S1(
        n2121), .Y(n1653) );
  MX4X1 U1137 ( .A(n1801), .B(n1799), .C(n1800), .D(n1798), .S0(n2113), .S1(
        n2121), .Y(n1652) );
  MXI4X1 U1138 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1797) );
  MXI2X1 U1139 ( .A(n1654), .B(n1655), .S0(n2107), .Y(N77) );
  MX4X1 U1140 ( .A(n1809), .B(n1807), .C(n1808), .D(n1806), .S0(n2114), .S1(
        n2122), .Y(n1654) );
  MX4X1 U1141 ( .A(n1805), .B(n1803), .C(n1804), .D(n1802), .S0(n2114), .S1(
        n2122), .Y(n1655) );
  MXI4X1 U1142 ( .A(\register[8][14] ), .B(\register[9][14] ), .C(
        \register[10][14] ), .D(\register[11][14] ), .S0(n2172), .S1(n2145), 
        .Y(n1807) );
  MXI2X1 U1143 ( .A(n1656), .B(n1657), .S0(n2107), .Y(N76) );
  MX4X1 U1144 ( .A(n1817), .B(n1815), .C(n1816), .D(n1814), .S0(n2114), .S1(
        n2122), .Y(n1656) );
  MX4X1 U1145 ( .A(n1813), .B(n1811), .C(n1812), .D(n1810), .S0(n2114), .S1(
        n2122), .Y(n1657) );
  MXI2X1 U1146 ( .A(n1658), .B(n1659), .S0(n2107), .Y(N75) );
  MX4X1 U1147 ( .A(n1821), .B(n1819), .C(n1820), .D(n1818), .S0(n2114), .S1(
        n2122), .Y(n1659) );
  MX4X1 U1148 ( .A(n1825), .B(n1823), .C(n1824), .D(n1822), .S0(n2114), .S1(
        n2122), .Y(n1658) );
  MXI4X1 U1149 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1821) );
  MXI2X1 U1150 ( .A(n1660), .B(n1661), .S0(n2107), .Y(N74) );
  MX4X1 U1151 ( .A(n1829), .B(n1827), .C(n1828), .D(n1826), .S0(n2114), .S1(
        n2122), .Y(n1661) );
  MX4X1 U1152 ( .A(n1833), .B(n1831), .C(n1832), .D(n1830), .S0(n2114), .S1(
        n2122), .Y(n1660) );
  MXI4X1 U1153 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1829) );
  MXI2X1 U1154 ( .A(n1662), .B(n1663), .S0(n2107), .Y(N73) );
  MX4X1 U1155 ( .A(n1837), .B(n1835), .C(n1836), .D(n1834), .S0(n2114), .S1(
        n2122), .Y(n1663) );
  MX4X1 U1156 ( .A(n1841), .B(n1839), .C(n1840), .D(n1838), .S0(n2114), .S1(
        n2122), .Y(n1662) );
  MXI4X1 U1157 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n2159), .S1(n2136), 
        .Y(n1837) );
  MXI2X1 U1158 ( .A(n1664), .B(n1665), .S0(n2107), .Y(N72) );
  MX4X1 U1159 ( .A(n1845), .B(n1843), .C(n1844), .D(n1842), .S0(n2114), .S1(
        n2122), .Y(n1665) );
  MX4X1 U1160 ( .A(n1849), .B(n1847), .C(n1848), .D(n1846), .S0(n2114), .S1(
        n2122), .Y(n1664) );
  MXI4X1 U1161 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n2159), .S1(n2137), 
        .Y(n1845) );
  MXI2X1 U1162 ( .A(n1666), .B(n1667), .S0(n2108), .Y(N71) );
  MX4X1 U1163 ( .A(n1853), .B(n1851), .C(n1852), .D(n1850), .S0(n2115), .S1(
        n2123), .Y(n1667) );
  MX4X1 U1164 ( .A(n1857), .B(n1855), .C(n1856), .D(n1854), .S0(n2115), .S1(
        n2123), .Y(n1666) );
  MXI2X1 U1165 ( .A(n1668), .B(n1669), .S0(n2108), .Y(N70) );
  MX4X1 U1166 ( .A(n1861), .B(n1859), .C(n1860), .D(n1858), .S0(n2115), .S1(
        n2123), .Y(n1669) );
  MX4X1 U1167 ( .A(n1865), .B(n1863), .C(n1864), .D(n1862), .S0(n2115), .S1(
        n2123), .Y(n1668) );
  MXI4X1 U1168 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1861) );
  MXI2X1 U1169 ( .A(n1670), .B(n1671), .S0(n2108), .Y(N69) );
  MX4X1 U1170 ( .A(n1869), .B(n1867), .C(n1868), .D(n1866), .S0(n2115), .S1(
        n2123), .Y(n1671) );
  MX4X1 U1171 ( .A(n1873), .B(n1871), .C(n1872), .D(n1870), .S0(n2115), .S1(
        n2123), .Y(n1670) );
  MXI4X1 U1172 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n2161), .S1(n2138), 
        .Y(n1869) );
  MXI2X1 U1173 ( .A(n1672), .B(n1673), .S0(n2108), .Y(N68) );
  MX4X1 U1174 ( .A(n1877), .B(n1875), .C(n1876), .D(n1874), .S0(n2115), .S1(
        n2123), .Y(n1673) );
  MX4X1 U1175 ( .A(n1881), .B(n1879), .C(n1880), .D(n1878), .S0(n2115), .S1(
        n2123), .Y(n1672) );
  MXI4X1 U1176 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1877) );
  MXI2X1 U1177 ( .A(n1674), .B(n1675), .S0(n2108), .Y(N67) );
  MX4X1 U1178 ( .A(n1885), .B(n1883), .C(n1884), .D(n1882), .S0(n2115), .S1(
        n2123), .Y(n1675) );
  MX4X1 U1179 ( .A(n1889), .B(n1887), .C(n1888), .D(n1886), .S0(n2115), .S1(
        n2123), .Y(n1674) );
  MXI4X1 U1180 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n2162), .S1(n2138), 
        .Y(n1885) );
  MXI2X1 U1181 ( .A(n1676), .B(n1677), .S0(n2108), .Y(N66) );
  MX4X1 U1182 ( .A(n1893), .B(n1891), .C(n1892), .D(n1890), .S0(n2115), .S1(
        n2123), .Y(n1677) );
  MX4X1 U1183 ( .A(n1897), .B(n1895), .C(n1896), .D(n1894), .S0(n2115), .S1(
        n2123), .Y(n1676) );
  MXI4X1 U1184 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n2162), .S1(n2139), 
        .Y(n1893) );
  MXI2X1 U1185 ( .A(n1678), .B(n1679), .S0(n2108), .Y(N65) );
  MX4X1 U1186 ( .A(n1901), .B(n1899), .C(n1900), .D(n1898), .S0(n2112), .S1(
        n2124), .Y(n1679) );
  MX4X1 U1187 ( .A(n1905), .B(n1903), .C(n1904), .D(n1902), .S0(n2112), .S1(
        n2124), .Y(n1678) );
  MXI4X1 U1188 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n2162), .S1(n2139), 
        .Y(n1901) );
  MXI2X1 U1189 ( .A(n1680), .B(n1681), .S0(n2108), .Y(N64) );
  MX4X1 U1190 ( .A(n1909), .B(n1907), .C(n1908), .D(n1906), .S0(n2112), .S1(
        n2124), .Y(n1681) );
  MX4X1 U1191 ( .A(n1913), .B(n1911), .C(n1912), .D(n1910), .S0(n2112), .S1(
        n2124), .Y(n1680) );
  MXI4X1 U1192 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1909) );
  MXI2X1 U1193 ( .A(n1682), .B(n1683), .S0(n2108), .Y(N63) );
  MX4X1 U1194 ( .A(n1917), .B(n1915), .C(n1916), .D(n1914), .S0(n2112), .S1(
        n2124), .Y(n1683) );
  MX4X1 U1195 ( .A(n1921), .B(n1919), .C(n1920), .D(n1918), .S0(n2112), .S1(
        n2124), .Y(n1682) );
  MXI4X1 U1196 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n2163), .S1(n2140), 
        .Y(n1917) );
  MXI2X1 U1197 ( .A(n1684), .B(n1685), .S0(n2108), .Y(N62) );
  MX4X1 U1198 ( .A(n1925), .B(n1923), .C(n1924), .D(n1922), .S0(n2112), .S1(
        n2124), .Y(n1685) );
  MX4X1 U1199 ( .A(n1929), .B(n1927), .C(n1928), .D(n1926), .S0(n2112), .S1(
        n2124), .Y(n1684) );
  MXI4X1 U1200 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1925) );
  MXI2X1 U1201 ( .A(n1686), .B(n1687), .S0(n2108), .Y(N61) );
  MX4X1 U1202 ( .A(n1933), .B(n1931), .C(n1932), .D(n1930), .S0(n2112), .S1(
        n2124), .Y(n1687) );
  MX4X1 U1203 ( .A(n1937), .B(n1935), .C(n1936), .D(n1934), .S0(n2112), .S1(
        n2124), .Y(n1686) );
  MXI4X1 U1204 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1933) );
  MXI2X1 U1205 ( .A(n1688), .B(n1689), .S0(n2108), .Y(N60) );
  MX4X1 U1206 ( .A(n1941), .B(n1939), .C(n1940), .D(n1938), .S0(n2112), .S1(
        n2124), .Y(n1689) );
  MX4X1 U1207 ( .A(n1945), .B(n1943), .C(n1944), .D(n1942), .S0(n2112), .S1(
        n2124), .Y(n1688) );
  MXI4X1 U1208 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n2165), .S1(n2140), 
        .Y(n1941) );
  MXI2X1 U1209 ( .A(n32), .B(n33), .S0(n1556), .Y(N56) );
  MX4X1 U1210 ( .A(n1143), .B(n1141), .C(n1142), .D(n1140), .S0(n1561), .S1(
        n1568), .Y(n33) );
  MX4X1 U1211 ( .A(n1147), .B(n1145), .C(n1146), .D(n1144), .S0(n1561), .S1(
        n1568), .Y(n32) );
  MXI4X1 U1212 ( .A(\register[16][0] ), .B(\register[17][0] ), .C(
        \register[18][0] ), .D(\register[19][0] ), .S0(n1615), .S1(n1590), .Y(
        n1143) );
  MXI2X1 U1213 ( .A(n34), .B(n35), .S0(n1556), .Y(N55) );
  MX4X1 U1214 ( .A(n1155), .B(n1153), .C(n1154), .D(n1152), .S0(n1561), .S1(
        n1568), .Y(n34) );
  MX4X1 U1215 ( .A(n1151), .B(n1149), .C(n1150), .D(n1148), .S0(n1561), .S1(
        n1568), .Y(n35) );
  MXI2X1 U1216 ( .A(n36), .B(n37), .S0(n1556), .Y(N54) );
  MX4X1 U1217 ( .A(n1163), .B(n1161), .C(n1162), .D(n1160), .S0(n1562), .S1(
        n1569), .Y(n36) );
  MX4X1 U1218 ( .A(n1159), .B(n1157), .C(n1158), .D(n1156), .S0(n1562), .S1(
        n1569), .Y(n37) );
  MXI4X1 U1219 ( .A(\register[8][2] ), .B(\register[9][2] ), .C(
        \register[10][2] ), .D(\register[11][2] ), .S0(n1616), .S1(n1590), .Y(
        n1161) );
  MXI2X1 U1220 ( .A(n38), .B(n39), .S0(n1556), .Y(N53) );
  MX4X1 U1221 ( .A(n1171), .B(n1169), .C(n1170), .D(n1168), .S0(n1562), .S1(
        n1569), .Y(n38) );
  MX4X1 U1222 ( .A(n1167), .B(n1165), .C(n1166), .D(n1164), .S0(n1562), .S1(
        n1569), .Y(n39) );
  MXI4X1 U1223 ( .A(\register[8][3] ), .B(\register[9][3] ), .C(
        \register[10][3] ), .D(\register[11][3] ), .S0(n1617), .S1(n1591), .Y(
        n1169) );
  MXI2X1 U1224 ( .A(n40), .B(n41), .S0(n1556), .Y(N52) );
  MX4X1 U1225 ( .A(n1179), .B(n1177), .C(n1178), .D(n1176), .S0(n1562), .S1(
        n1569), .Y(n40) );
  MX4X1 U1226 ( .A(n1175), .B(n1173), .C(n1174), .D(n1172), .S0(n1562), .S1(
        n1569), .Y(n41) );
  MXI4X1 U1227 ( .A(\register[8][4] ), .B(\register[9][4] ), .C(
        \register[10][4] ), .D(\register[11][4] ), .S0(n1617), .S1(n1591), .Y(
        n1177) );
  MXI2X1 U1228 ( .A(n42), .B(n43), .S0(n1556), .Y(N51) );
  MX4X1 U1229 ( .A(n1183), .B(n1181), .C(n1182), .D(n1180), .S0(n1562), .S1(
        n1569), .Y(n43) );
  MX4X1 U1230 ( .A(n1187), .B(n1185), .C(n1186), .D(n1184), .S0(n1562), .S1(
        n1569), .Y(n42) );
  MXI4X1 U1231 ( .A(\register[16][5] ), .B(\register[17][5] ), .C(
        \register[18][5] ), .D(\register[19][5] ), .S0(n1617), .S1(n1591), .Y(
        n1183) );
  MXI2X1 U1232 ( .A(n44), .B(n45), .S0(n1556), .Y(N50) );
  MX4X1 U1233 ( .A(n1195), .B(n1193), .C(n1194), .D(n1192), .S0(n1562), .S1(
        n1569), .Y(n44) );
  MX4X1 U1234 ( .A(n1191), .B(n1189), .C(n1190), .D(n1188), .S0(n1562), .S1(
        n1569), .Y(n45) );
  MXI4X1 U1235 ( .A(\register[8][6] ), .B(\register[9][6] ), .C(
        \register[10][6] ), .D(\register[11][6] ), .S0(n1623), .S1(n1592), .Y(
        n1193) );
  MXI2X1 U1236 ( .A(n46), .B(n67), .S0(n1556), .Y(N49) );
  MX4X1 U1237 ( .A(n1199), .B(n1197), .C(n1198), .D(n1196), .S0(n1562), .S1(
        n1569), .Y(n67) );
  MX4X1 U1238 ( .A(n1203), .B(n1201), .C(n1202), .D(n1200), .S0(n1562), .S1(
        n1569), .Y(n46) );
  MXI4X1 U1239 ( .A(\register[16][7] ), .B(\register[17][7] ), .C(
        \register[18][7] ), .D(\register[19][7] ), .S0(n1625), .S1(n1592), .Y(
        n1199) );
  MXI2X1 U1240 ( .A(n74), .B(n78), .S0(n1557), .Y(N48) );
  MX4X1 U1241 ( .A(n1211), .B(n1209), .C(n1210), .D(n1208), .S0(n1563), .S1(
        n1570), .Y(n74) );
  MX4X1 U1242 ( .A(n1207), .B(n1205), .C(n1206), .D(n1204), .S0(n1563), .S1(
        n1570), .Y(n78) );
  MXI4X1 U1243 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n1605), .S1(n1592), .Y(
        n1209) );
  MXI2X1 U1244 ( .A(n87), .B(n89), .S0(n1557), .Y(N47) );
  MX4X1 U1245 ( .A(n1215), .B(n1213), .C(n1214), .D(n1212), .S0(n1563), .S1(
        n1570), .Y(n89) );
  MX4X1 U1246 ( .A(n1219), .B(n1217), .C(n1218), .D(n1216), .S0(n1563), .S1(
        n1570), .Y(n87) );
  MXI2X1 U1247 ( .A(n96), .B(n98), .S0(n1557), .Y(N46) );
  MX4X1 U1248 ( .A(n1223), .B(n1221), .C(n1222), .D(n1220), .S0(n1563), .S1(
        n1570), .Y(n98) );
  MX4X1 U1249 ( .A(n1227), .B(n1225), .C(n1226), .D(n1224), .S0(n1563), .S1(
        n1570), .Y(n96) );
  MXI4X1 U1250 ( .A(\register[16][10] ), .B(\register[17][10] ), .C(
        \register[18][10] ), .D(\register[19][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1223) );
  MXI2X1 U1251 ( .A(n105), .B(n107), .S0(n1557), .Y(N45) );
  MX4X1 U1252 ( .A(n1231), .B(n1229), .C(n1230), .D(n1228), .S0(n1563), .S1(
        n1570), .Y(n107) );
  MX4X1 U1253 ( .A(n1235), .B(n1233), .C(n1234), .D(n1232), .S0(n1563), .S1(
        n1570), .Y(n105) );
  MXI4X1 U1254 ( .A(\register[16][11] ), .B(\register[17][11] ), .C(
        \register[18][11] ), .D(\register[19][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1231) );
  MXI2X1 U1255 ( .A(n1100), .B(n1101), .S0(n1557), .Y(N44) );
  MX4X1 U1256 ( .A(n1243), .B(n1241), .C(n1242), .D(n1240), .S0(n1563), .S1(
        n1570), .Y(n1100) );
  MX4X1 U1257 ( .A(n1239), .B(n1237), .C(n1238), .D(n1236), .S0(n1563), .S1(
        n1570), .Y(n1101) );
  MXI4X1 U1258 ( .A(\register[8][12] ), .B(\register[9][12] ), .C(
        \register[10][12] ), .D(\register[11][12] ), .S0(n1619), .S1(n1594), 
        .Y(n1241) );
  MXI2X1 U1259 ( .A(n1102), .B(n1103), .S0(n1557), .Y(N43) );
  MX4X1 U1260 ( .A(n1247), .B(n1245), .C(n1246), .D(n1244), .S0(n1563), .S1(
        n1570), .Y(n1103) );
  MX4X1 U1261 ( .A(n1251), .B(n1249), .C(n1250), .D(n1248), .S0(n1563), .S1(
        n1570), .Y(n1102) );
  MXI4X1 U1262 ( .A(\register[16][13] ), .B(\register[17][13] ), .C(
        \register[18][13] ), .D(\register[19][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1247) );
  MXI2X1 U1263 ( .A(n1104), .B(n1105), .S0(n1557), .Y(N42) );
  MX4X1 U1264 ( .A(n1259), .B(n1257), .C(n1258), .D(n1256), .S0(n1564), .S1(
        n1571), .Y(n1104) );
  MX4X1 U1265 ( .A(n1255), .B(n1253), .C(n1254), .D(n1252), .S0(n1564), .S1(
        n1571), .Y(n1105) );
  MXI2X1 U1266 ( .A(n1106), .B(n1107), .S0(n1557), .Y(N41) );
  MX4X1 U1267 ( .A(n1267), .B(n1265), .C(n1266), .D(n1264), .S0(n1564), .S1(
        n1571), .Y(n1106) );
  MX4X1 U1268 ( .A(n1263), .B(n1261), .C(n1262), .D(n1260), .S0(n1564), .S1(
        n1571), .Y(n1107) );
  MXI4X1 U1269 ( .A(\register[8][15] ), .B(\register[9][15] ), .C(
        \register[10][15] ), .D(\register[11][15] ), .S0(n1620), .S1(n1595), 
        .Y(n1265) );
  MXI2X1 U1270 ( .A(n1108), .B(n1109), .S0(n1557), .Y(N40) );
  MX4X1 U1271 ( .A(n1271), .B(n1269), .C(n1270), .D(n1268), .S0(n1564), .S1(
        n1571), .Y(n1109) );
  MX4X1 U1272 ( .A(n1275), .B(n1273), .C(n1274), .D(n1272), .S0(n1564), .S1(
        n1571), .Y(n1108) );
  MXI4X1 U1273 ( .A(\register[16][16] ), .B(\register[17][16] ), .C(
        \register[18][16] ), .D(\register[19][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1271) );
  MXI2X1 U1274 ( .A(n1110), .B(n1111), .S0(n1557), .Y(N39) );
  MX4X1 U1275 ( .A(n1279), .B(n1277), .C(n1278), .D(n1276), .S0(n1564), .S1(
        n1571), .Y(n1111) );
  MX4X1 U1276 ( .A(n1283), .B(n1281), .C(n1282), .D(n1280), .S0(n1564), .S1(
        n1571), .Y(n1110) );
  MXI4X1 U1277 ( .A(\register[16][17] ), .B(\register[17][17] ), .C(
        \register[18][17] ), .D(\register[19][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1279) );
  MXI2X1 U1278 ( .A(n1112), .B(n1113), .S0(n1557), .Y(N38) );
  MX4X1 U1279 ( .A(n1287), .B(n1285), .C(n1286), .D(n1284), .S0(n1564), .S1(
        n1571), .Y(n1113) );
  MX4X1 U1280 ( .A(n1291), .B(n1289), .C(n1290), .D(n1288), .S0(n1564), .S1(
        n1571), .Y(n1112) );
  MXI4X1 U1281 ( .A(\register[16][18] ), .B(\register[17][18] ), .C(
        \register[18][18] ), .D(\register[19][18] ), .S0(n1609), .S1(n1585), 
        .Y(n1287) );
  MXI2X1 U1282 ( .A(n1114), .B(n1115), .S0(n1557), .Y(N37) );
  MX4X1 U1283 ( .A(n1295), .B(n1293), .C(n1294), .D(n1292), .S0(n1564), .S1(
        n1571), .Y(n1115) );
  MX4X1 U1284 ( .A(n1299), .B(n1297), .C(n1298), .D(n1296), .S0(n1564), .S1(
        n1571), .Y(n1114) );
  MXI4X1 U1285 ( .A(\register[16][19] ), .B(\register[17][19] ), .C(
        \register[18][19] ), .D(\register[19][19] ), .S0(n1609), .S1(n1586), 
        .Y(n1295) );
  MXI2X1 U1286 ( .A(n1116), .B(n1117), .S0(n1558), .Y(N36) );
  MX4X1 U1287 ( .A(n1303), .B(n1301), .C(n1302), .D(n1300), .S0(n1565), .S1(
        n1572), .Y(n1117) );
  MX4X1 U1288 ( .A(n1307), .B(n1305), .C(n1306), .D(n1304), .S0(n1565), .S1(
        n1572), .Y(n1116) );
  MXI4X1 U1289 ( .A(\register[16][20] ), .B(\register[17][20] ), .C(
        \register[18][20] ), .D(\register[19][20] ), .S0(n1610), .S1(n1586), 
        .Y(n1303) );
  MXI2X1 U1290 ( .A(n1118), .B(n1119), .S0(n1558), .Y(N35) );
  MX4X1 U1291 ( .A(n1311), .B(n1309), .C(n1310), .D(n1308), .S0(n1565), .S1(
        n1572), .Y(n1119) );
  MX4X1 U1292 ( .A(n1315), .B(n1313), .C(n1314), .D(n1312), .S0(n1565), .S1(
        n1572), .Y(n1118) );
  MXI4X1 U1293 ( .A(\register[16][21] ), .B(\register[17][21] ), .C(
        \register[18][21] ), .D(\register[19][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1311) );
  MXI2X1 U1294 ( .A(n1120), .B(n1121), .S0(n1558), .Y(N34) );
  MX4X1 U1295 ( .A(n1319), .B(n1317), .C(n1318), .D(n1316), .S0(n1565), .S1(
        n1572), .Y(n1121) );
  MX4X1 U1296 ( .A(n1323), .B(n1321), .C(n1322), .D(n1320), .S0(n1565), .S1(
        n1572), .Y(n1120) );
  MXI4X1 U1297 ( .A(\register[16][22] ), .B(\register[17][22] ), .C(
        \register[18][22] ), .D(\register[19][22] ), .S0(n1611), .S1(n1587), 
        .Y(n1319) );
  MXI2X1 U1298 ( .A(n1122), .B(n1123), .S0(n1558), .Y(N33) );
  MX4X1 U1299 ( .A(n1327), .B(n1325), .C(n1326), .D(n1324), .S0(n1565), .S1(
        n1572), .Y(n1123) );
  MX4X1 U1300 ( .A(n1331), .B(n1329), .C(n1330), .D(n1328), .S0(n1565), .S1(
        n1572), .Y(n1122) );
  MXI4X1 U1301 ( .A(\register[16][23] ), .B(\register[17][23] ), .C(
        \register[18][23] ), .D(\register[19][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1327) );
  MXI2X1 U1302 ( .A(n1124), .B(n1125), .S0(n1558), .Y(N32) );
  MX4X1 U1303 ( .A(n1335), .B(n1333), .C(n1334), .D(n1332), .S0(n1565), .S1(
        n1572), .Y(n1125) );
  MX4X1 U1304 ( .A(n1339), .B(n1337), .C(n1338), .D(n1336), .S0(n1565), .S1(
        n1572), .Y(n1124) );
  MXI4X1 U1305 ( .A(\register[16][24] ), .B(\register[17][24] ), .C(
        \register[18][24] ), .D(\register[19][24] ), .S0(n1612), .S1(n1587), 
        .Y(n1335) );
  MXI2X1 U1306 ( .A(n1126), .B(n1127), .S0(n1558), .Y(N31) );
  MX4X1 U1307 ( .A(n1343), .B(n1341), .C(n1342), .D(n1340), .S0(n1565), .S1(
        n1572), .Y(n1127) );
  MX4X1 U1308 ( .A(n1347), .B(n1345), .C(n1346), .D(n1344), .S0(n1565), .S1(
        n1572), .Y(n1126) );
  MXI4X1 U1309 ( .A(\register[16][25] ), .B(\register[17][25] ), .C(
        \register[18][25] ), .D(\register[19][25] ), .S0(n1612), .S1(n1588), 
        .Y(n1343) );
  MXI2X1 U1310 ( .A(n1128), .B(n1129), .S0(n1558), .Y(N30) );
  MX4X1 U1311 ( .A(n1351), .B(n1349), .C(n1350), .D(n1348), .S0(n1566), .S1(
        n1573), .Y(n1129) );
  MX4X1 U1312 ( .A(n1355), .B(n1353), .C(n1354), .D(n1352), .S0(n1566), .S1(
        n1573), .Y(n1128) );
  MXI4X1 U1313 ( .A(\register[16][26] ), .B(\register[17][26] ), .C(
        \register[18][26] ), .D(\register[19][26] ), .S0(n1612), .S1(n1588), 
        .Y(n1351) );
  MXI2X1 U1314 ( .A(n1130), .B(n1131), .S0(n1558), .Y(N29) );
  MX4X1 U1315 ( .A(n1359), .B(n1357), .C(n1358), .D(n1356), .S0(n1566), .S1(
        n1573), .Y(n1131) );
  MX4X1 U1316 ( .A(n1363), .B(n1361), .C(n1362), .D(n1360), .S0(n1566), .S1(
        n1573), .Y(n1130) );
  MXI4X1 U1317 ( .A(\register[16][27] ), .B(\register[17][27] ), .C(
        \register[18][27] ), .D(\register[19][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1359) );
  MXI2X1 U1318 ( .A(n1132), .B(n1133), .S0(n1558), .Y(N28) );
  MX4X1 U1319 ( .A(n1367), .B(n1365), .C(n1366), .D(n1364), .S0(n1566), .S1(
        n1573), .Y(n1133) );
  MX4X1 U1320 ( .A(n1371), .B(n1369), .C(n1370), .D(n1368), .S0(n1566), .S1(
        n1573), .Y(n1132) );
  MXI4X1 U1321 ( .A(\register[16][28] ), .B(\register[17][28] ), .C(
        \register[18][28] ), .D(\register[19][28] ), .S0(n1613), .S1(n1589), 
        .Y(n1367) );
  MXI2X1 U1322 ( .A(n1134), .B(n1135), .S0(n1558), .Y(N27) );
  MX4X1 U1323 ( .A(n1375), .B(n1373), .C(n1374), .D(n1372), .S0(n1566), .S1(
        n1573), .Y(n1135) );
  MX4X1 U1324 ( .A(n1379), .B(n1377), .C(n1378), .D(n1376), .S0(n1566), .S1(
        n1573), .Y(n1134) );
  MXI4X1 U1325 ( .A(\register[16][29] ), .B(\register[17][29] ), .C(
        \register[18][29] ), .D(\register[19][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1375) );
  MXI2X1 U1326 ( .A(n1136), .B(n1137), .S0(n1558), .Y(N26) );
  MX4X1 U1327 ( .A(n1383), .B(n1381), .C(n1382), .D(n1380), .S0(n1566), .S1(
        n1573), .Y(n1137) );
  MX4X1 U1328 ( .A(n1387), .B(n1385), .C(n1386), .D(n1384), .S0(n1566), .S1(
        n1573), .Y(n1136) );
  MXI4X1 U1329 ( .A(\register[16][30] ), .B(\register[17][30] ), .C(
        \register[18][30] ), .D(\register[19][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1383) );
  MXI2X1 U1330 ( .A(n1138), .B(n1139), .S0(n1558), .Y(N25) );
  MX4X1 U1331 ( .A(n1391), .B(n1389), .C(n1390), .D(n1388), .S0(n1566), .S1(
        n1573), .Y(n1139) );
  MX4X1 U1332 ( .A(n1395), .B(n1393), .C(n1394), .D(n1392), .S0(n1566), .S1(
        n1573), .Y(n1138) );
  MXI4X1 U1333 ( .A(\register[16][31] ), .B(\register[17][31] ), .C(
        \register[18][31] ), .D(\register[19][31] ), .S0(n1615), .S1(n1589), 
        .Y(n1391) );
  OAI2BB2XL U1334 ( .B0(n2308), .B1(n2515), .A0N(\register[4][23] ), .A1N(
        n2515), .Y(n227) );
  OAI2BB2XL U1335 ( .B0(n2304), .B1(n2515), .A0N(\register[4][25] ), .A1N(
        n2516), .Y(n229) );
  OAI2BB2XL U1336 ( .B0(n2302), .B1(n2515), .A0N(\register[4][26] ), .A1N(
        n2516), .Y(n230) );
  OAI2BB2XL U1337 ( .B0(n2300), .B1(n2515), .A0N(\register[4][27] ), .A1N(
        n2516), .Y(n231) );
  OAI2BB2XL U1338 ( .B0(n2297), .B1(n2515), .A0N(\register[4][28] ), .A1N(
        n2516), .Y(n232) );
  OAI2BB2XL U1339 ( .B0(n2295), .B1(n2515), .A0N(\register[4][29] ), .A1N(
        n2516), .Y(n233) );
  OAI2BB2XL U1340 ( .B0(n2293), .B1(n2515), .A0N(\register[4][30] ), .A1N(
        n2513), .Y(n234) );
  OAI2BB2XL U1341 ( .B0(n2291), .B1(n2515), .A0N(\register[4][31] ), .A1N(
        n2513), .Y(n235) );
  OAI2BB2XL U1342 ( .B0(n2308), .B1(n2506), .A0N(\register[6][23] ), .A1N(
        n2506), .Y(n291) );
  OAI2BB2XL U1343 ( .B0(n2304), .B1(n2506), .A0N(\register[6][25] ), .A1N(
        n2507), .Y(n293) );
  OAI2BB2XL U1344 ( .B0(n2302), .B1(n2506), .A0N(\register[6][26] ), .A1N(
        n2507), .Y(n294) );
  OAI2BB2XL U1345 ( .B0(n2300), .B1(n2506), .A0N(\register[6][27] ), .A1N(
        n2507), .Y(n295) );
  OAI2BB2XL U1346 ( .B0(n2297), .B1(n2506), .A0N(\register[6][28] ), .A1N(
        n2507), .Y(n296) );
  OAI2BB2XL U1347 ( .B0(n2295), .B1(n2506), .A0N(\register[6][29] ), .A1N(
        n2507), .Y(n297) );
  OAI2BB2XL U1348 ( .B0(n2293), .B1(n2506), .A0N(\register[6][30] ), .A1N(
        n2503), .Y(n298) );
  OAI2BB2XL U1349 ( .B0(n2291), .B1(n2506), .A0N(\register[6][31] ), .A1N(
        n2503), .Y(n299) );
  OAI2BB2XL U1350 ( .B0(n2307), .B1(n2471), .A0N(\register[12][23] ), .A1N(
        n2471), .Y(n483) );
  OAI2BB2XL U1351 ( .B0(n2303), .B1(n2471), .A0N(\register[12][25] ), .A1N(
        n2472), .Y(n485) );
  OAI2BB2XL U1352 ( .B0(n2301), .B1(n2471), .A0N(\register[12][26] ), .A1N(
        n2472), .Y(n486) );
  OAI2BB2XL U1353 ( .B0(n2299), .B1(n2471), .A0N(\register[12][27] ), .A1N(
        n2472), .Y(n487) );
  OAI2BB2XL U1354 ( .B0(n2296), .B1(n2471), .A0N(\register[12][28] ), .A1N(
        n2472), .Y(n488) );
  OAI2BB2XL U1355 ( .B0(n2294), .B1(n2471), .A0N(\register[12][29] ), .A1N(
        n2472), .Y(n489) );
  OAI2BB2XL U1356 ( .B0(n2292), .B1(n2471), .A0N(\register[12][30] ), .A1N(
        n2473), .Y(n490) );
  OAI2BB2XL U1357 ( .B0(n2290), .B1(n2471), .A0N(\register[12][31] ), .A1N(
        n2473), .Y(n491) );
  OAI2BB2XL U1358 ( .B0(n2307), .B1(n2461), .A0N(\register[14][23] ), .A1N(
        n2461), .Y(n547) );
  OAI2BB2XL U1359 ( .B0(n2303), .B1(n2461), .A0N(\register[14][25] ), .A1N(
        n2462), .Y(n549) );
  OAI2BB2XL U1360 ( .B0(n2301), .B1(n2461), .A0N(\register[14][26] ), .A1N(
        n2462), .Y(n550) );
  OAI2BB2XL U1361 ( .B0(n2299), .B1(n2461), .A0N(\register[14][27] ), .A1N(
        n2462), .Y(n551) );
  OAI2BB2XL U1362 ( .B0(n2296), .B1(n2461), .A0N(\register[14][28] ), .A1N(
        n2462), .Y(n552) );
  OAI2BB2XL U1363 ( .B0(n2294), .B1(n2461), .A0N(\register[14][29] ), .A1N(
        n2462), .Y(n553) );
  OAI2BB2XL U1364 ( .B0(n2292), .B1(n2461), .A0N(\register[14][30] ), .A1N(
        n2458), .Y(n554) );
  OAI2BB2XL U1365 ( .B0(n2290), .B1(n2461), .A0N(\register[14][31] ), .A1N(
        n2458), .Y(n555) );
  OAI2BB2XL U1366 ( .B0(n2307), .B1(n2426), .A0N(\register[20][23] ), .A1N(
        n2426), .Y(n739) );
  OAI2BB2XL U1367 ( .B0(n2303), .B1(n2426), .A0N(\register[20][25] ), .A1N(
        n2427), .Y(n741) );
  OAI2BB2XL U1368 ( .B0(n2301), .B1(n2426), .A0N(\register[20][26] ), .A1N(
        n2427), .Y(n742) );
  OAI2BB2XL U1369 ( .B0(n2298), .B1(n2426), .A0N(\register[20][27] ), .A1N(
        n2427), .Y(n743) );
  OAI2BB2XL U1370 ( .B0(n2296), .B1(n2426), .A0N(\register[20][28] ), .A1N(
        n2427), .Y(n744) );
  OAI2BB2XL U1371 ( .B0(n2294), .B1(n2426), .A0N(\register[20][29] ), .A1N(
        n2427), .Y(n745) );
  OAI2BB2XL U1372 ( .B0(n2292), .B1(n2426), .A0N(\register[20][30] ), .A1N(
        n2424), .Y(n746) );
  OAI2BB2XL U1373 ( .B0(n2290), .B1(n2426), .A0N(\register[20][31] ), .A1N(
        n2424), .Y(n747) );
  OAI2BB2XL U1374 ( .B0(n2307), .B1(n2416), .A0N(\register[22][23] ), .A1N(
        n2416), .Y(n803) );
  OAI2BB2XL U1375 ( .B0(n2303), .B1(n2416), .A0N(\register[22][25] ), .A1N(
        n2417), .Y(n805) );
  OAI2BB2XL U1376 ( .B0(n2301), .B1(n2416), .A0N(\register[22][26] ), .A1N(
        n2417), .Y(n806) );
  OAI2BB2XL U1377 ( .B0(n2298), .B1(n2416), .A0N(\register[22][27] ), .A1N(
        n2417), .Y(n807) );
  OAI2BB2XL U1378 ( .B0(n2296), .B1(n2416), .A0N(\register[22][28] ), .A1N(
        n2417), .Y(n808) );
  OAI2BB2XL U1379 ( .B0(n2294), .B1(n2416), .A0N(\register[22][29] ), .A1N(
        n2417), .Y(n809) );
  OAI2BB2XL U1380 ( .B0(n2292), .B1(n2416), .A0N(\register[22][30] ), .A1N(
        n2413), .Y(n810) );
  OAI2BB2XL U1381 ( .B0(n2290), .B1(n2416), .A0N(\register[22][31] ), .A1N(
        n2413), .Y(n811) );
  OAI2BB2XL U1382 ( .B0(n2307), .B1(n2383), .A0N(\register[28][23] ), .A1N(
        n2383), .Y(n995) );
  OAI2BB2XL U1383 ( .B0(n2303), .B1(n2383), .A0N(\register[28][25] ), .A1N(
        n2384), .Y(n997) );
  OAI2BB2XL U1384 ( .B0(n2301), .B1(n2383), .A0N(\register[28][26] ), .A1N(
        n2384), .Y(n998) );
  OAI2BB2XL U1385 ( .B0(n2298), .B1(n2383), .A0N(\register[28][27] ), .A1N(
        n2384), .Y(n999) );
  OAI2BB2XL U1386 ( .B0(n2296), .B1(n2383), .A0N(\register[28][28] ), .A1N(
        n2384), .Y(n1000) );
  OAI2BB2XL U1387 ( .B0(n2294), .B1(n2383), .A0N(\register[28][29] ), .A1N(
        n2384), .Y(n1001) );
  OAI2BB2XL U1388 ( .B0(n2292), .B1(n2383), .A0N(\register[28][30] ), .A1N(
        n2385), .Y(n1002) );
  OAI2BB2XL U1389 ( .B0(n2290), .B1(n2383), .A0N(\register[28][31] ), .A1N(
        n2385), .Y(n1003) );
  OAI2BB2XL U1390 ( .B0(n2307), .B1(n2374), .A0N(\register[30][23] ), .A1N(
        n2374), .Y(n1059) );
  OAI2BB2XL U1391 ( .B0(n2303), .B1(n2374), .A0N(\register[30][25] ), .A1N(
        n2375), .Y(n1061) );
  OAI2BB2XL U1392 ( .B0(n2301), .B1(n2374), .A0N(\register[30][26] ), .A1N(
        n2375), .Y(n1062) );
  OAI2BB2XL U1393 ( .B0(n2298), .B1(n2374), .A0N(\register[30][27] ), .A1N(
        n2375), .Y(n1063) );
  OAI2BB2XL U1394 ( .B0(n2296), .B1(n2374), .A0N(\register[30][28] ), .A1N(
        n2375), .Y(n1064) );
  OAI2BB2XL U1395 ( .B0(n2294), .B1(n2374), .A0N(\register[30][29] ), .A1N(
        n2375), .Y(n1065) );
  OAI2BB2XL U1396 ( .B0(n2292), .B1(n2374), .A0N(\register[30][30] ), .A1N(
        n2371), .Y(n1066) );
  OAI2BB2XL U1397 ( .B0(n2290), .B1(n2374), .A0N(\register[30][31] ), .A1N(
        n2371), .Y(n1067) );
  OAI2BB2XL U1398 ( .B0(n2308), .B1(n2525), .A0N(\register[2][23] ), .A1N(
        n2525), .Y(n163) );
  OAI2BB2XL U1399 ( .B0(n2304), .B1(n2525), .A0N(\register[2][25] ), .A1N(
        n2526), .Y(n165) );
  OAI2BB2XL U1400 ( .B0(n2302), .B1(n2525), .A0N(\register[2][26] ), .A1N(
        n2526), .Y(n166) );
  OAI2BB2XL U1401 ( .B0(n2300), .B1(n2525), .A0N(\register[2][27] ), .A1N(
        n2526), .Y(n167) );
  OAI2BB2XL U1402 ( .B0(n2297), .B1(n2525), .A0N(\register[2][28] ), .A1N(
        n2526), .Y(n168) );
  OAI2BB2XL U1403 ( .B0(n2295), .B1(n2525), .A0N(\register[2][29] ), .A1N(
        n2526), .Y(n169) );
  OAI2BB2XL U1404 ( .B0(n2293), .B1(n2525), .A0N(\register[2][30] ), .A1N(
        n2522), .Y(n170) );
  OAI2BB2XL U1405 ( .B0(n2291), .B1(n2525), .A0N(\register[2][31] ), .A1N(
        n2522), .Y(n171) );
  OAI2BB2XL U1406 ( .B0(n2307), .B1(n2484), .A0N(\register[10][23] ), .A1N(
        n2484), .Y(n419) );
  OAI2BB2XL U1407 ( .B0(n2303), .B1(n2484), .A0N(\register[10][25] ), .A1N(
        n2485), .Y(n421) );
  OAI2BB2XL U1408 ( .B0(n2301), .B1(n2484), .A0N(\register[10][26] ), .A1N(
        n2485), .Y(n422) );
  OAI2BB2XL U1409 ( .B0(n2299), .B1(n2484), .A0N(\register[10][27] ), .A1N(
        n2485), .Y(n423) );
  OAI2BB2XL U1410 ( .B0(n2296), .B1(n2484), .A0N(\register[10][28] ), .A1N(
        n2485), .Y(n424) );
  OAI2BB2XL U1411 ( .B0(n2294), .B1(n2484), .A0N(\register[10][29] ), .A1N(
        n2485), .Y(n425) );
  OAI2BB2XL U1412 ( .B0(n2292), .B1(n2484), .A0N(\register[10][30] ), .A1N(
        n2481), .Y(n426) );
  OAI2BB2XL U1413 ( .B0(n2290), .B1(n2484), .A0N(\register[10][31] ), .A1N(
        n2481), .Y(n427) );
  OAI2BB2XL U1414 ( .B0(n2307), .B1(n2438), .A0N(\register[18][23] ), .A1N(
        n2438), .Y(n675) );
  OAI2BB2XL U1415 ( .B0(n2303), .B1(n2438), .A0N(\register[18][25] ), .A1N(
        n2439), .Y(n677) );
  OAI2BB2XL U1416 ( .B0(n2301), .B1(n2438), .A0N(\register[18][26] ), .A1N(
        n2439), .Y(n678) );
  OAI2BB2XL U1417 ( .B0(n2299), .B1(n2438), .A0N(\register[18][27] ), .A1N(
        n2439), .Y(n679) );
  OAI2BB2XL U1418 ( .B0(n2296), .B1(n2438), .A0N(\register[18][28] ), .A1N(
        n2439), .Y(n680) );
  OAI2BB2XL U1419 ( .B0(n2294), .B1(n2438), .A0N(\register[18][29] ), .A1N(
        n2439), .Y(n681) );
  OAI2BB2XL U1420 ( .B0(n2292), .B1(n2438), .A0N(\register[18][30] ), .A1N(
        n2435), .Y(n682) );
  OAI2BB2XL U1421 ( .B0(n2290), .B1(n2438), .A0N(\register[18][31] ), .A1N(
        n2435), .Y(n683) );
  OAI2BB2XL U1422 ( .B0(n2307), .B1(n2394), .A0N(\register[26][23] ), .A1N(
        n2394), .Y(n931) );
  OAI2BB2XL U1423 ( .B0(n2303), .B1(n2394), .A0N(\register[26][25] ), .A1N(
        n2395), .Y(n933) );
  OAI2BB2XL U1424 ( .B0(n2301), .B1(n2394), .A0N(\register[26][26] ), .A1N(
        n2395), .Y(n934) );
  OAI2BB2XL U1425 ( .B0(n2298), .B1(n2394), .A0N(\register[26][27] ), .A1N(
        n2395), .Y(n935) );
  OAI2BB2XL U1426 ( .B0(n2296), .B1(n2394), .A0N(\register[26][28] ), .A1N(
        n2395), .Y(n936) );
  OAI2BB2XL U1427 ( .B0(n2294), .B1(n2394), .A0N(\register[26][29] ), .A1N(
        n2395), .Y(n937) );
  OAI2BB2XL U1428 ( .B0(n2292), .B1(n2394), .A0N(\register[26][30] ), .A1N(
        n2391), .Y(n938) );
  OAI2BB2XL U1429 ( .B0(n2290), .B1(n2394), .A0N(\register[26][31] ), .A1N(
        n2391), .Y(n939) );
  OAI2BB2XL U1430 ( .B0(n2308), .B1(n2500), .A0N(\register[7][23] ), .A1N(
        n2500), .Y(n323) );
  OAI2BB2XL U1431 ( .B0(n2304), .B1(n2500), .A0N(\register[7][25] ), .A1N(
        n2501), .Y(n325) );
  OAI2BB2XL U1432 ( .B0(n2302), .B1(n2500), .A0N(\register[7][26] ), .A1N(
        n2501), .Y(n326) );
  OAI2BB2XL U1433 ( .B0(n2300), .B1(n2500), .A0N(\register[7][27] ), .A1N(
        n2501), .Y(n327) );
  OAI2BB2XL U1434 ( .B0(n2297), .B1(n2500), .A0N(\register[7][28] ), .A1N(
        n2501), .Y(n328) );
  OAI2BB2XL U1435 ( .B0(n2295), .B1(n2500), .A0N(\register[7][29] ), .A1N(
        n2501), .Y(n329) );
  OAI2BB2XL U1436 ( .B0(n2293), .B1(n2500), .A0N(\register[7][30] ), .A1N(
        n2498), .Y(n330) );
  OAI2BB2XL U1437 ( .B0(n2291), .B1(n2500), .A0N(\register[7][31] ), .A1N(
        n2499), .Y(n331) );
  OAI2BB2XL U1438 ( .B0(n2307), .B1(n2455), .A0N(\register[15][23] ), .A1N(
        n2455), .Y(n579) );
  OAI2BB2XL U1439 ( .B0(n2303), .B1(n2455), .A0N(\register[15][25] ), .A1N(
        n2456), .Y(n581) );
  OAI2BB2XL U1440 ( .B0(n2301), .B1(n2455), .A0N(\register[15][26] ), .A1N(
        n2456), .Y(n582) );
  OAI2BB2XL U1441 ( .B0(n2299), .B1(n2455), .A0N(\register[15][27] ), .A1N(
        n2456), .Y(n583) );
  OAI2BB2XL U1442 ( .B0(n2296), .B1(n2455), .A0N(\register[15][28] ), .A1N(
        n2456), .Y(n584) );
  OAI2BB2XL U1443 ( .B0(n2294), .B1(n2455), .A0N(\register[15][29] ), .A1N(
        n2456), .Y(n585) );
  OAI2BB2XL U1444 ( .B0(n2292), .B1(n2455), .A0N(\register[15][30] ), .A1N(
        n2453), .Y(n586) );
  OAI2BB2XL U1445 ( .B0(n2290), .B1(n2455), .A0N(\register[15][31] ), .A1N(
        n2454), .Y(n587) );
  OAI2BB2XL U1446 ( .B0(n2307), .B1(n2409), .A0N(\register[23][23] ), .A1N(
        n2409), .Y(n835) );
  OAI2BB2XL U1447 ( .B0(n2303), .B1(n2409), .A0N(\register[23][25] ), .A1N(
        n2410), .Y(n837) );
  OAI2BB2XL U1448 ( .B0(n2301), .B1(n2409), .A0N(\register[23][26] ), .A1N(
        n2410), .Y(n838) );
  OAI2BB2XL U1449 ( .B0(n2298), .B1(n2409), .A0N(\register[23][27] ), .A1N(
        n2410), .Y(n839) );
  OAI2BB2XL U1450 ( .B0(n2296), .B1(n2409), .A0N(\register[23][28] ), .A1N(
        n2410), .Y(n840) );
  OAI2BB2XL U1451 ( .B0(n2294), .B1(n2409), .A0N(\register[23][29] ), .A1N(
        n2410), .Y(n841) );
  OAI2BB2XL U1452 ( .B0(n2292), .B1(n2409), .A0N(\register[23][30] ), .A1N(
        n2411), .Y(n842) );
  OAI2BB2XL U1453 ( .B0(n2290), .B1(n2409), .A0N(\register[23][31] ), .A1N(
        n2411), .Y(n843) );
  OAI2BB2XL U1454 ( .B0(n2307), .B1(n2368), .A0N(\register[31][23] ), .A1N(
        n2368), .Y(n1091) );
  OAI2BB2XL U1455 ( .B0(n2303), .B1(n2368), .A0N(\register[31][25] ), .A1N(
        n2369), .Y(n1093) );
  OAI2BB2XL U1456 ( .B0(n2301), .B1(n2368), .A0N(\register[31][26] ), .A1N(
        n2369), .Y(n1094) );
  OAI2BB2XL U1457 ( .B0(n2298), .B1(n2368), .A0N(\register[31][27] ), .A1N(
        n2369), .Y(n1095) );
  OAI2BB2XL U1458 ( .B0(n2296), .B1(n2368), .A0N(\register[31][28] ), .A1N(
        n2369), .Y(n1096) );
  OAI2BB2XL U1459 ( .B0(n2294), .B1(n2368), .A0N(\register[31][29] ), .A1N(
        n2369), .Y(n1097) );
  OAI2BB2XL U1460 ( .B0(n2292), .B1(n2368), .A0N(\register[31][30] ), .A1N(
        n2366), .Y(n1098) );
  OAI2BB2XL U1461 ( .B0(n2290), .B1(n2368), .A0N(\register[31][31] ), .A1N(
        n2367), .Y(n1099) );
  OAI2BB2XL U1462 ( .B0(n2308), .B1(n2511), .A0N(\register[5][23] ), .A1N(
        n2511), .Y(n259) );
  OAI2BB2XL U1463 ( .B0(n2304), .B1(n2511), .A0N(\register[5][25] ), .A1N(
        n2512), .Y(n261) );
  OAI2BB2XL U1464 ( .B0(n2302), .B1(n2511), .A0N(\register[5][26] ), .A1N(
        n2512), .Y(n262) );
  OAI2BB2XL U1465 ( .B0(n2300), .B1(n2511), .A0N(\register[5][27] ), .A1N(
        n2512), .Y(n263) );
  OAI2BB2XL U1466 ( .B0(n2297), .B1(n2511), .A0N(\register[5][28] ), .A1N(
        n2512), .Y(n264) );
  OAI2BB2XL U1467 ( .B0(n2295), .B1(n2511), .A0N(\register[5][29] ), .A1N(
        n2512), .Y(n265) );
  OAI2BB2XL U1468 ( .B0(n2293), .B1(n2511), .A0N(\register[5][30] ), .A1N(
        n2509), .Y(n266) );
  OAI2BB2XL U1469 ( .B0(n2291), .B1(n2511), .A0N(\register[5][31] ), .A1N(
        n2510), .Y(n267) );
  OAI2BB2XL U1470 ( .B0(n2307), .B1(n2494), .A0N(\register[8][23] ), .A1N(
        n2494), .Y(n355) );
  OAI2BB2XL U1471 ( .B0(n2303), .B1(n2494), .A0N(\register[8][25] ), .A1N(
        n2495), .Y(n357) );
  OAI2BB2XL U1472 ( .B0(n2301), .B1(n2494), .A0N(\register[8][26] ), .A1N(
        n2495), .Y(n358) );
  OAI2BB2XL U1473 ( .B0(n2299), .B1(n2494), .A0N(\register[8][27] ), .A1N(
        n2495), .Y(n359) );
  OAI2BB2XL U1474 ( .B0(n2296), .B1(n2494), .A0N(\register[8][28] ), .A1N(
        n2495), .Y(n360) );
  OAI2BB2XL U1475 ( .B0(n2294), .B1(n2494), .A0N(\register[8][29] ), .A1N(
        n2495), .Y(n361) );
  OAI2BB2XL U1476 ( .B0(n2292), .B1(n2494), .A0N(\register[8][30] ), .A1N(
        n2492), .Y(n362) );
  OAI2BB2XL U1477 ( .B0(n2290), .B1(n2494), .A0N(\register[8][31] ), .A1N(
        n2493), .Y(n363) );
  OAI2BB2XL U1478 ( .B0(n2307), .B1(n2449), .A0N(\register[16][23] ), .A1N(
        n2449), .Y(n611) );
  OAI2BB2XL U1479 ( .B0(n2303), .B1(n2449), .A0N(\register[16][25] ), .A1N(
        n2450), .Y(n613) );
  OAI2BB2XL U1480 ( .B0(n2301), .B1(n2449), .A0N(\register[16][26] ), .A1N(
        n2450), .Y(n614) );
  OAI2BB2XL U1481 ( .B0(n2299), .B1(n2449), .A0N(\register[16][27] ), .A1N(
        n2450), .Y(n615) );
  OAI2BB2XL U1482 ( .B0(n2296), .B1(n2449), .A0N(\register[16][28] ), .A1N(
        n2450), .Y(n616) );
  OAI2BB2XL U1483 ( .B0(n2294), .B1(n2449), .A0N(\register[16][29] ), .A1N(
        n2450), .Y(n617) );
  OAI2BB2XL U1484 ( .B0(n2292), .B1(n2449), .A0N(\register[16][30] ), .A1N(
        n2446), .Y(n618) );
  OAI2BB2XL U1485 ( .B0(n2290), .B1(n2449), .A0N(\register[16][31] ), .A1N(
        n2446), .Y(n619) );
  OAI2BB2XL U1486 ( .B0(n2308), .B1(n2404), .A0N(\register[24][23] ), .A1N(
        n2404), .Y(n867) );
  OAI2BB2XL U1487 ( .B0(n2304), .B1(n2404), .A0N(\register[24][25] ), .A1N(
        n2405), .Y(n869) );
  OAI2BB2XL U1488 ( .B0(n2302), .B1(n2404), .A0N(\register[24][26] ), .A1N(
        n2405), .Y(n870) );
  OAI2BB2XL U1489 ( .B0(n2298), .B1(n2404), .A0N(\register[24][27] ), .A1N(
        n2405), .Y(n871) );
  OAI2BB2XL U1490 ( .B0(n2297), .B1(n2404), .A0N(\register[24][28] ), .A1N(
        n2405), .Y(n872) );
  OAI2BB2XL U1491 ( .B0(n2295), .B1(n2404), .A0N(\register[24][29] ), .A1N(
        n2405), .Y(n873) );
  OAI2BB2XL U1492 ( .B0(n2293), .B1(n2404), .A0N(\register[24][30] ), .A1N(
        n2403), .Y(n874) );
  OAI2BB2XL U1493 ( .B0(n2291), .B1(n2404), .A0N(\register[24][31] ), .A1N(
        n2402), .Y(n875) );
  OAI2BB2XL U1494 ( .B0(n2307), .B1(n2467), .A0N(\register[13][23] ), .A1N(
        n2467), .Y(n515) );
  OAI2BB2XL U1495 ( .B0(n2308), .B1(n2421), .A0N(\register[21][23] ), .A1N(
        n2421), .Y(n771) );
  OAI2BB2XL U1496 ( .B0(n2308), .B1(n2379), .A0N(\register[29][23] ), .A1N(
        n2379), .Y(n1027) );
  OAI2BB2XL U1497 ( .B0(n2303), .B1(n2467), .A0N(\register[13][25] ), .A1N(
        n2468), .Y(n517) );
  OAI2BB2XL U1498 ( .B0(n2301), .B1(n2467), .A0N(\register[13][26] ), .A1N(
        n2468), .Y(n518) );
  OAI2BB2XL U1499 ( .B0(n2299), .B1(n2467), .A0N(\register[13][27] ), .A1N(
        n2468), .Y(n519) );
  OAI2BB2XL U1500 ( .B0(n2296), .B1(n2467), .A0N(\register[13][28] ), .A1N(
        n2468), .Y(n520) );
  OAI2BB2XL U1501 ( .B0(n2294), .B1(n2467), .A0N(\register[13][29] ), .A1N(
        n2468), .Y(n521) );
  OAI2BB2XL U1502 ( .B0(n2304), .B1(n2421), .A0N(\register[21][25] ), .A1N(
        n2422), .Y(n773) );
  OAI2BB2XL U1503 ( .B0(n2302), .B1(n2421), .A0N(\register[21][26] ), .A1N(
        n2422), .Y(n774) );
  OAI2BB2XL U1504 ( .B0(n2298), .B1(n2421), .A0N(\register[21][27] ), .A1N(
        n2422), .Y(n775) );
  OAI2BB2XL U1505 ( .B0(n2297), .B1(n2421), .A0N(\register[21][28] ), .A1N(
        n2422), .Y(n776) );
  OAI2BB2XL U1506 ( .B0(n2295), .B1(n2421), .A0N(\register[21][29] ), .A1N(
        n2422), .Y(n777) );
  OAI2BB2XL U1507 ( .B0(n2304), .B1(n2379), .A0N(\register[29][25] ), .A1N(
        n2380), .Y(n1029) );
  OAI2BB2XL U1508 ( .B0(n2302), .B1(n2379), .A0N(\register[29][26] ), .A1N(
        n2380), .Y(n1030) );
  OAI2BB2XL U1509 ( .B0(n2298), .B1(n2379), .A0N(\register[29][27] ), .A1N(
        n2380), .Y(n1031) );
  OAI2BB2XL U1510 ( .B0(n2297), .B1(n2379), .A0N(\register[29][28] ), .A1N(
        n2380), .Y(n1032) );
  OAI2BB2XL U1511 ( .B0(n2295), .B1(n2379), .A0N(\register[29][29] ), .A1N(
        n2380), .Y(n1033) );
  OAI2BB2XL U1512 ( .B0(n2292), .B1(n2467), .A0N(\register[13][30] ), .A1N(
        n2465), .Y(n522) );
  OAI2BB2XL U1513 ( .B0(n2290), .B1(n2467), .A0N(\register[13][31] ), .A1N(
        n2466), .Y(n523) );
  OAI2BB2XL U1514 ( .B0(n2293), .B1(n2421), .A0N(\register[21][30] ), .A1N(
        n2423), .Y(n778) );
  OAI2BB2XL U1515 ( .B0(n2291), .B1(n2421), .A0N(\register[21][31] ), .A1N(
        n2423), .Y(n779) );
  OAI2BB2XL U1516 ( .B0(n2293), .B1(n2379), .A0N(\register[29][30] ), .A1N(
        n2377), .Y(n1034) );
  OAI2BB2XL U1517 ( .B0(n2291), .B1(n2379), .A0N(\register[29][31] ), .A1N(
        n2378), .Y(n1035) );
  OAI2BB2XL U1518 ( .B0(n2362), .B1(n2470), .A0N(\register[12][0] ), .A1N(
        n2473), .Y(n460) );
  OAI2BB2XL U1519 ( .B0(n2361), .B1(n2469), .A0N(\register[12][1] ), .A1N(
        n2473), .Y(n461) );
  OAI2BB2XL U1520 ( .B0(n2359), .B1(n2469), .A0N(\register[12][2] ), .A1N(
        n2473), .Y(n462) );
  OAI2BB2XL U1521 ( .B0(n2356), .B1(n2469), .A0N(\register[12][3] ), .A1N(
        n2472), .Y(n463) );
  OAI2BB2XL U1522 ( .B0(n2354), .B1(n2469), .A0N(\register[12][4] ), .A1N(
        n2473), .Y(n464) );
  OAI2BB2XL U1523 ( .B0(n2351), .B1(n2469), .A0N(\register[12][5] ), .A1N(
        n2472), .Y(n465) );
  OAI2BB2XL U1524 ( .B0(n2349), .B1(n2469), .A0N(\register[12][6] ), .A1N(
        n2472), .Y(n466) );
  OAI2BB2XL U1525 ( .B0(n2346), .B1(n2469), .A0N(\register[12][7] ), .A1N(
        n2472), .Y(n467) );
  OAI2BB2XL U1526 ( .B0(n2344), .B1(n2469), .A0N(\register[12][8] ), .A1N(
        n2472), .Y(n468) );
  OAI2BB2XL U1527 ( .B0(n2342), .B1(n2469), .A0N(\register[12][9] ), .A1N(
        n2472), .Y(n469) );
  OAI2BB2XL U1528 ( .B0(n2339), .B1(n2469), .A0N(\register[12][10] ), .A1N(
        n2472), .Y(n470) );
  OAI2BB2XL U1529 ( .B0(n2337), .B1(n2469), .A0N(\register[12][11] ), .A1N(
        n2472), .Y(n471) );
  OAI2BB2XL U1530 ( .B0(n2335), .B1(n2469), .A0N(\register[12][12] ), .A1N(
        n2472), .Y(n472) );
  OAI2BB2XL U1531 ( .B0(n2332), .B1(n2470), .A0N(\register[12][13] ), .A1N(
        n2472), .Y(n473) );
  OAI2BB2XL U1532 ( .B0(n2330), .B1(n2470), .A0N(\register[12][14] ), .A1N(
        n2472), .Y(n474) );
  OAI2BB2XL U1533 ( .B0(n2327), .B1(n2470), .A0N(\register[12][15] ), .A1N(
        n2471), .Y(n475) );
  OAI2BB2XL U1534 ( .B0(n2324), .B1(n2470), .A0N(\register[12][16] ), .A1N(
        n2472), .Y(n476) );
  OAI2BB2XL U1535 ( .B0(n2322), .B1(n2470), .A0N(\register[12][17] ), .A1N(
        n2471), .Y(n477) );
  OAI2BB2XL U1536 ( .B0(n2319), .B1(n2470), .A0N(\register[12][18] ), .A1N(
        n2471), .Y(n478) );
  OAI2BB2XL U1537 ( .B0(n2316), .B1(n2470), .A0N(\register[12][19] ), .A1N(
        n2471), .Y(n479) );
  OAI2BB2XL U1538 ( .B0(n2314), .B1(n2470), .A0N(\register[12][20] ), .A1N(
        n2471), .Y(n480) );
  OAI2BB2XL U1539 ( .B0(n2312), .B1(n2470), .A0N(\register[12][21] ), .A1N(
        n2471), .Y(n481) );
  OAI2BB2XL U1540 ( .B0(n2310), .B1(n2470), .A0N(\register[12][22] ), .A1N(
        n2472), .Y(n482) );
  OAI2BB2XL U1541 ( .B0(n2305), .B1(n2470), .A0N(\register[12][24] ), .A1N(
        n2472), .Y(n484) );
  OAI2BB2XL U1542 ( .B0(n2362), .B1(n2460), .A0N(\register[14][0] ), .A1N(
        n2458), .Y(n524) );
  OAI2BB2XL U1543 ( .B0(n2361), .B1(n2459), .A0N(\register[14][1] ), .A1N(
        n2458), .Y(n525) );
  OAI2BB2XL U1544 ( .B0(n2359), .B1(n2459), .A0N(\register[14][2] ), .A1N(
        n2458), .Y(n526) );
  OAI2BB2XL U1545 ( .B0(n2356), .B1(n2459), .A0N(\register[14][3] ), .A1N(
        n2462), .Y(n527) );
  OAI2BB2XL U1546 ( .B0(n2354), .B1(n2459), .A0N(\register[14][4] ), .A1N(
        n2458), .Y(n528) );
  OAI2BB2XL U1547 ( .B0(n2351), .B1(n2459), .A0N(\register[14][5] ), .A1N(
        n2462), .Y(n529) );
  OAI2BB2XL U1548 ( .B0(n2349), .B1(n2459), .A0N(\register[14][6] ), .A1N(
        n2462), .Y(n530) );
  OAI2BB2XL U1549 ( .B0(n2346), .B1(n2459), .A0N(\register[14][7] ), .A1N(
        n2462), .Y(n531) );
  OAI2BB2XL U1550 ( .B0(n2344), .B1(n2459), .A0N(\register[14][8] ), .A1N(
        n2462), .Y(n532) );
  OAI2BB2XL U1551 ( .B0(n2342), .B1(n2459), .A0N(\register[14][9] ), .A1N(
        n2462), .Y(n533) );
  OAI2BB2XL U1552 ( .B0(n2339), .B1(n2459), .A0N(\register[14][10] ), .A1N(
        n2462), .Y(n534) );
  OAI2BB2XL U1553 ( .B0(n2337), .B1(n2459), .A0N(\register[14][11] ), .A1N(
        n2462), .Y(n535) );
  OAI2BB2XL U1554 ( .B0(n2335), .B1(n2459), .A0N(\register[14][12] ), .A1N(
        n2462), .Y(n536) );
  OAI2BB2XL U1555 ( .B0(n2332), .B1(n2460), .A0N(\register[14][13] ), .A1N(
        n2462), .Y(n537) );
  OAI2BB2XL U1556 ( .B0(n2330), .B1(n2460), .A0N(\register[14][14] ), .A1N(
        n2462), .Y(n538) );
  OAI2BB2XL U1557 ( .B0(n2327), .B1(n2460), .A0N(\register[14][15] ), .A1N(
        n2461), .Y(n539) );
  OAI2BB2XL U1558 ( .B0(n2324), .B1(n2460), .A0N(\register[14][16] ), .A1N(
        n2462), .Y(n540) );
  OAI2BB2XL U1559 ( .B0(n2322), .B1(n2460), .A0N(\register[14][17] ), .A1N(
        n2461), .Y(n541) );
  OAI2BB2XL U1560 ( .B0(n2319), .B1(n2460), .A0N(\register[14][18] ), .A1N(
        n2461), .Y(n542) );
  OAI2BB2XL U1561 ( .B0(n2316), .B1(n2460), .A0N(\register[14][19] ), .A1N(
        n2461), .Y(n543) );
  OAI2BB2XL U1562 ( .B0(n2314), .B1(n2460), .A0N(\register[14][20] ), .A1N(
        n2461), .Y(n544) );
  OAI2BB2XL U1563 ( .B0(n2312), .B1(n2460), .A0N(\register[14][21] ), .A1N(
        n2461), .Y(n545) );
  OAI2BB2XL U1564 ( .B0(n2310), .B1(n2460), .A0N(\register[14][22] ), .A1N(
        n2462), .Y(n546) );
  OAI2BB2XL U1565 ( .B0(n2305), .B1(n2460), .A0N(\register[14][24] ), .A1N(
        n2462), .Y(n548) );
  OAI2BB2XL U1566 ( .B0(n2362), .B1(n2425), .A0N(\register[20][0] ), .A1N(
        n2424), .Y(n716) );
  OAI2BB2XL U1567 ( .B0(n2360), .B1(n2424), .A0N(\register[20][1] ), .A1N(
        n2424), .Y(n717) );
  OAI2BB2XL U1568 ( .B0(n2358), .B1(n2424), .A0N(\register[20][2] ), .A1N(
        n2424), .Y(n718) );
  OAI2BB2XL U1569 ( .B0(n2355), .B1(n2424), .A0N(\register[20][3] ), .A1N(
        n2427), .Y(n719) );
  OAI2BB2XL U1570 ( .B0(n2353), .B1(n2425), .A0N(\register[20][4] ), .A1N(
        n2424), .Y(n720) );
  OAI2BB2XL U1571 ( .B0(n2351), .B1(n2424), .A0N(\register[20][5] ), .A1N(
        n2427), .Y(n721) );
  OAI2BB2XL U1572 ( .B0(n2348), .B1(n2425), .A0N(\register[20][6] ), .A1N(
        n2427), .Y(n722) );
  OAI2BB2XL U1573 ( .B0(n2346), .B1(n2424), .A0N(\register[20][7] ), .A1N(
        n2427), .Y(n723) );
  OAI2BB2XL U1574 ( .B0(n2344), .B1(n2424), .A0N(\register[20][8] ), .A1N(
        n2427), .Y(n724) );
  OAI2BB2XL U1575 ( .B0(n2341), .B1(n2425), .A0N(\register[20][9] ), .A1N(
        n2427), .Y(n725) );
  OAI2BB2XL U1576 ( .B0(n2339), .B1(n2424), .A0N(\register[20][10] ), .A1N(
        n2427), .Y(n726) );
  OAI2BB2XL U1577 ( .B0(n2337), .B1(n2424), .A0N(\register[20][11] ), .A1N(
        n2427), .Y(n727) );
  OAI2BB2XL U1578 ( .B0(n2334), .B1(n2425), .A0N(\register[20][12] ), .A1N(
        n2427), .Y(n728) );
  OAI2BB2XL U1579 ( .B0(n2332), .B1(n2425), .A0N(\register[20][13] ), .A1N(
        n2427), .Y(n729) );
  OAI2BB2XL U1580 ( .B0(n2329), .B1(n2425), .A0N(\register[20][14] ), .A1N(
        n2427), .Y(n730) );
  OAI2BB2XL U1581 ( .B0(n2326), .B1(n2425), .A0N(\register[20][15] ), .A1N(
        n2426), .Y(n731) );
  OAI2BB2XL U1582 ( .B0(n2324), .B1(n2425), .A0N(\register[20][16] ), .A1N(
        n2427), .Y(n732) );
  OAI2BB2XL U1583 ( .B0(n2321), .B1(n2425), .A0N(\register[20][17] ), .A1N(
        n2426), .Y(n733) );
  OAI2BB2XL U1584 ( .B0(n2318), .B1(n2425), .A0N(\register[20][18] ), .A1N(
        n2426), .Y(n734) );
  OAI2BB2XL U1585 ( .B0(n2316), .B1(n2425), .A0N(\register[20][19] ), .A1N(
        n2426), .Y(n735) );
  OAI2BB2XL U1586 ( .B0(n2314), .B1(n2425), .A0N(\register[20][20] ), .A1N(
        n2426), .Y(n736) );
  OAI2BB2XL U1587 ( .B0(n2312), .B1(n2425), .A0N(\register[20][21] ), .A1N(
        n2426), .Y(n737) );
  OAI2BB2XL U1588 ( .B0(n2309), .B1(n2425), .A0N(\register[20][22] ), .A1N(
        n2427), .Y(n738) );
  OAI2BB2XL U1589 ( .B0(n2305), .B1(n2425), .A0N(\register[20][24] ), .A1N(
        n2427), .Y(n740) );
  OAI2BB2XL U1590 ( .B0(n2362), .B1(n2415), .A0N(\register[22][0] ), .A1N(
        n2413), .Y(n780) );
  OAI2BB2XL U1591 ( .B0(n2360), .B1(n2414), .A0N(\register[22][1] ), .A1N(
        n2413), .Y(n781) );
  OAI2BB2XL U1592 ( .B0(n2358), .B1(n2414), .A0N(\register[22][2] ), .A1N(
        n2413), .Y(n782) );
  OAI2BB2XL U1593 ( .B0(n2355), .B1(n2414), .A0N(\register[22][3] ), .A1N(
        n2417), .Y(n783) );
  OAI2BB2XL U1594 ( .B0(n2353), .B1(n2414), .A0N(\register[22][4] ), .A1N(
        n2413), .Y(n784) );
  OAI2BB2XL U1595 ( .B0(n2351), .B1(n2414), .A0N(\register[22][5] ), .A1N(
        n2417), .Y(n785) );
  OAI2BB2XL U1596 ( .B0(n2348), .B1(n2414), .A0N(\register[22][6] ), .A1N(
        n2417), .Y(n786) );
  OAI2BB2XL U1597 ( .B0(n2346), .B1(n2414), .A0N(\register[22][7] ), .A1N(
        n2417), .Y(n787) );
  OAI2BB2XL U1598 ( .B0(n2344), .B1(n2414), .A0N(\register[22][8] ), .A1N(
        n2417), .Y(n788) );
  OAI2BB2XL U1599 ( .B0(n2341), .B1(n2414), .A0N(\register[22][9] ), .A1N(
        n2417), .Y(n789) );
  OAI2BB2XL U1600 ( .B0(n2339), .B1(n2414), .A0N(\register[22][10] ), .A1N(
        n2417), .Y(n790) );
  OAI2BB2XL U1601 ( .B0(n2337), .B1(n2414), .A0N(\register[22][11] ), .A1N(
        n2417), .Y(n791) );
  OAI2BB2XL U1602 ( .B0(n2334), .B1(n2414), .A0N(\register[22][12] ), .A1N(
        n2417), .Y(n792) );
  OAI2BB2XL U1603 ( .B0(n2332), .B1(n2415), .A0N(\register[22][13] ), .A1N(
        n2417), .Y(n793) );
  OAI2BB2XL U1604 ( .B0(n2329), .B1(n2415), .A0N(\register[22][14] ), .A1N(
        n2417), .Y(n794) );
  OAI2BB2XL U1605 ( .B0(n2326), .B1(n2415), .A0N(\register[22][15] ), .A1N(
        n2416), .Y(n795) );
  OAI2BB2XL U1606 ( .B0(n2324), .B1(n2415), .A0N(\register[22][16] ), .A1N(
        n2417), .Y(n796) );
  OAI2BB2XL U1607 ( .B0(n2321), .B1(n2415), .A0N(\register[22][17] ), .A1N(
        n2416), .Y(n797) );
  OAI2BB2XL U1608 ( .B0(n2318), .B1(n2415), .A0N(\register[22][18] ), .A1N(
        n2416), .Y(n798) );
  OAI2BB2XL U1609 ( .B0(n2316), .B1(n2415), .A0N(\register[22][19] ), .A1N(
        n2416), .Y(n799) );
  OAI2BB2XL U1610 ( .B0(n2314), .B1(n2415), .A0N(\register[22][20] ), .A1N(
        n2416), .Y(n800) );
  OAI2BB2XL U1611 ( .B0(n2312), .B1(n2415), .A0N(\register[22][21] ), .A1N(
        n2416), .Y(n801) );
  OAI2BB2XL U1612 ( .B0(n2309), .B1(n2415), .A0N(\register[22][22] ), .A1N(
        n2417), .Y(n802) );
  OAI2BB2XL U1613 ( .B0(n2305), .B1(n2415), .A0N(\register[22][24] ), .A1N(
        n2417), .Y(n804) );
  OAI2BB2XL U1614 ( .B0(n2362), .B1(n2382), .A0N(\register[28][0] ), .A1N(
        n2385), .Y(n972) );
  OAI2BB2XL U1615 ( .B0(n2360), .B1(n2381), .A0N(\register[28][1] ), .A1N(
        n2385), .Y(n973) );
  OAI2BB2XL U1616 ( .B0(n2358), .B1(n2381), .A0N(\register[28][2] ), .A1N(
        n2385), .Y(n974) );
  OAI2BB2XL U1617 ( .B0(n2355), .B1(n2381), .A0N(\register[28][3] ), .A1N(
        n2384), .Y(n975) );
  OAI2BB2XL U1618 ( .B0(n2353), .B1(n2381), .A0N(\register[28][4] ), .A1N(
        n2385), .Y(n976) );
  OAI2BB2XL U1619 ( .B0(n2351), .B1(n2381), .A0N(\register[28][5] ), .A1N(
        n2384), .Y(n977) );
  OAI2BB2XL U1620 ( .B0(n2348), .B1(n2381), .A0N(\register[28][6] ), .A1N(
        n2384), .Y(n978) );
  OAI2BB2XL U1621 ( .B0(n2346), .B1(n2381), .A0N(\register[28][7] ), .A1N(
        n2384), .Y(n979) );
  OAI2BB2XL U1622 ( .B0(n2344), .B1(n2381), .A0N(\register[28][8] ), .A1N(
        n2384), .Y(n980) );
  OAI2BB2XL U1623 ( .B0(n2341), .B1(n2381), .A0N(\register[28][9] ), .A1N(
        n2384), .Y(n981) );
  OAI2BB2XL U1624 ( .B0(n2339), .B1(n2381), .A0N(\register[28][10] ), .A1N(
        n2384), .Y(n982) );
  OAI2BB2XL U1625 ( .B0(n2337), .B1(n2381), .A0N(\register[28][11] ), .A1N(
        n2384), .Y(n983) );
  OAI2BB2XL U1626 ( .B0(n2334), .B1(n2381), .A0N(\register[28][12] ), .A1N(
        n2384), .Y(n984) );
  OAI2BB2XL U1627 ( .B0(n2332), .B1(n2382), .A0N(\register[28][13] ), .A1N(
        n2384), .Y(n985) );
  OAI2BB2XL U1628 ( .B0(n2329), .B1(n2382), .A0N(\register[28][14] ), .A1N(
        n2384), .Y(n986) );
  OAI2BB2XL U1629 ( .B0(n2326), .B1(n2382), .A0N(\register[28][15] ), .A1N(
        n2383), .Y(n987) );
  OAI2BB2XL U1630 ( .B0(n2324), .B1(n2382), .A0N(\register[28][16] ), .A1N(
        n2384), .Y(n988) );
  OAI2BB2XL U1631 ( .B0(n2321), .B1(n2382), .A0N(\register[28][17] ), .A1N(
        n2383), .Y(n989) );
  OAI2BB2XL U1632 ( .B0(n2318), .B1(n2382), .A0N(\register[28][18] ), .A1N(
        n2383), .Y(n990) );
  OAI2BB2XL U1633 ( .B0(n2316), .B1(n2382), .A0N(\register[28][19] ), .A1N(
        n2383), .Y(n991) );
  OAI2BB2XL U1634 ( .B0(n2314), .B1(n2382), .A0N(\register[28][20] ), .A1N(
        n2383), .Y(n992) );
  OAI2BB2XL U1635 ( .B0(n2312), .B1(n2382), .A0N(\register[28][21] ), .A1N(
        n2383), .Y(n993) );
  OAI2BB2XL U1636 ( .B0(n2309), .B1(n2382), .A0N(\register[28][22] ), .A1N(
        n2384), .Y(n994) );
  OAI2BB2XL U1637 ( .B0(n2305), .B1(n2382), .A0N(\register[28][24] ), .A1N(
        n2384), .Y(n996) );
  OAI2BB2XL U1638 ( .B0(n2362), .B1(n2373), .A0N(\register[30][0] ), .A1N(
        n2371), .Y(n1036) );
  OAI2BB2XL U1639 ( .B0(n2360), .B1(n2372), .A0N(\register[30][1] ), .A1N(
        n2371), .Y(n1037) );
  OAI2BB2XL U1640 ( .B0(n2358), .B1(n2372), .A0N(\register[30][2] ), .A1N(
        n2371), .Y(n1038) );
  OAI2BB2XL U1641 ( .B0(n2355), .B1(n2372), .A0N(\register[30][3] ), .A1N(
        n2375), .Y(n1039) );
  OAI2BB2XL U1642 ( .B0(n2353), .B1(n2372), .A0N(\register[30][4] ), .A1N(
        n2371), .Y(n1040) );
  OAI2BB2XL U1643 ( .B0(n2351), .B1(n2372), .A0N(\register[30][5] ), .A1N(
        n2375), .Y(n1041) );
  OAI2BB2XL U1644 ( .B0(n2348), .B1(n2372), .A0N(\register[30][6] ), .A1N(
        n2375), .Y(n1042) );
  OAI2BB2XL U1645 ( .B0(n2346), .B1(n2372), .A0N(\register[30][7] ), .A1N(
        n2375), .Y(n1043) );
  OAI2BB2XL U1646 ( .B0(n2344), .B1(n2372), .A0N(\register[30][8] ), .A1N(
        n2375), .Y(n1044) );
  OAI2BB2XL U1647 ( .B0(n2341), .B1(n2372), .A0N(\register[30][9] ), .A1N(
        n2375), .Y(n1045) );
  OAI2BB2XL U1648 ( .B0(n2339), .B1(n2372), .A0N(\register[30][10] ), .A1N(
        n2375), .Y(n1046) );
  OAI2BB2XL U1649 ( .B0(n2337), .B1(n2372), .A0N(\register[30][11] ), .A1N(
        n2375), .Y(n1047) );
  OAI2BB2XL U1650 ( .B0(n2334), .B1(n2372), .A0N(\register[30][12] ), .A1N(
        n2375), .Y(n1048) );
  OAI2BB2XL U1651 ( .B0(n2332), .B1(n2373), .A0N(\register[30][13] ), .A1N(
        n2375), .Y(n1049) );
  OAI2BB2XL U1652 ( .B0(n2329), .B1(n2373), .A0N(\register[30][14] ), .A1N(
        n2375), .Y(n1050) );
  OAI2BB2XL U1653 ( .B0(n2326), .B1(n2373), .A0N(\register[30][15] ), .A1N(
        n2374), .Y(n1051) );
  OAI2BB2XL U1654 ( .B0(n2324), .B1(n2373), .A0N(\register[30][16] ), .A1N(
        n2375), .Y(n1052) );
  OAI2BB2XL U1655 ( .B0(n2321), .B1(n2373), .A0N(\register[30][17] ), .A1N(
        n2374), .Y(n1053) );
  OAI2BB2XL U1656 ( .B0(n2318), .B1(n2373), .A0N(\register[30][18] ), .A1N(
        n2374), .Y(n1054) );
  OAI2BB2XL U1657 ( .B0(n2316), .B1(n2373), .A0N(\register[30][19] ), .A1N(
        n2374), .Y(n1055) );
  OAI2BB2XL U1658 ( .B0(n2314), .B1(n2373), .A0N(\register[30][20] ), .A1N(
        n2374), .Y(n1056) );
  OAI2BB2XL U1659 ( .B0(n2312), .B1(n2373), .A0N(\register[30][21] ), .A1N(
        n2374), .Y(n1057) );
  OAI2BB2XL U1660 ( .B0(n2309), .B1(n2373), .A0N(\register[30][22] ), .A1N(
        n2375), .Y(n1058) );
  OAI2BB2XL U1661 ( .B0(n2305), .B1(n2373), .A0N(\register[30][24] ), .A1N(
        n2375), .Y(n1060) );
  OAI2BB2XL U1662 ( .B0(n2362), .B1(n2483), .A0N(\register[10][0] ), .A1N(
        n2481), .Y(n396) );
  OAI2BB2XL U1663 ( .B0(n2361), .B1(n2482), .A0N(\register[10][1] ), .A1N(
        n2481), .Y(n397) );
  OAI2BB2XL U1664 ( .B0(n2359), .B1(n2482), .A0N(\register[10][2] ), .A1N(
        n2481), .Y(n398) );
  OAI2BB2XL U1665 ( .B0(n2356), .B1(n2482), .A0N(\register[10][3] ), .A1N(
        n2485), .Y(n399) );
  OAI2BB2XL U1666 ( .B0(n2354), .B1(n2482), .A0N(\register[10][4] ), .A1N(
        n2481), .Y(n400) );
  OAI2BB2XL U1667 ( .B0(n2351), .B1(n2482), .A0N(\register[10][5] ), .A1N(
        n2485), .Y(n401) );
  OAI2BB2XL U1668 ( .B0(n2349), .B1(n2482), .A0N(\register[10][6] ), .A1N(
        n2485), .Y(n402) );
  OAI2BB2XL U1669 ( .B0(n2346), .B1(n2482), .A0N(\register[10][7] ), .A1N(
        n2485), .Y(n403) );
  OAI2BB2XL U1670 ( .B0(n2344), .B1(n2482), .A0N(\register[10][8] ), .A1N(
        n2485), .Y(n404) );
  OAI2BB2XL U1671 ( .B0(n2342), .B1(n2482), .A0N(\register[10][9] ), .A1N(
        n2485), .Y(n405) );
  OAI2BB2XL U1672 ( .B0(n2339), .B1(n2482), .A0N(\register[10][10] ), .A1N(
        n2485), .Y(n406) );
  OAI2BB2XL U1673 ( .B0(n2337), .B1(n2482), .A0N(\register[10][11] ), .A1N(
        n2485), .Y(n407) );
  OAI2BB2XL U1674 ( .B0(n2335), .B1(n2482), .A0N(\register[10][12] ), .A1N(
        n2485), .Y(n408) );
  OAI2BB2XL U1675 ( .B0(n2332), .B1(n2483), .A0N(\register[10][13] ), .A1N(
        n2485), .Y(n409) );
  OAI2BB2XL U1676 ( .B0(n2330), .B1(n2483), .A0N(\register[10][14] ), .A1N(
        n2485), .Y(n410) );
  OAI2BB2XL U1677 ( .B0(n2327), .B1(n2483), .A0N(\register[10][15] ), .A1N(
        n2484), .Y(n411) );
  OAI2BB2XL U1678 ( .B0(n2324), .B1(n2483), .A0N(\register[10][16] ), .A1N(
        n2485), .Y(n412) );
  OAI2BB2XL U1679 ( .B0(n2322), .B1(n2483), .A0N(\register[10][17] ), .A1N(
        n2484), .Y(n413) );
  OAI2BB2XL U1680 ( .B0(n2319), .B1(n2483), .A0N(\register[10][18] ), .A1N(
        n2484), .Y(n414) );
  OAI2BB2XL U1681 ( .B0(n2316), .B1(n2483), .A0N(\register[10][19] ), .A1N(
        n2484), .Y(n415) );
  OAI2BB2XL U1682 ( .B0(n2314), .B1(n2483), .A0N(\register[10][20] ), .A1N(
        n2484), .Y(n416) );
  OAI2BB2XL U1683 ( .B0(n2312), .B1(n2483), .A0N(\register[10][21] ), .A1N(
        n2484), .Y(n417) );
  OAI2BB2XL U1684 ( .B0(n2310), .B1(n2483), .A0N(\register[10][22] ), .A1N(
        n2485), .Y(n418) );
  OAI2BB2XL U1685 ( .B0(n2305), .B1(n2483), .A0N(\register[10][24] ), .A1N(
        n2485), .Y(n420) );
  OAI2BB2XL U1686 ( .B0(n2362), .B1(n2437), .A0N(\register[18][0] ), .A1N(
        n2435), .Y(n652) );
  OAI2BB2XL U1687 ( .B0(n2361), .B1(n2436), .A0N(\register[18][1] ), .A1N(
        n2435), .Y(n653) );
  OAI2BB2XL U1688 ( .B0(n2359), .B1(n2436), .A0N(\register[18][2] ), .A1N(
        n2435), .Y(n654) );
  OAI2BB2XL U1689 ( .B0(n2356), .B1(n2436), .A0N(\register[18][3] ), .A1N(
        n2439), .Y(n655) );
  OAI2BB2XL U1690 ( .B0(n2354), .B1(n2436), .A0N(\register[18][4] ), .A1N(
        n2435), .Y(n656) );
  OAI2BB2XL U1691 ( .B0(n2351), .B1(n2436), .A0N(\register[18][5] ), .A1N(
        n2439), .Y(n657) );
  OAI2BB2XL U1692 ( .B0(n2349), .B1(n2436), .A0N(\register[18][6] ), .A1N(
        n2439), .Y(n658) );
  OAI2BB2XL U1693 ( .B0(n2346), .B1(n2436), .A0N(\register[18][7] ), .A1N(
        n2439), .Y(n659) );
  OAI2BB2XL U1694 ( .B0(n2344), .B1(n2436), .A0N(\register[18][8] ), .A1N(
        n2439), .Y(n660) );
  OAI2BB2XL U1695 ( .B0(n2342), .B1(n2436), .A0N(\register[18][9] ), .A1N(
        n2439), .Y(n661) );
  OAI2BB2XL U1696 ( .B0(n2339), .B1(n2436), .A0N(\register[18][10] ), .A1N(
        n2439), .Y(n662) );
  OAI2BB2XL U1697 ( .B0(n2337), .B1(n2436), .A0N(\register[18][11] ), .A1N(
        n2439), .Y(n663) );
  OAI2BB2XL U1698 ( .B0(n2335), .B1(n2436), .A0N(\register[18][12] ), .A1N(
        n2439), .Y(n664) );
  OAI2BB2XL U1699 ( .B0(n2332), .B1(n2437), .A0N(\register[18][13] ), .A1N(
        n2439), .Y(n665) );
  OAI2BB2XL U1700 ( .B0(n2330), .B1(n2437), .A0N(\register[18][14] ), .A1N(
        n2439), .Y(n666) );
  OAI2BB2XL U1701 ( .B0(n2327), .B1(n2437), .A0N(\register[18][15] ), .A1N(
        n2438), .Y(n667) );
  OAI2BB2XL U1702 ( .B0(n2324), .B1(n2437), .A0N(\register[18][16] ), .A1N(
        n2439), .Y(n668) );
  OAI2BB2XL U1703 ( .B0(n2322), .B1(n2437), .A0N(\register[18][17] ), .A1N(
        n2438), .Y(n669) );
  OAI2BB2XL U1704 ( .B0(n2319), .B1(n2437), .A0N(\register[18][18] ), .A1N(
        n2438), .Y(n670) );
  OAI2BB2XL U1705 ( .B0(n2316), .B1(n2437), .A0N(\register[18][19] ), .A1N(
        n2438), .Y(n671) );
  OAI2BB2XL U1706 ( .B0(n2314), .B1(n2437), .A0N(\register[18][20] ), .A1N(
        n2438), .Y(n672) );
  OAI2BB2XL U1707 ( .B0(n2312), .B1(n2437), .A0N(\register[18][21] ), .A1N(
        n2438), .Y(n673) );
  OAI2BB2XL U1708 ( .B0(n2310), .B1(n2437), .A0N(\register[18][22] ), .A1N(
        n2439), .Y(n674) );
  OAI2BB2XL U1709 ( .B0(n2305), .B1(n2437), .A0N(\register[18][24] ), .A1N(
        n2439), .Y(n676) );
  OAI2BB2XL U1710 ( .B0(n2362), .B1(n2393), .A0N(\register[26][0] ), .A1N(
        n2391), .Y(n908) );
  OAI2BB2XL U1711 ( .B0(n2360), .B1(n2392), .A0N(\register[26][1] ), .A1N(
        n2391), .Y(n909) );
  OAI2BB2XL U1712 ( .B0(n2358), .B1(n2392), .A0N(\register[26][2] ), .A1N(
        n2391), .Y(n910) );
  OAI2BB2XL U1713 ( .B0(n2355), .B1(n2392), .A0N(\register[26][3] ), .A1N(
        n2395), .Y(n911) );
  OAI2BB2XL U1714 ( .B0(n2353), .B1(n2392), .A0N(\register[26][4] ), .A1N(
        n2391), .Y(n912) );
  OAI2BB2XL U1715 ( .B0(n2351), .B1(n2392), .A0N(\register[26][5] ), .A1N(
        n2395), .Y(n913) );
  OAI2BB2XL U1716 ( .B0(n2348), .B1(n2392), .A0N(\register[26][6] ), .A1N(
        n2395), .Y(n914) );
  OAI2BB2XL U1717 ( .B0(n2346), .B1(n2392), .A0N(\register[26][7] ), .A1N(
        n2395), .Y(n915) );
  OAI2BB2XL U1718 ( .B0(n2344), .B1(n2392), .A0N(\register[26][8] ), .A1N(
        n2395), .Y(n916) );
  OAI2BB2XL U1719 ( .B0(n2341), .B1(n2392), .A0N(\register[26][9] ), .A1N(
        n2395), .Y(n917) );
  OAI2BB2XL U1720 ( .B0(n2339), .B1(n2392), .A0N(\register[26][10] ), .A1N(
        n2395), .Y(n918) );
  OAI2BB2XL U1721 ( .B0(n2337), .B1(n2392), .A0N(\register[26][11] ), .A1N(
        n2395), .Y(n919) );
  OAI2BB2XL U1722 ( .B0(n2334), .B1(n2392), .A0N(\register[26][12] ), .A1N(
        n2395), .Y(n920) );
  OAI2BB2XL U1723 ( .B0(n2332), .B1(n2393), .A0N(\register[26][13] ), .A1N(
        n2395), .Y(n921) );
  OAI2BB2XL U1724 ( .B0(n2329), .B1(n2393), .A0N(\register[26][14] ), .A1N(
        n2395), .Y(n922) );
  OAI2BB2XL U1725 ( .B0(n2326), .B1(n2393), .A0N(\register[26][15] ), .A1N(
        n2394), .Y(n923) );
  OAI2BB2XL U1726 ( .B0(n2324), .B1(n2393), .A0N(\register[26][16] ), .A1N(
        n2395), .Y(n924) );
  OAI2BB2XL U1727 ( .B0(n2321), .B1(n2393), .A0N(\register[26][17] ), .A1N(
        n2394), .Y(n925) );
  OAI2BB2XL U1728 ( .B0(n2318), .B1(n2393), .A0N(\register[26][18] ), .A1N(
        n2394), .Y(n926) );
  OAI2BB2XL U1729 ( .B0(n2316), .B1(n2393), .A0N(\register[26][19] ), .A1N(
        n2394), .Y(n927) );
  OAI2BB2XL U1730 ( .B0(n2314), .B1(n2393), .A0N(\register[26][20] ), .A1N(
        n2394), .Y(n928) );
  OAI2BB2XL U1731 ( .B0(n2312), .B1(n2393), .A0N(\register[26][21] ), .A1N(
        n2394), .Y(n929) );
  OAI2BB2XL U1732 ( .B0(n2309), .B1(n2393), .A0N(\register[26][22] ), .A1N(
        n2395), .Y(n930) );
  OAI2BB2XL U1733 ( .B0(n2305), .B1(n2393), .A0N(\register[26][24] ), .A1N(
        n2395), .Y(n932) );
  OAI2BB2XL U1734 ( .B0(n2362), .B1(n2454), .A0N(\register[15][0] ), .A1N(
        n2451), .Y(n556) );
  OAI2BB2XL U1735 ( .B0(n2361), .B1(n2453), .A0N(\register[15][1] ), .A1N(
        n2451), .Y(n557) );
  OAI2BB2XL U1736 ( .B0(n2359), .B1(n2453), .A0N(\register[15][2] ), .A1N(
        n2451), .Y(n558) );
  OAI2BB2XL U1737 ( .B0(n2356), .B1(n2453), .A0N(\register[15][3] ), .A1N(
        n2456), .Y(n559) );
  OAI2BB2XL U1738 ( .B0(n2354), .B1(n2453), .A0N(\register[15][4] ), .A1N(
        n2451), .Y(n560) );
  OAI2BB2XL U1739 ( .B0(n2351), .B1(n2453), .A0N(\register[15][5] ), .A1N(
        n2456), .Y(n561) );
  OAI2BB2XL U1740 ( .B0(n2349), .B1(n2453), .A0N(\register[15][6] ), .A1N(
        n2456), .Y(n562) );
  OAI2BB2XL U1741 ( .B0(n2346), .B1(n2453), .A0N(\register[15][7] ), .A1N(
        n2456), .Y(n563) );
  OAI2BB2XL U1742 ( .B0(n2344), .B1(n2453), .A0N(\register[15][8] ), .A1N(
        n2456), .Y(n564) );
  OAI2BB2XL U1743 ( .B0(n2342), .B1(n2453), .A0N(\register[15][9] ), .A1N(
        n2456), .Y(n565) );
  OAI2BB2XL U1744 ( .B0(n2339), .B1(n2453), .A0N(\register[15][10] ), .A1N(
        n2456), .Y(n566) );
  OAI2BB2XL U1745 ( .B0(n2337), .B1(n2453), .A0N(\register[15][11] ), .A1N(
        n2456), .Y(n567) );
  OAI2BB2XL U1746 ( .B0(n2335), .B1(n2453), .A0N(\register[15][12] ), .A1N(
        n2456), .Y(n568) );
  OAI2BB2XL U1747 ( .B0(n2332), .B1(n2454), .A0N(\register[15][13] ), .A1N(
        n2456), .Y(n569) );
  OAI2BB2XL U1748 ( .B0(n2330), .B1(n2454), .A0N(\register[15][14] ), .A1N(
        n2456), .Y(n570) );
  OAI2BB2XL U1749 ( .B0(n2327), .B1(n2454), .A0N(\register[15][15] ), .A1N(
        n2455), .Y(n571) );
  OAI2BB2XL U1750 ( .B0(n2324), .B1(n2454), .A0N(\register[15][16] ), .A1N(
        n2456), .Y(n572) );
  OAI2BB2XL U1751 ( .B0(n2322), .B1(n2454), .A0N(\register[15][17] ), .A1N(
        n2455), .Y(n573) );
  OAI2BB2XL U1752 ( .B0(n2319), .B1(n2454), .A0N(\register[15][18] ), .A1N(
        n2455), .Y(n574) );
  OAI2BB2XL U1753 ( .B0(n2316), .B1(n2454), .A0N(\register[15][19] ), .A1N(
        n2455), .Y(n575) );
  OAI2BB2XL U1754 ( .B0(n2314), .B1(n2454), .A0N(\register[15][20] ), .A1N(
        n2455), .Y(n576) );
  OAI2BB2XL U1755 ( .B0(n2312), .B1(n2454), .A0N(\register[15][21] ), .A1N(
        n2455), .Y(n577) );
  OAI2BB2XL U1756 ( .B0(n2310), .B1(n2454), .A0N(\register[15][22] ), .A1N(
        n2456), .Y(n578) );
  OAI2BB2XL U1757 ( .B0(n2305), .B1(n2454), .A0N(\register[15][24] ), .A1N(
        n2456), .Y(n580) );
  OAI2BB2XL U1758 ( .B0(n2363), .B1(n2408), .A0N(\register[23][0] ), .A1N(
        n2411), .Y(n812) );
  OAI2BB2XL U1759 ( .B0(n2360), .B1(n2407), .A0N(\register[23][1] ), .A1N(
        n2411), .Y(n813) );
  OAI2BB2XL U1760 ( .B0(n2358), .B1(n2407), .A0N(\register[23][2] ), .A1N(
        n2411), .Y(n814) );
  OAI2BB2XL U1761 ( .B0(n2355), .B1(n2407), .A0N(\register[23][3] ), .A1N(
        n2410), .Y(n815) );
  OAI2BB2XL U1762 ( .B0(n2353), .B1(n2407), .A0N(\register[23][4] ), .A1N(
        n2411), .Y(n816) );
  OAI2BB2XL U1763 ( .B0(n2351), .B1(n2407), .A0N(\register[23][5] ), .A1N(
        n2410), .Y(n817) );
  OAI2BB2XL U1764 ( .B0(n2348), .B1(n2407), .A0N(\register[23][6] ), .A1N(
        n2410), .Y(n818) );
  OAI2BB2XL U1765 ( .B0(n2346), .B1(n2407), .A0N(\register[23][7] ), .A1N(
        n2410), .Y(n819) );
  OAI2BB2XL U1766 ( .B0(n2344), .B1(n2407), .A0N(\register[23][8] ), .A1N(
        n2410), .Y(n820) );
  OAI2BB2XL U1767 ( .B0(n2341), .B1(n2407), .A0N(\register[23][9] ), .A1N(
        n2410), .Y(n821) );
  OAI2BB2XL U1768 ( .B0(n2339), .B1(n2407), .A0N(\register[23][10] ), .A1N(
        n2410), .Y(n822) );
  OAI2BB2XL U1769 ( .B0(n2337), .B1(n2407), .A0N(\register[23][11] ), .A1N(
        n2410), .Y(n823) );
  OAI2BB2XL U1770 ( .B0(n2334), .B1(n2407), .A0N(\register[23][12] ), .A1N(
        n2410), .Y(n824) );
  OAI2BB2XL U1771 ( .B0(n2332), .B1(n2408), .A0N(\register[23][13] ), .A1N(
        n2410), .Y(n825) );
  OAI2BB2XL U1772 ( .B0(n2329), .B1(n2408), .A0N(\register[23][14] ), .A1N(
        n2410), .Y(n826) );
  OAI2BB2XL U1773 ( .B0(n2326), .B1(n2408), .A0N(\register[23][15] ), .A1N(
        n2409), .Y(n827) );
  OAI2BB2XL U1774 ( .B0(n2324), .B1(n2408), .A0N(\register[23][16] ), .A1N(
        n2410), .Y(n828) );
  OAI2BB2XL U1775 ( .B0(n2321), .B1(n2408), .A0N(\register[23][17] ), .A1N(
        n2409), .Y(n829) );
  OAI2BB2XL U1776 ( .B0(n2318), .B1(n2408), .A0N(\register[23][18] ), .A1N(
        n2409), .Y(n830) );
  OAI2BB2XL U1777 ( .B0(n2316), .B1(n2408), .A0N(\register[23][19] ), .A1N(
        n2409), .Y(n831) );
  OAI2BB2XL U1778 ( .B0(n2314), .B1(n2408), .A0N(\register[23][20] ), .A1N(
        n2409), .Y(n832) );
  OAI2BB2XL U1779 ( .B0(n2312), .B1(n2408), .A0N(\register[23][21] ), .A1N(
        n2409), .Y(n833) );
  OAI2BB2XL U1780 ( .B0(n2309), .B1(n2408), .A0N(\register[23][22] ), .A1N(
        n2410), .Y(n834) );
  OAI2BB2XL U1781 ( .B0(n2305), .B1(n2408), .A0N(\register[23][24] ), .A1N(
        n2410), .Y(n836) );
  OAI2BB2XL U1782 ( .B0(n2362), .B1(n2367), .A0N(\register[31][0] ), .A1N(
        n2364), .Y(n1068) );
  OAI2BB2XL U1783 ( .B0(n2360), .B1(n2366), .A0N(\register[31][1] ), .A1N(
        n2364), .Y(n1069) );
  OAI2BB2XL U1784 ( .B0(n2358), .B1(n2366), .A0N(\register[31][2] ), .A1N(
        n2364), .Y(n1070) );
  OAI2BB2XL U1785 ( .B0(n2355), .B1(n2366), .A0N(\register[31][3] ), .A1N(
        n2369), .Y(n1071) );
  OAI2BB2XL U1786 ( .B0(n2353), .B1(n2366), .A0N(\register[31][4] ), .A1N(
        n2364), .Y(n1072) );
  OAI2BB2XL U1787 ( .B0(n2351), .B1(n2366), .A0N(\register[31][5] ), .A1N(
        n2369), .Y(n1073) );
  OAI2BB2XL U1788 ( .B0(n2348), .B1(n2366), .A0N(\register[31][6] ), .A1N(
        n2369), .Y(n1074) );
  OAI2BB2XL U1789 ( .B0(n2346), .B1(n2366), .A0N(\register[31][7] ), .A1N(
        n2369), .Y(n1075) );
  OAI2BB2XL U1790 ( .B0(n2344), .B1(n2366), .A0N(\register[31][8] ), .A1N(
        n2369), .Y(n1076) );
  OAI2BB2XL U1791 ( .B0(n2341), .B1(n2366), .A0N(\register[31][9] ), .A1N(
        n2369), .Y(n1077) );
  OAI2BB2XL U1792 ( .B0(n2339), .B1(n2366), .A0N(\register[31][10] ), .A1N(
        n2369), .Y(n1078) );
  OAI2BB2XL U1793 ( .B0(n2337), .B1(n2366), .A0N(\register[31][11] ), .A1N(
        n2369), .Y(n1079) );
  OAI2BB2XL U1794 ( .B0(n2334), .B1(n2366), .A0N(\register[31][12] ), .A1N(
        n2369), .Y(n1080) );
  OAI2BB2XL U1795 ( .B0(n2332), .B1(n2367), .A0N(\register[31][13] ), .A1N(
        n2369), .Y(n1081) );
  OAI2BB2XL U1796 ( .B0(n2329), .B1(n2367), .A0N(\register[31][14] ), .A1N(
        n2369), .Y(n1082) );
  OAI2BB2XL U1797 ( .B0(n2326), .B1(n2367), .A0N(\register[31][15] ), .A1N(
        n2368), .Y(n1083) );
  OAI2BB2XL U1798 ( .B0(n2324), .B1(n2367), .A0N(\register[31][16] ), .A1N(
        n2369), .Y(n1084) );
  OAI2BB2XL U1799 ( .B0(n2321), .B1(n2367), .A0N(\register[31][17] ), .A1N(
        n2368), .Y(n1085) );
  OAI2BB2XL U1800 ( .B0(n2318), .B1(n2367), .A0N(\register[31][18] ), .A1N(
        n2368), .Y(n1086) );
  OAI2BB2XL U1801 ( .B0(n2316), .B1(n2367), .A0N(\register[31][19] ), .A1N(
        n2368), .Y(n1087) );
  OAI2BB2XL U1802 ( .B0(n2314), .B1(n2367), .A0N(\register[31][20] ), .A1N(
        n2368), .Y(n1088) );
  OAI2BB2XL U1803 ( .B0(n2312), .B1(n2367), .A0N(\register[31][21] ), .A1N(
        n2368), .Y(n1089) );
  OAI2BB2XL U1804 ( .B0(n2309), .B1(n2367), .A0N(\register[31][22] ), .A1N(
        n2369), .Y(n1090) );
  OAI2BB2XL U1805 ( .B0(n2305), .B1(n2367), .A0N(\register[31][24] ), .A1N(
        n2369), .Y(n1092) );
  OAI2BB2XL U1806 ( .B0(n2362), .B1(n2493), .A0N(\register[8][0] ), .A1N(n2492), .Y(n332) );
  OAI2BB2XL U1807 ( .B0(n2361), .B1(n2492), .A0N(\register[8][1] ), .A1N(n2493), .Y(n333) );
  OAI2BB2XL U1808 ( .B0(n2359), .B1(n2492), .A0N(\register[8][2] ), .A1N(n2492), .Y(n334) );
  OAI2BB2XL U1809 ( .B0(n2356), .B1(n2492), .A0N(\register[8][3] ), .A1N(n2495), .Y(n335) );
  OAI2BB2XL U1810 ( .B0(n2354), .B1(n2492), .A0N(\register[8][4] ), .A1N(n2493), .Y(n336) );
  OAI2BB2XL U1811 ( .B0(n2351), .B1(n2492), .A0N(\register[8][5] ), .A1N(n2495), .Y(n337) );
  OAI2BB2XL U1812 ( .B0(n2349), .B1(n2492), .A0N(\register[8][6] ), .A1N(n2495), .Y(n338) );
  OAI2BB2XL U1813 ( .B0(n2346), .B1(n2492), .A0N(\register[8][7] ), .A1N(n2495), .Y(n339) );
  OAI2BB2XL U1814 ( .B0(n2344), .B1(n2492), .A0N(\register[8][8] ), .A1N(n2495), .Y(n340) );
  OAI2BB2XL U1815 ( .B0(n2342), .B1(n2492), .A0N(\register[8][9] ), .A1N(n2495), .Y(n341) );
  OAI2BB2XL U1816 ( .B0(n2339), .B1(n2492), .A0N(\register[8][10] ), .A1N(
        n2495), .Y(n342) );
  OAI2BB2XL U1817 ( .B0(n2337), .B1(n2492), .A0N(\register[8][11] ), .A1N(
        n2495), .Y(n343) );
  OAI2BB2XL U1818 ( .B0(n2335), .B1(n2492), .A0N(\register[8][12] ), .A1N(
        n2495), .Y(n344) );
  OAI2BB2XL U1819 ( .B0(n2332), .B1(n2493), .A0N(\register[8][13] ), .A1N(
        n2495), .Y(n345) );
  OAI2BB2XL U1820 ( .B0(n2330), .B1(n2493), .A0N(\register[8][14] ), .A1N(
        n2495), .Y(n346) );
  OAI2BB2XL U1821 ( .B0(n2327), .B1(n2493), .A0N(\register[8][15] ), .A1N(
        n2494), .Y(n347) );
  OAI2BB2XL U1822 ( .B0(n2324), .B1(n2493), .A0N(\register[8][16] ), .A1N(
        n2495), .Y(n348) );
  OAI2BB2XL U1823 ( .B0(n2322), .B1(n2493), .A0N(\register[8][17] ), .A1N(
        n2494), .Y(n349) );
  OAI2BB2XL U1824 ( .B0(n2319), .B1(n2493), .A0N(\register[8][18] ), .A1N(
        n2494), .Y(n350) );
  OAI2BB2XL U1825 ( .B0(n2316), .B1(n2493), .A0N(\register[8][19] ), .A1N(
        n2494), .Y(n351) );
  OAI2BB2XL U1826 ( .B0(n2314), .B1(n2493), .A0N(\register[8][20] ), .A1N(
        n2494), .Y(n352) );
  OAI2BB2XL U1827 ( .B0(n2312), .B1(n2493), .A0N(\register[8][21] ), .A1N(
        n2494), .Y(n353) );
  OAI2BB2XL U1828 ( .B0(n2310), .B1(n2493), .A0N(\register[8][22] ), .A1N(
        n2495), .Y(n354) );
  OAI2BB2XL U1829 ( .B0(n2305), .B1(n2493), .A0N(\register[8][24] ), .A1N(
        n2495), .Y(n356) );
  OAI2BB2XL U1830 ( .B0(n2362), .B1(n2448), .A0N(\register[16][0] ), .A1N(
        n2446), .Y(n588) );
  OAI2BB2XL U1831 ( .B0(n2361), .B1(n2447), .A0N(\register[16][1] ), .A1N(
        n2446), .Y(n589) );
  OAI2BB2XL U1832 ( .B0(n2359), .B1(n2447), .A0N(\register[16][2] ), .A1N(
        n2446), .Y(n590) );
  OAI2BB2XL U1833 ( .B0(n2356), .B1(n2447), .A0N(\register[16][3] ), .A1N(
        n2450), .Y(n591) );
  OAI2BB2XL U1834 ( .B0(n2354), .B1(n2447), .A0N(\register[16][4] ), .A1N(
        n2446), .Y(n592) );
  OAI2BB2XL U1835 ( .B0(n2351), .B1(n2447), .A0N(\register[16][5] ), .A1N(
        n2450), .Y(n593) );
  OAI2BB2XL U1836 ( .B0(n2349), .B1(n2447), .A0N(\register[16][6] ), .A1N(
        n2450), .Y(n594) );
  OAI2BB2XL U1837 ( .B0(n2346), .B1(n2447), .A0N(\register[16][7] ), .A1N(
        n2450), .Y(n595) );
  OAI2BB2XL U1838 ( .B0(n2344), .B1(n2447), .A0N(\register[16][8] ), .A1N(
        n2450), .Y(n596) );
  OAI2BB2XL U1839 ( .B0(n2342), .B1(n2447), .A0N(\register[16][9] ), .A1N(
        n2450), .Y(n597) );
  OAI2BB2XL U1840 ( .B0(n2339), .B1(n2447), .A0N(\register[16][10] ), .A1N(
        n2450), .Y(n598) );
  OAI2BB2XL U1841 ( .B0(n2337), .B1(n2447), .A0N(\register[16][11] ), .A1N(
        n2450), .Y(n599) );
  OAI2BB2XL U1842 ( .B0(n2335), .B1(n2447), .A0N(\register[16][12] ), .A1N(
        n2450), .Y(n600) );
  OAI2BB2XL U1843 ( .B0(n2332), .B1(n2448), .A0N(\register[16][13] ), .A1N(
        n2450), .Y(n601) );
  OAI2BB2XL U1844 ( .B0(n2330), .B1(n2448), .A0N(\register[16][14] ), .A1N(
        n2450), .Y(n602) );
  OAI2BB2XL U1845 ( .B0(n2327), .B1(n2448), .A0N(\register[16][15] ), .A1N(
        n2449), .Y(n603) );
  OAI2BB2XL U1846 ( .B0(n2324), .B1(n2448), .A0N(\register[16][16] ), .A1N(
        n2450), .Y(n604) );
  OAI2BB2XL U1847 ( .B0(n2322), .B1(n2448), .A0N(\register[16][17] ), .A1N(
        n2449), .Y(n605) );
  OAI2BB2XL U1848 ( .B0(n2319), .B1(n2448), .A0N(\register[16][18] ), .A1N(
        n2449), .Y(n606) );
  OAI2BB2XL U1849 ( .B0(n2316), .B1(n2448), .A0N(\register[16][19] ), .A1N(
        n2449), .Y(n607) );
  OAI2BB2XL U1850 ( .B0(n2314), .B1(n2448), .A0N(\register[16][20] ), .A1N(
        n2449), .Y(n608) );
  OAI2BB2XL U1851 ( .B0(n2312), .B1(n2448), .A0N(\register[16][21] ), .A1N(
        n2449), .Y(n609) );
  OAI2BB2XL U1852 ( .B0(n2310), .B1(n2448), .A0N(\register[16][22] ), .A1N(
        n2450), .Y(n610) );
  OAI2BB2XL U1853 ( .B0(n2305), .B1(n2448), .A0N(\register[16][24] ), .A1N(
        n2450), .Y(n612) );
  OAI2BB2XL U1854 ( .B0(n2363), .B1(n2403), .A0N(\register[24][0] ), .A1N(
        n2402), .Y(n844) );
  OAI2BB2XL U1855 ( .B0(n2360), .B1(n2402), .A0N(\register[24][1] ), .A1N(
        n2403), .Y(n845) );
  OAI2BB2XL U1856 ( .B0(n2358), .B1(n2402), .A0N(\register[24][2] ), .A1N(
        n2403), .Y(n846) );
  OAI2BB2XL U1857 ( .B0(n2355), .B1(n2402), .A0N(\register[24][3] ), .A1N(
        n2405), .Y(n847) );
  OAI2BB2XL U1858 ( .B0(n2353), .B1(n2402), .A0N(\register[24][4] ), .A1N(
        n2402), .Y(n848) );
  OAI2BB2XL U1859 ( .B0(n2352), .B1(n2402), .A0N(\register[24][5] ), .A1N(
        n2405), .Y(n849) );
  OAI2BB2XL U1860 ( .B0(n2348), .B1(n2402), .A0N(\register[24][6] ), .A1N(
        n2405), .Y(n850) );
  OAI2BB2XL U1861 ( .B0(n2347), .B1(n2402), .A0N(\register[24][7] ), .A1N(
        n2405), .Y(n851) );
  OAI2BB2XL U1862 ( .B0(n2345), .B1(n2402), .A0N(\register[24][8] ), .A1N(
        n2405), .Y(n852) );
  OAI2BB2XL U1863 ( .B0(n2341), .B1(n2402), .A0N(\register[24][9] ), .A1N(
        n2405), .Y(n853) );
  OAI2BB2XL U1864 ( .B0(n2340), .B1(n2402), .A0N(\register[24][10] ), .A1N(
        n2405), .Y(n854) );
  OAI2BB2XL U1865 ( .B0(n2338), .B1(n2402), .A0N(\register[24][11] ), .A1N(
        n2405), .Y(n855) );
  OAI2BB2XL U1866 ( .B0(n2334), .B1(n2402), .A0N(\register[24][12] ), .A1N(
        n2405), .Y(n856) );
  OAI2BB2XL U1867 ( .B0(n2333), .B1(n2403), .A0N(\register[24][13] ), .A1N(
        n2405), .Y(n857) );
  OAI2BB2XL U1868 ( .B0(n2329), .B1(n2403), .A0N(\register[24][14] ), .A1N(
        n2405), .Y(n858) );
  OAI2BB2XL U1869 ( .B0(n2326), .B1(n2403), .A0N(\register[24][15] ), .A1N(
        n2404), .Y(n859) );
  OAI2BB2XL U1870 ( .B0(n2325), .B1(n2403), .A0N(\register[24][16] ), .A1N(
        n2405), .Y(n860) );
  OAI2BB2XL U1871 ( .B0(n2321), .B1(n2403), .A0N(\register[24][17] ), .A1N(
        n2404), .Y(n861) );
  OAI2BB2XL U1872 ( .B0(n2318), .B1(n2403), .A0N(\register[24][18] ), .A1N(
        n2404), .Y(n862) );
  OAI2BB2XL U1873 ( .B0(n2317), .B1(n2403), .A0N(\register[24][19] ), .A1N(
        n2404), .Y(n863) );
  OAI2BB2XL U1874 ( .B0(n2315), .B1(n2403), .A0N(\register[24][20] ), .A1N(
        n2404), .Y(n864) );
  OAI2BB2XL U1875 ( .B0(n2313), .B1(n2403), .A0N(\register[24][21] ), .A1N(
        n2404), .Y(n865) );
  OAI2BB2XL U1876 ( .B0(n2309), .B1(n2403), .A0N(\register[24][22] ), .A1N(
        n2405), .Y(n866) );
  OAI2BB2XL U1877 ( .B0(n2306), .B1(n2403), .A0N(\register[24][24] ), .A1N(
        n2405), .Y(n868) );
  OAI2BB2XL U1878 ( .B0(n2327), .B1(n2466), .A0N(\register[13][15] ), .A1N(
        n2467), .Y(n507) );
  OAI2BB2XL U1879 ( .B0(n2322), .B1(n2466), .A0N(\register[13][17] ), .A1N(
        n2467), .Y(n509) );
  OAI2BB2XL U1880 ( .B0(n2319), .B1(n2466), .A0N(\register[13][18] ), .A1N(
        n2467), .Y(n510) );
  OAI2BB2XL U1881 ( .B0(n2316), .B1(n2466), .A0N(\register[13][19] ), .A1N(
        n2467), .Y(n511) );
  OAI2BB2XL U1882 ( .B0(n2314), .B1(n2466), .A0N(\register[13][20] ), .A1N(
        n2467), .Y(n512) );
  OAI2BB2XL U1883 ( .B0(n2312), .B1(n2466), .A0N(\register[13][21] ), .A1N(
        n2467), .Y(n513) );
  OAI2BB2XL U1884 ( .B0(n2326), .B1(n2420), .A0N(\register[21][15] ), .A1N(
        n2421), .Y(n763) );
  OAI2BB2XL U1885 ( .B0(n2321), .B1(n2420), .A0N(\register[21][17] ), .A1N(
        n2421), .Y(n765) );
  OAI2BB2XL U1886 ( .B0(n2318), .B1(n2420), .A0N(\register[21][18] ), .A1N(
        n2421), .Y(n766) );
  OAI2BB2XL U1887 ( .B0(n2317), .B1(n2420), .A0N(\register[21][19] ), .A1N(
        n2421), .Y(n767) );
  OAI2BB2XL U1888 ( .B0(n2315), .B1(n2420), .A0N(\register[21][20] ), .A1N(
        n2421), .Y(n768) );
  OAI2BB2XL U1889 ( .B0(n2313), .B1(n2420), .A0N(\register[21][21] ), .A1N(
        n2421), .Y(n769) );
  OAI2BB2XL U1890 ( .B0(n2326), .B1(n2378), .A0N(\register[29][15] ), .A1N(
        n2379), .Y(n1019) );
  OAI2BB2XL U1891 ( .B0(n2321), .B1(n2378), .A0N(\register[29][17] ), .A1N(
        n2379), .Y(n1021) );
  OAI2BB2XL U1892 ( .B0(n2318), .B1(n2378), .A0N(\register[29][18] ), .A1N(
        n2379), .Y(n1022) );
  OAI2BB2XL U1893 ( .B0(n2317), .B1(n2378), .A0N(\register[29][19] ), .A1N(
        n2379), .Y(n1023) );
  OAI2BB2XL U1894 ( .B0(n2315), .B1(n2378), .A0N(\register[29][20] ), .A1N(
        n2379), .Y(n1024) );
  OAI2BB2XL U1895 ( .B0(n2313), .B1(n2378), .A0N(\register[29][21] ), .A1N(
        n2379), .Y(n1025) );
  OAI2BB2XL U1896 ( .B0(n2356), .B1(n2465), .A0N(\register[13][3] ), .A1N(
        n2468), .Y(n495) );
  OAI2BB2XL U1897 ( .B0(n2351), .B1(n2465), .A0N(\register[13][5] ), .A1N(
        n2468), .Y(n497) );
  OAI2BB2XL U1898 ( .B0(n2349), .B1(n2465), .A0N(\register[13][6] ), .A1N(
        n2468), .Y(n498) );
  OAI2BB2XL U1899 ( .B0(n2346), .B1(n2465), .A0N(\register[13][7] ), .A1N(
        n2468), .Y(n499) );
  OAI2BB2XL U1900 ( .B0(n2344), .B1(n2465), .A0N(\register[13][8] ), .A1N(
        n2468), .Y(n500) );
  OAI2BB2XL U1901 ( .B0(n2342), .B1(n2465), .A0N(\register[13][9] ), .A1N(
        n2468), .Y(n501) );
  OAI2BB2XL U1902 ( .B0(n2339), .B1(n2465), .A0N(\register[13][10] ), .A1N(
        n2468), .Y(n502) );
  OAI2BB2XL U1903 ( .B0(n2337), .B1(n2465), .A0N(\register[13][11] ), .A1N(
        n2468), .Y(n503) );
  OAI2BB2XL U1904 ( .B0(n2335), .B1(n2465), .A0N(\register[13][12] ), .A1N(
        n2468), .Y(n504) );
  OAI2BB2XL U1905 ( .B0(n2332), .B1(n2466), .A0N(\register[13][13] ), .A1N(
        n2468), .Y(n505) );
  OAI2BB2XL U1906 ( .B0(n2330), .B1(n2466), .A0N(\register[13][14] ), .A1N(
        n2468), .Y(n506) );
  OAI2BB2XL U1907 ( .B0(n2324), .B1(n2466), .A0N(\register[13][16] ), .A1N(
        n2468), .Y(n508) );
  OAI2BB2XL U1908 ( .B0(n2310), .B1(n2466), .A0N(\register[13][22] ), .A1N(
        n2468), .Y(n514) );
  OAI2BB2XL U1909 ( .B0(n2305), .B1(n2466), .A0N(\register[13][24] ), .A1N(
        n2468), .Y(n516) );
  OAI2BB2XL U1910 ( .B0(n2355), .B1(n2419), .A0N(\register[21][3] ), .A1N(
        n2422), .Y(n751) );
  OAI2BB2XL U1911 ( .B0(n2352), .B1(n2419), .A0N(\register[21][5] ), .A1N(
        n2422), .Y(n753) );
  OAI2BB2XL U1912 ( .B0(n2348), .B1(n2419), .A0N(\register[21][6] ), .A1N(
        n2422), .Y(n754) );
  OAI2BB2XL U1913 ( .B0(n2347), .B1(n2419), .A0N(\register[21][7] ), .A1N(
        n2422), .Y(n755) );
  OAI2BB2XL U1914 ( .B0(n2345), .B1(n2419), .A0N(\register[21][8] ), .A1N(
        n2422), .Y(n756) );
  OAI2BB2XL U1915 ( .B0(n2341), .B1(n2419), .A0N(\register[21][9] ), .A1N(
        n2422), .Y(n757) );
  OAI2BB2XL U1916 ( .B0(n2340), .B1(n2419), .A0N(\register[21][10] ), .A1N(
        n2422), .Y(n758) );
  OAI2BB2XL U1917 ( .B0(n2338), .B1(n2419), .A0N(\register[21][11] ), .A1N(
        n2422), .Y(n759) );
  OAI2BB2XL U1918 ( .B0(n2334), .B1(n2419), .A0N(\register[21][12] ), .A1N(
        n2422), .Y(n760) );
  OAI2BB2XL U1919 ( .B0(n2333), .B1(n2420), .A0N(\register[21][13] ), .A1N(
        n2422), .Y(n761) );
  OAI2BB2XL U1920 ( .B0(n2329), .B1(n2420), .A0N(\register[21][14] ), .A1N(
        n2422), .Y(n762) );
  OAI2BB2XL U1921 ( .B0(n2325), .B1(n2420), .A0N(\register[21][16] ), .A1N(
        n2422), .Y(n764) );
  OAI2BB2XL U1922 ( .B0(n2309), .B1(n2420), .A0N(\register[21][22] ), .A1N(
        n2422), .Y(n770) );
  OAI2BB2XL U1923 ( .B0(n2306), .B1(n2420), .A0N(\register[21][24] ), .A1N(
        n2422), .Y(n772) );
  OAI2BB2XL U1924 ( .B0(n2355), .B1(n2377), .A0N(\register[29][3] ), .A1N(
        n2380), .Y(n1007) );
  OAI2BB2XL U1925 ( .B0(n2352), .B1(n2377), .A0N(\register[29][5] ), .A1N(
        n2380), .Y(n1009) );
  OAI2BB2XL U1926 ( .B0(n2348), .B1(n2377), .A0N(\register[29][6] ), .A1N(
        n2380), .Y(n1010) );
  OAI2BB2XL U1927 ( .B0(n2347), .B1(n2377), .A0N(\register[29][7] ), .A1N(
        n2380), .Y(n1011) );
  OAI2BB2XL U1928 ( .B0(n2345), .B1(n2377), .A0N(\register[29][8] ), .A1N(
        n2380), .Y(n1012) );
  OAI2BB2XL U1929 ( .B0(n2341), .B1(n2377), .A0N(\register[29][9] ), .A1N(
        n2380), .Y(n1013) );
  OAI2BB2XL U1930 ( .B0(n2340), .B1(n2377), .A0N(\register[29][10] ), .A1N(
        n2380), .Y(n1014) );
  OAI2BB2XL U1931 ( .B0(n2338), .B1(n2377), .A0N(\register[29][11] ), .A1N(
        n2380), .Y(n1015) );
  OAI2BB2XL U1932 ( .B0(n2334), .B1(n2377), .A0N(\register[29][12] ), .A1N(
        n2380), .Y(n1016) );
  OAI2BB2XL U1933 ( .B0(n2333), .B1(n2378), .A0N(\register[29][13] ), .A1N(
        n2380), .Y(n1017) );
  OAI2BB2XL U1934 ( .B0(n2329), .B1(n2378), .A0N(\register[29][14] ), .A1N(
        n2380), .Y(n1018) );
  OAI2BB2XL U1935 ( .B0(n2325), .B1(n2378), .A0N(\register[29][16] ), .A1N(
        n2380), .Y(n1020) );
  OAI2BB2XL U1936 ( .B0(n2309), .B1(n2378), .A0N(\register[29][22] ), .A1N(
        n2380), .Y(n1026) );
  OAI2BB2XL U1937 ( .B0(n2306), .B1(n2378), .A0N(\register[29][24] ), .A1N(
        n2380), .Y(n1028) );
  OAI2BB2XL U1938 ( .B0(n2362), .B1(n2466), .A0N(\register[13][0] ), .A1N(
        n2463), .Y(n492) );
  OAI2BB2XL U1939 ( .B0(n2361), .B1(n2465), .A0N(\register[13][1] ), .A1N(
        n2463), .Y(n493) );
  OAI2BB2XL U1940 ( .B0(n2359), .B1(n2465), .A0N(\register[13][2] ), .A1N(
        n2463), .Y(n494) );
  OAI2BB2XL U1941 ( .B0(n2354), .B1(n2465), .A0N(\register[13][4] ), .A1N(
        n2463), .Y(n496) );
  OAI2BB2XL U1942 ( .B0(n2363), .B1(n2420), .A0N(\register[21][0] ), .A1N(
        n2423), .Y(n748) );
  OAI2BB2XL U1943 ( .B0(n2360), .B1(n2419), .A0N(\register[21][1] ), .A1N(
        n2423), .Y(n749) );
  OAI2BB2XL U1944 ( .B0(n2358), .B1(n2419), .A0N(\register[21][2] ), .A1N(
        n2423), .Y(n750) );
  OAI2BB2XL U1945 ( .B0(n2353), .B1(n2419), .A0N(\register[21][4] ), .A1N(
        n2423), .Y(n752) );
  OAI2BB2XL U1946 ( .B0(n2362), .B1(n2378), .A0N(\register[29][0] ), .A1N(
        n2376), .Y(n1004) );
  OAI2BB2XL U1947 ( .B0(n2360), .B1(n2377), .A0N(\register[29][1] ), .A1N(
        n2376), .Y(n1005) );
  OAI2BB2XL U1948 ( .B0(n2358), .B1(n2377), .A0N(\register[29][2] ), .A1N(
        n2376), .Y(n1006) );
  OAI2BB2XL U1949 ( .B0(n2353), .B1(n2377), .A0N(\register[29][4] ), .A1N(
        n2376), .Y(n1008) );
  OAI2BB2XL U1950 ( .B0(n2363), .B1(n2514), .A0N(\register[4][0] ), .A1N(n2513), .Y(n204) );
  OAI2BB2XL U1951 ( .B0(n2361), .B1(n2513), .A0N(\register[4][1] ), .A1N(n2513), .Y(n205) );
  OAI2BB2XL U1952 ( .B0(n2612), .B1(n2513), .A0N(\register[4][2] ), .A1N(n2513), .Y(n206) );
  OAI2BB2XL U1953 ( .B0(n2357), .B1(n2513), .A0N(\register[4][3] ), .A1N(n2516), .Y(n207) );
  OAI2BB2XL U1954 ( .B0(n2610), .B1(n2513), .A0N(\register[4][4] ), .A1N(n2513), .Y(n208) );
  OAI2BB2XL U1955 ( .B0(n2352), .B1(n2513), .A0N(\register[4][5] ), .A1N(n2516), .Y(n209) );
  OAI2BB2XL U1956 ( .B0(n2350), .B1(n2513), .A0N(\register[4][6] ), .A1N(n2516), .Y(n210) );
  OAI2BB2XL U1957 ( .B0(n2347), .B1(n2513), .A0N(\register[4][7] ), .A1N(n2516), .Y(n211) );
  OAI2BB2XL U1958 ( .B0(n2345), .B1(n2513), .A0N(\register[4][8] ), .A1N(n2516), .Y(n212) );
  OAI2BB2XL U1959 ( .B0(n2343), .B1(n2514), .A0N(\register[4][9] ), .A1N(n2516), .Y(n213) );
  OAI2BB2XL U1960 ( .B0(n2340), .B1(n2514), .A0N(\register[4][10] ), .A1N(
        n2516), .Y(n214) );
  OAI2BB2XL U1961 ( .B0(n2338), .B1(n2514), .A0N(\register[4][11] ), .A1N(
        n2516), .Y(n215) );
  OAI2BB2XL U1962 ( .B0(n2336), .B1(n2514), .A0N(\register[4][12] ), .A1N(
        n2516), .Y(n216) );
  OAI2BB2XL U1963 ( .B0(n2333), .B1(n2514), .A0N(\register[4][13] ), .A1N(
        n2516), .Y(n217) );
  OAI2BB2XL U1964 ( .B0(n2331), .B1(n2514), .A0N(\register[4][14] ), .A1N(
        n2516), .Y(n218) );
  OAI2BB2XL U1965 ( .B0(n2328), .B1(n2514), .A0N(\register[4][15] ), .A1N(
        n2515), .Y(n219) );
  OAI2BB2XL U1966 ( .B0(n2325), .B1(n2514), .A0N(\register[4][16] ), .A1N(
        n2516), .Y(n220) );
  OAI2BB2XL U1967 ( .B0(n2323), .B1(n2514), .A0N(\register[4][17] ), .A1N(
        n2515), .Y(n221) );
  OAI2BB2XL U1968 ( .B0(n2320), .B1(n2514), .A0N(\register[4][18] ), .A1N(
        n2515), .Y(n222) );
  OAI2BB2XL U1969 ( .B0(n2317), .B1(n2514), .A0N(\register[4][19] ), .A1N(
        n2515), .Y(n223) );
  OAI2BB2XL U1970 ( .B0(n2315), .B1(n2514), .A0N(\register[4][20] ), .A1N(
        n2515), .Y(n224) );
  OAI2BB2XL U1971 ( .B0(n2313), .B1(n2514), .A0N(\register[4][21] ), .A1N(
        n2515), .Y(n225) );
  OAI2BB2XL U1972 ( .B0(n2311), .B1(n2514), .A0N(\register[4][22] ), .A1N(
        n2516), .Y(n226) );
  OAI2BB2XL U1973 ( .B0(n2306), .B1(n2514), .A0N(\register[4][24] ), .A1N(
        n2516), .Y(n228) );
  OAI2BB2XL U1974 ( .B0(n2363), .B1(n2505), .A0N(\register[6][0] ), .A1N(n2503), .Y(n268) );
  OAI2BB2XL U1975 ( .B0(n2360), .B1(n2504), .A0N(\register[6][1] ), .A1N(n2503), .Y(n269) );
  OAI2BB2XL U1976 ( .B0(n2612), .B1(n2504), .A0N(\register[6][2] ), .A1N(n2503), .Y(n270) );
  OAI2BB2XL U1977 ( .B0(n2357), .B1(n2504), .A0N(\register[6][3] ), .A1N(n2507), .Y(n271) );
  OAI2BB2XL U1978 ( .B0(n2610), .B1(n2504), .A0N(\register[6][4] ), .A1N(n2503), .Y(n272) );
  OAI2BB2XL U1979 ( .B0(n2352), .B1(n2504), .A0N(\register[6][5] ), .A1N(n2507), .Y(n273) );
  OAI2BB2XL U1980 ( .B0(n2350), .B1(n2504), .A0N(\register[6][6] ), .A1N(n2507), .Y(n274) );
  OAI2BB2XL U1981 ( .B0(n2347), .B1(n2504), .A0N(\register[6][7] ), .A1N(n2507), .Y(n275) );
  OAI2BB2XL U1982 ( .B0(n2345), .B1(n2504), .A0N(\register[6][8] ), .A1N(n2507), .Y(n276) );
  OAI2BB2XL U1983 ( .B0(n2343), .B1(n2504), .A0N(\register[6][9] ), .A1N(n2507), .Y(n277) );
  OAI2BB2XL U1984 ( .B0(n2340), .B1(n2504), .A0N(\register[6][10] ), .A1N(
        n2507), .Y(n278) );
  OAI2BB2XL U1985 ( .B0(n2338), .B1(n2504), .A0N(\register[6][11] ), .A1N(
        n2507), .Y(n279) );
  OAI2BB2XL U1986 ( .B0(n2336), .B1(n2504), .A0N(\register[6][12] ), .A1N(
        n2507), .Y(n280) );
  OAI2BB2XL U1987 ( .B0(n2333), .B1(n2505), .A0N(\register[6][13] ), .A1N(
        n2507), .Y(n281) );
  OAI2BB2XL U1988 ( .B0(n2331), .B1(n2505), .A0N(\register[6][14] ), .A1N(
        n2507), .Y(n282) );
  OAI2BB2XL U1989 ( .B0(n2328), .B1(n2505), .A0N(\register[6][15] ), .A1N(
        n2506), .Y(n283) );
  OAI2BB2XL U1990 ( .B0(n2325), .B1(n2505), .A0N(\register[6][16] ), .A1N(
        n2507), .Y(n284) );
  OAI2BB2XL U1991 ( .B0(n2323), .B1(n2505), .A0N(\register[6][17] ), .A1N(
        n2506), .Y(n285) );
  OAI2BB2XL U1992 ( .B0(n2320), .B1(n2505), .A0N(\register[6][18] ), .A1N(
        n2506), .Y(n286) );
  OAI2BB2XL U1993 ( .B0(n2317), .B1(n2505), .A0N(\register[6][19] ), .A1N(
        n2506), .Y(n287) );
  OAI2BB2XL U1994 ( .B0(n2315), .B1(n2505), .A0N(\register[6][20] ), .A1N(
        n2506), .Y(n288) );
  OAI2BB2XL U1995 ( .B0(n2313), .B1(n2505), .A0N(\register[6][21] ), .A1N(
        n2506), .Y(n289) );
  OAI2BB2XL U1996 ( .B0(n2311), .B1(n2505), .A0N(\register[6][22] ), .A1N(
        n2507), .Y(n290) );
  OAI2BB2XL U1997 ( .B0(n2306), .B1(n2505), .A0N(\register[6][24] ), .A1N(
        n2507), .Y(n292) );
  OAI2BB2XL U1998 ( .B0(n2363), .B1(n2524), .A0N(\register[2][0] ), .A1N(n2522), .Y(n140) );
  OAI2BB2XL U1999 ( .B0(n2613), .B1(n2523), .A0N(\register[2][1] ), .A1N(n2522), .Y(n141) );
  OAI2BB2XL U2000 ( .B0(n2612), .B1(n2523), .A0N(\register[2][2] ), .A1N(n2522), .Y(n142) );
  OAI2BB2XL U2001 ( .B0(n2357), .B1(n2523), .A0N(\register[2][3] ), .A1N(n2526), .Y(n143) );
  OAI2BB2XL U2002 ( .B0(n2610), .B1(n2523), .A0N(\register[2][4] ), .A1N(n2522), .Y(n144) );
  OAI2BB2XL U2003 ( .B0(n2352), .B1(n2523), .A0N(\register[2][5] ), .A1N(n2526), .Y(n145) );
  OAI2BB2XL U2004 ( .B0(n2350), .B1(n2523), .A0N(\register[2][6] ), .A1N(n2526), .Y(n146) );
  OAI2BB2XL U2005 ( .B0(n2347), .B1(n2523), .A0N(\register[2][7] ), .A1N(n2526), .Y(n147) );
  OAI2BB2XL U2006 ( .B0(n2345), .B1(n2523), .A0N(\register[2][8] ), .A1N(n2526), .Y(n148) );
  OAI2BB2XL U2007 ( .B0(n2343), .B1(n2523), .A0N(\register[2][9] ), .A1N(n2526), .Y(n149) );
  OAI2BB2XL U2008 ( .B0(n2340), .B1(n2523), .A0N(\register[2][10] ), .A1N(
        n2526), .Y(n150) );
  OAI2BB2XL U2009 ( .B0(n2338), .B1(n2523), .A0N(\register[2][11] ), .A1N(
        n2526), .Y(n151) );
  OAI2BB2XL U2010 ( .B0(n2336), .B1(n2523), .A0N(\register[2][12] ), .A1N(
        n2526), .Y(n152) );
  OAI2BB2XL U2011 ( .B0(n2333), .B1(n2524), .A0N(\register[2][13] ), .A1N(
        n2526), .Y(n153) );
  OAI2BB2XL U2012 ( .B0(n2331), .B1(n2524), .A0N(\register[2][14] ), .A1N(
        n2526), .Y(n154) );
  OAI2BB2XL U2013 ( .B0(n2328), .B1(n2524), .A0N(\register[2][15] ), .A1N(
        n2525), .Y(n155) );
  OAI2BB2XL U2014 ( .B0(n2325), .B1(n2524), .A0N(\register[2][16] ), .A1N(
        n2526), .Y(n156) );
  OAI2BB2XL U2015 ( .B0(n2323), .B1(n2524), .A0N(\register[2][17] ), .A1N(
        n2525), .Y(n157) );
  OAI2BB2XL U2016 ( .B0(n2320), .B1(n2524), .A0N(\register[2][18] ), .A1N(
        n2525), .Y(n158) );
  OAI2BB2XL U2017 ( .B0(n2317), .B1(n2524), .A0N(\register[2][19] ), .A1N(
        n2525), .Y(n159) );
  OAI2BB2XL U2018 ( .B0(n2315), .B1(n2524), .A0N(\register[2][20] ), .A1N(
        n2525), .Y(n160) );
  OAI2BB2XL U2019 ( .B0(n2313), .B1(n2524), .A0N(\register[2][21] ), .A1N(
        n2525), .Y(n161) );
  OAI2BB2XL U2020 ( .B0(n2311), .B1(n2524), .A0N(\register[2][22] ), .A1N(
        n2526), .Y(n162) );
  OAI2BB2XL U2021 ( .B0(n2306), .B1(n2524), .A0N(\register[2][24] ), .A1N(
        n2526), .Y(n164) );
  OAI2BB2XL U2022 ( .B0(n2363), .B1(n2499), .A0N(\register[7][0] ), .A1N(n2496), .Y(n300) );
  OAI2BB2XL U2023 ( .B0(n2361), .B1(n2498), .A0N(\register[7][1] ), .A1N(n2496), .Y(n301) );
  OAI2BB2XL U2024 ( .B0(n2612), .B1(n2498), .A0N(\register[7][2] ), .A1N(n2496), .Y(n302) );
  OAI2BB2XL U2025 ( .B0(n2357), .B1(n2498), .A0N(\register[7][3] ), .A1N(n2501), .Y(n303) );
  OAI2BB2XL U2026 ( .B0(n2610), .B1(n2498), .A0N(\register[7][4] ), .A1N(n2496), .Y(n304) );
  OAI2BB2XL U2027 ( .B0(n2352), .B1(n2498), .A0N(\register[7][5] ), .A1N(n2501), .Y(n305) );
  OAI2BB2XL U2028 ( .B0(n2350), .B1(n2498), .A0N(\register[7][6] ), .A1N(n2501), .Y(n306) );
  OAI2BB2XL U2029 ( .B0(n2347), .B1(n2498), .A0N(\register[7][7] ), .A1N(n2501), .Y(n307) );
  OAI2BB2XL U2030 ( .B0(n2345), .B1(n2498), .A0N(\register[7][8] ), .A1N(n2501), .Y(n308) );
  OAI2BB2XL U2031 ( .B0(n2343), .B1(n2498), .A0N(\register[7][9] ), .A1N(n2501), .Y(n309) );
  OAI2BB2XL U2032 ( .B0(n2340), .B1(n2498), .A0N(\register[7][10] ), .A1N(
        n2501), .Y(n310) );
  OAI2BB2XL U2033 ( .B0(n2338), .B1(n2498), .A0N(\register[7][11] ), .A1N(
        n2501), .Y(n311) );
  OAI2BB2XL U2034 ( .B0(n2336), .B1(n2498), .A0N(\register[7][12] ), .A1N(
        n2501), .Y(n312) );
  OAI2BB2XL U2035 ( .B0(n2333), .B1(n2499), .A0N(\register[7][13] ), .A1N(
        n2501), .Y(n313) );
  OAI2BB2XL U2036 ( .B0(n2331), .B1(n2499), .A0N(\register[7][14] ), .A1N(
        n2501), .Y(n314) );
  OAI2BB2XL U2037 ( .B0(n2328), .B1(n2499), .A0N(\register[7][15] ), .A1N(
        n2500), .Y(n315) );
  OAI2BB2XL U2038 ( .B0(n2325), .B1(n2499), .A0N(\register[7][16] ), .A1N(
        n2501), .Y(n316) );
  OAI2BB2XL U2039 ( .B0(n2323), .B1(n2499), .A0N(\register[7][17] ), .A1N(
        n2500), .Y(n317) );
  OAI2BB2XL U2040 ( .B0(n2320), .B1(n2499), .A0N(\register[7][18] ), .A1N(
        n2500), .Y(n318) );
  OAI2BB2XL U2041 ( .B0(n2317), .B1(n2499), .A0N(\register[7][19] ), .A1N(
        n2500), .Y(n319) );
  OAI2BB2XL U2042 ( .B0(n2315), .B1(n2499), .A0N(\register[7][20] ), .A1N(
        n2500), .Y(n320) );
  OAI2BB2XL U2043 ( .B0(n2313), .B1(n2499), .A0N(\register[7][21] ), .A1N(
        n2500), .Y(n321) );
  OAI2BB2XL U2044 ( .B0(n2311), .B1(n2499), .A0N(\register[7][22] ), .A1N(
        n2501), .Y(n322) );
  OAI2BB2XL U2045 ( .B0(n2306), .B1(n2499), .A0N(\register[7][24] ), .A1N(
        n2501), .Y(n324) );
  OAI2BB2XL U2046 ( .B0(n2363), .B1(n2510), .A0N(\register[5][0] ), .A1N(n2508), .Y(n236) );
  OAI2BB2XL U2047 ( .B0(n2360), .B1(n2509), .A0N(\register[5][1] ), .A1N(n2508), .Y(n237) );
  OAI2BB2XL U2048 ( .B0(n2612), .B1(n2509), .A0N(\register[5][2] ), .A1N(n2508), .Y(n238) );
  OAI2BB2XL U2049 ( .B0(n2357), .B1(n2509), .A0N(\register[5][3] ), .A1N(n2512), .Y(n239) );
  OAI2BB2XL U2050 ( .B0(n2610), .B1(n2509), .A0N(\register[5][4] ), .A1N(n2508), .Y(n240) );
  OAI2BB2XL U2051 ( .B0(n2352), .B1(n2509), .A0N(\register[5][5] ), .A1N(n2512), .Y(n241) );
  OAI2BB2XL U2052 ( .B0(n2350), .B1(n2509), .A0N(\register[5][6] ), .A1N(n2512), .Y(n242) );
  OAI2BB2XL U2053 ( .B0(n2347), .B1(n2509), .A0N(\register[5][7] ), .A1N(n2512), .Y(n243) );
  OAI2BB2XL U2054 ( .B0(n2345), .B1(n2509), .A0N(\register[5][8] ), .A1N(n2512), .Y(n244) );
  OAI2BB2XL U2055 ( .B0(n2343), .B1(n2509), .A0N(\register[5][9] ), .A1N(n2512), .Y(n245) );
  OAI2BB2XL U2056 ( .B0(n2340), .B1(n2509), .A0N(\register[5][10] ), .A1N(
        n2512), .Y(n246) );
  OAI2BB2XL U2057 ( .B0(n2338), .B1(n2509), .A0N(\register[5][11] ), .A1N(
        n2512), .Y(n247) );
  OAI2BB2XL U2058 ( .B0(n2336), .B1(n2509), .A0N(\register[5][12] ), .A1N(
        n2512), .Y(n248) );
  OAI2BB2XL U2059 ( .B0(n2333), .B1(n2510), .A0N(\register[5][13] ), .A1N(
        n2512), .Y(n249) );
  OAI2BB2XL U2060 ( .B0(n2331), .B1(n2510), .A0N(\register[5][14] ), .A1N(
        n2512), .Y(n250) );
  OAI2BB2XL U2061 ( .B0(n2328), .B1(n2510), .A0N(\register[5][15] ), .A1N(
        n2511), .Y(n251) );
  OAI2BB2XL U2062 ( .B0(n2325), .B1(n2510), .A0N(\register[5][16] ), .A1N(
        n2512), .Y(n252) );
  OAI2BB2XL U2063 ( .B0(n2323), .B1(n2510), .A0N(\register[5][17] ), .A1N(
        n2511), .Y(n253) );
  OAI2BB2XL U2064 ( .B0(n2320), .B1(n2510), .A0N(\register[5][18] ), .A1N(
        n2511), .Y(n254) );
  OAI2BB2XL U2065 ( .B0(n2317), .B1(n2510), .A0N(\register[5][19] ), .A1N(
        n2511), .Y(n255) );
  OAI2BB2XL U2066 ( .B0(n2315), .B1(n2510), .A0N(\register[5][20] ), .A1N(
        n2511), .Y(n256) );
  OAI2BB2XL U2067 ( .B0(n2313), .B1(n2510), .A0N(\register[5][21] ), .A1N(
        n2511), .Y(n257) );
  OAI2BB2XL U2068 ( .B0(n2311), .B1(n2510), .A0N(\register[5][22] ), .A1N(
        n2512), .Y(n258) );
  OAI2BB2XL U2069 ( .B0(n2306), .B1(n2510), .A0N(\register[5][24] ), .A1N(
        n2512), .Y(n260) );
  NOR2BX1 U2070 ( .AN(n2147), .B(\register[3][0] ), .Y(n2101) );
  NOR2BX1 U2071 ( .AN(n2147), .B(\register[3][1] ), .Y(n2096) );
  NOR2BX1 U2072 ( .AN(n2147), .B(\register[3][2] ), .Y(n2091) );
  NOR2BX1 U2073 ( .AN(n2147), .B(\register[3][3] ), .Y(n2086) );
  NOR2BX1 U2074 ( .AN(n2147), .B(\register[3][4] ), .Y(n2081) );
  NOR2BX1 U2075 ( .AN(n2146), .B(\register[3][5] ), .Y(n2076) );
  NOR2BX1 U2076 ( .AN(n2147), .B(\register[3][6] ), .Y(n2071) );
  NOR2BX1 U2077 ( .AN(n2146), .B(\register[3][8] ), .Y(n2061) );
  NOR2BX1 U2078 ( .AN(n2146), .B(\register[3][9] ), .Y(n2056) );
  NOR2BX1 U2079 ( .AN(n2146), .B(\register[3][10] ), .Y(n2051) );
  NOR2BX1 U2080 ( .AN(n2146), .B(\register[3][11] ), .Y(n2046) );
  NOR2BX1 U2081 ( .AN(n2147), .B(\register[3][12] ), .Y(n2041) );
  NOR2BX1 U2082 ( .AN(n2146), .B(\register[3][13] ), .Y(n2036) );
  NOR2BX1 U2083 ( .AN(n2146), .B(\register[3][14] ), .Y(n2031) );
  NOR2BX1 U2084 ( .AN(n2146), .B(\register[3][15] ), .Y(n2026) );
  NOR2BX1 U2085 ( .AN(n2146), .B(\register[3][16] ), .Y(n2021) );
  NOR2BX1 U2086 ( .AN(n2146), .B(\register[3][17] ), .Y(n2016) );
  NOR2BX1 U2087 ( .AN(n2146), .B(\register[3][18] ), .Y(n2011) );
  NOR2BX1 U2088 ( .AN(n2146), .B(\register[3][19] ), .Y(n2006) );
  NOR2BX1 U2089 ( .AN(n2146), .B(\register[3][21] ), .Y(n1996) );
  NOR2BX1 U2090 ( .AN(n2146), .B(\register[3][22] ), .Y(n1991) );
  NOR2BX1 U2091 ( .AN(n2146), .B(\register[3][23] ), .Y(n1986) );
  NOR2BX1 U2092 ( .AN(n2146), .B(\register[3][24] ), .Y(n1981) );
  NOR2BX1 U2093 ( .AN(n2147), .B(\register[3][25] ), .Y(n1976) );
  NOR2BX1 U2094 ( .AN(n2147), .B(\register[3][26] ), .Y(n1971) );
  NOR2BX1 U2095 ( .AN(n2147), .B(\register[3][27] ), .Y(n1966) );
  NOR2BX1 U2096 ( .AN(n2147), .B(\register[3][28] ), .Y(n1961) );
  NOR2BX1 U2097 ( .AN(n2147), .B(\register[3][29] ), .Y(n1956) );
  NOR2BX1 U2098 ( .AN(n2147), .B(\register[3][30] ), .Y(n1951) );
  NOR2BX1 U2099 ( .AN(n2147), .B(\register[3][31] ), .Y(n1946) );
  NOR2BX1 U2100 ( .AN(n1596), .B(\register[3][0] ), .Y(n1551) );
  NOR2BX1 U2101 ( .AN(n1596), .B(\register[3][2] ), .Y(n1541) );
  NOR2BX1 U2102 ( .AN(n1595), .B(\register[3][8] ), .Y(n1511) );
  NOR2BX1 U2103 ( .AN(n1595), .B(\register[3][10] ), .Y(n1501) );
  NOR2BX1 U2104 ( .AN(n1595), .B(\register[3][11] ), .Y(n1496) );
  NOR2BX1 U2105 ( .AN(n1596), .B(\register[3][12] ), .Y(n1491) );
  NOR2BX1 U2106 ( .AN(n1595), .B(\register[3][13] ), .Y(n1486) );
  NOR2BX1 U2107 ( .AN(n1595), .B(\register[3][15] ), .Y(n1476) );
  NOR2BX1 U2108 ( .AN(n1595), .B(\register[3][16] ), .Y(n1471) );
  NOR2BX1 U2109 ( .AN(n1595), .B(\register[3][17] ), .Y(n1466) );
  NOR2BX1 U2110 ( .AN(n1595), .B(\register[3][18] ), .Y(n1461) );
  NOR2BX1 U2111 ( .AN(n1595), .B(\register[3][19] ), .Y(n1456) );
  NOR2BX1 U2112 ( .AN(n1595), .B(\register[3][20] ), .Y(n1451) );
  NOR2BX1 U2113 ( .AN(n1595), .B(\register[3][21] ), .Y(n1446) );
  NOR2BX1 U2114 ( .AN(n1595), .B(\register[3][22] ), .Y(n1441) );
  NOR2BX1 U2115 ( .AN(n1595), .B(\register[3][23] ), .Y(n1436) );
  NOR2BX1 U2116 ( .AN(n1595), .B(\register[3][24] ), .Y(n1431) );
  NOR2BX1 U2117 ( .AN(n1596), .B(\register[3][25] ), .Y(n1426) );
  NOR2BX1 U2118 ( .AN(n1596), .B(\register[3][26] ), .Y(n1421) );
  NOR2BX1 U2119 ( .AN(n1596), .B(\register[3][27] ), .Y(n1416) );
  NOR2BX1 U2120 ( .AN(n1596), .B(\register[3][28] ), .Y(n1411) );
  NOR2BX1 U2121 ( .AN(n1596), .B(\register[3][29] ), .Y(n1406) );
  NOR2BX1 U2122 ( .AN(n1596), .B(\register[3][30] ), .Y(n1401) );
  NOR2BX1 U2123 ( .AN(n1596), .B(\register[3][31] ), .Y(n1396) );
  NOR2X1 U2124 ( .A(n1600), .B(\register[1][26] ), .Y(n1423) );
  NAND2X1 U2125 ( .A(n2100), .B(n2099), .Y(n1705) );
  NOR2X1 U2126 ( .A(n2098), .B(n2097), .Y(n2100) );
  MXI2X1 U2127 ( .A(n2552), .B(n2096), .S0(n2172), .Y(n2099) );
  NOR2X1 U2128 ( .A(n2149), .B(\register[1][1] ), .Y(n2098) );
  NAND2X1 U2129 ( .A(n1550), .B(n1549), .Y(n1155) );
  NOR2X1 U2130 ( .A(n1548), .B(n1547), .Y(n1550) );
  NOR2X1 U2131 ( .A(n1598), .B(\register[1][1] ), .Y(n1548) );
  NAND2X1 U2132 ( .A(n2095), .B(n2094), .Y(n1713) );
  NOR2X1 U2133 ( .A(n2093), .B(n2092), .Y(n2095) );
  MXI2X1 U2134 ( .A(n2553), .B(n2091), .S0(n2173), .Y(n2094) );
  NOR2X1 U2135 ( .A(n2149), .B(\register[1][2] ), .Y(n2093) );
  NAND2X1 U2136 ( .A(n2090), .B(n2089), .Y(n1721) );
  NOR2X1 U2137 ( .A(n2088), .B(n2087), .Y(n2090) );
  MXI2X1 U2138 ( .A(n2554), .B(n2086), .S0(n2173), .Y(n2089) );
  NOR2X1 U2139 ( .A(n2148), .B(\register[1][3] ), .Y(n2088) );
  NAND2X1 U2140 ( .A(n2085), .B(n2084), .Y(n1729) );
  NOR2X1 U2141 ( .A(n2083), .B(n2082), .Y(n2085) );
  MXI2X1 U2142 ( .A(n2555), .B(n2081), .S0(n2173), .Y(n2084) );
  NOR2X1 U2143 ( .A(n2147), .B(\register[1][4] ), .Y(n2083) );
  NAND2X1 U2144 ( .A(n2080), .B(n2079), .Y(n1737) );
  NOR2X1 U2145 ( .A(n2078), .B(n2077), .Y(n2080) );
  MXI2X1 U2146 ( .A(n2556), .B(n2076), .S0(n2173), .Y(n2079) );
  NOR2X1 U2147 ( .A(n2148), .B(\register[1][5] ), .Y(n2078) );
  NAND2X1 U2148 ( .A(n2075), .B(n2074), .Y(n1745) );
  NOR2X1 U2149 ( .A(n2073), .B(n2072), .Y(n2075) );
  MXI2X1 U2150 ( .A(n2557), .B(n2071), .S0(n2173), .Y(n2074) );
  NOR2X1 U2151 ( .A(n2147), .B(\register[1][6] ), .Y(n2073) );
  NAND2X1 U2152 ( .A(n2070), .B(n2069), .Y(n1753) );
  NOR2X1 U2153 ( .A(n2068), .B(n2067), .Y(n2070) );
  NOR2X1 U2154 ( .A(n2148), .B(\register[1][7] ), .Y(n2068) );
  NAND2X1 U2155 ( .A(n2065), .B(n2064), .Y(n1761) );
  NOR2X1 U2156 ( .A(n2063), .B(n2062), .Y(n2065) );
  MXI2X1 U2157 ( .A(n2559), .B(n2061), .S0(n2173), .Y(n2064) );
  NOR2X1 U2158 ( .A(n2149), .B(\register[1][8] ), .Y(n2063) );
  NAND2X1 U2159 ( .A(n2060), .B(n2059), .Y(n1769) );
  NOR2X1 U2160 ( .A(n2058), .B(n2057), .Y(n2060) );
  MXI2X1 U2161 ( .A(n2560), .B(n2056), .S0(n2173), .Y(n2059) );
  NOR2X1 U2162 ( .A(n2148), .B(\register[1][9] ), .Y(n2058) );
  NAND2X1 U2163 ( .A(n2055), .B(n2054), .Y(n1777) );
  NOR2X1 U2164 ( .A(n2053), .B(n2052), .Y(n2055) );
  MXI2X1 U2165 ( .A(n2561), .B(n2051), .S0(n2173), .Y(n2054) );
  NOR2X1 U2166 ( .A(n2148), .B(\register[1][10] ), .Y(n2053) );
  NAND2X1 U2167 ( .A(n2050), .B(n2049), .Y(n1785) );
  NOR2X1 U2168 ( .A(n2048), .B(n2047), .Y(n2050) );
  MXI2X1 U2169 ( .A(n2562), .B(n2046), .S0(n2173), .Y(n2049) );
  NOR2X1 U2170 ( .A(n2149), .B(\register[1][11] ), .Y(n2048) );
  NAND2X1 U2171 ( .A(n2045), .B(n2044), .Y(n1793) );
  NOR2X1 U2172 ( .A(n2043), .B(n2042), .Y(n2045) );
  MXI2X1 U2173 ( .A(n2563), .B(n2041), .S0(n2173), .Y(n2044) );
  NOR2X1 U2174 ( .A(n2149), .B(\register[1][12] ), .Y(n2043) );
  NAND2X1 U2175 ( .A(n2040), .B(n2039), .Y(n1801) );
  NOR2X1 U2176 ( .A(n2038), .B(n2037), .Y(n2040) );
  MXI2X1 U2177 ( .A(n2564), .B(n2036), .S0(n2173), .Y(n2039) );
  NOR2X1 U2178 ( .A(n2149), .B(\register[1][13] ), .Y(n2038) );
  NAND2X1 U2179 ( .A(n2035), .B(n2034), .Y(n1809) );
  NOR2X1 U2180 ( .A(n2033), .B(n2032), .Y(n2035) );
  MXI2X1 U2181 ( .A(n2565), .B(n2031), .S0(n2173), .Y(n2034) );
  NOR2X1 U2182 ( .A(n2149), .B(\register[1][14] ), .Y(n2033) );
  NAND2X1 U2183 ( .A(n2030), .B(n2029), .Y(n1817) );
  NOR2X1 U2184 ( .A(n2028), .B(n2027), .Y(n2030) );
  MXI2X1 U2185 ( .A(n2566), .B(n2026), .S0(n2174), .Y(n2029) );
  NOR2X1 U2186 ( .A(n2150), .B(\register[1][15] ), .Y(n2028) );
  NAND2X1 U2187 ( .A(n2025), .B(n2024), .Y(n1825) );
  NOR2X1 U2188 ( .A(n2023), .B(n2022), .Y(n2025) );
  MXI2X1 U2189 ( .A(n2567), .B(n2021), .S0(n2174), .Y(n2024) );
  NOR2X1 U2190 ( .A(n2150), .B(\register[1][16] ), .Y(n2023) );
  NAND2X1 U2191 ( .A(n2020), .B(n2019), .Y(n1833) );
  NOR2X1 U2192 ( .A(n2018), .B(n2017), .Y(n2020) );
  MXI2X1 U2193 ( .A(n2568), .B(n2016), .S0(n2174), .Y(n2019) );
  NOR2X1 U2194 ( .A(n2150), .B(\register[1][17] ), .Y(n2018) );
  NAND2X1 U2195 ( .A(n2015), .B(n2014), .Y(n1841) );
  NOR2X1 U2196 ( .A(n2013), .B(n2012), .Y(n2015) );
  MXI2X1 U2197 ( .A(n2569), .B(n2011), .S0(n2174), .Y(n2014) );
  NOR2X1 U2198 ( .A(n2150), .B(\register[1][18] ), .Y(n2013) );
  NAND2X1 U2199 ( .A(n2010), .B(n2009), .Y(n1849) );
  NOR2X1 U2200 ( .A(n2008), .B(n2007), .Y(n2010) );
  MXI2X1 U2201 ( .A(n2570), .B(n2006), .S0(n2174), .Y(n2009) );
  NOR2X1 U2202 ( .A(n2150), .B(\register[1][19] ), .Y(n2008) );
  NAND2X1 U2203 ( .A(n2005), .B(n2004), .Y(n1857) );
  NOR2X1 U2204 ( .A(n2003), .B(n2002), .Y(n2005) );
  NAND2X1 U2205 ( .A(n2000), .B(n1999), .Y(n1865) );
  NOR2X1 U2206 ( .A(n1998), .B(n1997), .Y(n2000) );
  MXI2X1 U2207 ( .A(n2572), .B(n1996), .S0(n2174), .Y(n1999) );
  NOR2X1 U2208 ( .A(n2151), .B(\register[1][21] ), .Y(n1998) );
  NAND2X1 U2209 ( .A(n1995), .B(n1994), .Y(n1873) );
  NOR2X1 U2210 ( .A(n1993), .B(n1992), .Y(n1995) );
  MXI2X1 U2211 ( .A(n2573), .B(n1991), .S0(n2174), .Y(n1994) );
  NOR2X1 U2212 ( .A(n2151), .B(\register[1][22] ), .Y(n1993) );
  NAND2X1 U2213 ( .A(n1990), .B(n1989), .Y(n1881) );
  NOR2X1 U2214 ( .A(n1988), .B(n1987), .Y(n1990) );
  MXI2X1 U2215 ( .A(n2574), .B(n1986), .S0(n2174), .Y(n1989) );
  NOR2X1 U2216 ( .A(n2151), .B(\register[1][23] ), .Y(n1988) );
  NAND2X1 U2217 ( .A(n1985), .B(n1984), .Y(n1889) );
  NOR2X1 U2218 ( .A(n1983), .B(n1982), .Y(n1985) );
  MXI2X1 U2219 ( .A(n2575), .B(n1981), .S0(n2174), .Y(n1984) );
  NOR2X1 U2220 ( .A(n2151), .B(\register[1][24] ), .Y(n1983) );
  NAND2X1 U2221 ( .A(n1975), .B(n1974), .Y(n1905) );
  NOR2X1 U2222 ( .A(n1973), .B(n1972), .Y(n1975) );
  MXI2X1 U2223 ( .A(n2577), .B(n1971), .S0(n2174), .Y(n1974) );
  NOR2X1 U2224 ( .A(n2151), .B(\register[1][26] ), .Y(n1973) );
  NAND2X1 U2225 ( .A(n1960), .B(n1959), .Y(n1929) );
  NOR2X1 U2226 ( .A(n1958), .B(n1957), .Y(n1960) );
  MXI2X1 U2227 ( .A(n2580), .B(n1956), .S0(n2174), .Y(n1959) );
  NOR2X1 U2228 ( .A(n2129), .B(\register[1][29] ), .Y(n1958) );
  NAND2X1 U2229 ( .A(n1950), .B(n1949), .Y(n1945) );
  NOR2X1 U2230 ( .A(n1948), .B(n1947), .Y(n1950) );
  MXI2X1 U2231 ( .A(n2582), .B(n1946), .S0(n2174), .Y(n1949) );
  NOR2X1 U2232 ( .A(n2137), .B(\register[1][31] ), .Y(n1948) );
  NAND2X1 U2233 ( .A(n1545), .B(n1544), .Y(n1163) );
  NOR2X1 U2234 ( .A(n1543), .B(n1542), .Y(n1545) );
  MXI2X1 U2235 ( .A(n2553), .B(n1541), .S0(n1621), .Y(n1544) );
  NOR2X1 U2236 ( .A(n1598), .B(\register[1][2] ), .Y(n1543) );
  NAND2X1 U2237 ( .A(n1540), .B(n1539), .Y(n1171) );
  NOR2X1 U2238 ( .A(n1538), .B(n1537), .Y(n1540) );
  NAND2X1 U2239 ( .A(n1535), .B(n1534), .Y(n1179) );
  NOR2X1 U2240 ( .A(n1533), .B(n1532), .Y(n1535) );
  MXI2X1 U2241 ( .A(n2555), .B(n1531), .S0(n1621), .Y(n1534) );
  NAND2X1 U2242 ( .A(n1530), .B(n1529), .Y(n1187) );
  NOR2X1 U2243 ( .A(n1528), .B(n1527), .Y(n1530) );
  NAND2X1 U2244 ( .A(n1525), .B(n1524), .Y(n1195) );
  NOR2X1 U2245 ( .A(n1523), .B(n1522), .Y(n1525) );
  MXI2X1 U2246 ( .A(n2557), .B(n1521), .S0(n1621), .Y(n1524) );
  NAND2X1 U2247 ( .A(n1520), .B(n1519), .Y(n1203) );
  NOR2X1 U2248 ( .A(n1518), .B(n1517), .Y(n1520) );
  NAND2X1 U2249 ( .A(n1515), .B(n1514), .Y(n1211) );
  NOR2X1 U2250 ( .A(n1513), .B(n1512), .Y(n1515) );
  MXI2X1 U2251 ( .A(n2559), .B(n1511), .S0(n1621), .Y(n1514) );
  NOR2X1 U2252 ( .A(n1598), .B(\register[1][8] ), .Y(n1513) );
  NAND2X1 U2253 ( .A(n1510), .B(n1509), .Y(n1219) );
  NOR2X1 U2254 ( .A(n1508), .B(n1507), .Y(n1510) );
  NAND2X1 U2255 ( .A(n1505), .B(n1504), .Y(n1227) );
  NOR2X1 U2256 ( .A(n1503), .B(n1502), .Y(n1505) );
  MXI2X1 U2257 ( .A(n2561), .B(n1501), .S0(n1621), .Y(n1504) );
  NOR2X1 U2258 ( .A(n1597), .B(\register[1][10] ), .Y(n1503) );
  NAND2X1 U2259 ( .A(n1500), .B(n1499), .Y(n1235) );
  NOR2X1 U2260 ( .A(n1498), .B(n1497), .Y(n1500) );
  MXI2X1 U2261 ( .A(n2562), .B(n1496), .S0(n1621), .Y(n1499) );
  NOR2X1 U2262 ( .A(n1598), .B(\register[1][11] ), .Y(n1498) );
  NAND2X1 U2263 ( .A(n1495), .B(n1494), .Y(n1243) );
  NOR2X1 U2264 ( .A(n1493), .B(n1492), .Y(n1495) );
  MXI2X1 U2265 ( .A(n2563), .B(n1491), .S0(n1621), .Y(n1494) );
  NOR2X1 U2266 ( .A(n1598), .B(\register[1][12] ), .Y(n1493) );
  NAND2X1 U2267 ( .A(n1490), .B(n1489), .Y(n1251) );
  NOR2X1 U2268 ( .A(n1488), .B(n1487), .Y(n1490) );
  MXI2X1 U2269 ( .A(n2564), .B(n1486), .S0(n1621), .Y(n1489) );
  NOR2X1 U2270 ( .A(n1598), .B(\register[1][13] ), .Y(n1488) );
  NAND2X1 U2271 ( .A(n1485), .B(n1484), .Y(n1259) );
  NOR2X1 U2272 ( .A(n1483), .B(n1482), .Y(n1485) );
  NOR2X1 U2273 ( .A(n1598), .B(\register[1][14] ), .Y(n1483) );
  NAND2X1 U2274 ( .A(n1480), .B(n1479), .Y(n1267) );
  NOR2X1 U2275 ( .A(n1478), .B(n1477), .Y(n1480) );
  MXI2X1 U2276 ( .A(n2566), .B(n1476), .S0(n1622), .Y(n1479) );
  NOR2X1 U2277 ( .A(n1599), .B(\register[1][15] ), .Y(n1478) );
  NAND2X1 U2278 ( .A(n1475), .B(n1474), .Y(n1275) );
  NOR2X1 U2279 ( .A(n1473), .B(n1472), .Y(n1475) );
  MXI2X1 U2280 ( .A(n2567), .B(n1471), .S0(n1622), .Y(n1474) );
  NOR2X1 U2281 ( .A(n1599), .B(\register[1][16] ), .Y(n1473) );
  NAND2X1 U2282 ( .A(n1470), .B(n1469), .Y(n1283) );
  NOR2X1 U2283 ( .A(n1468), .B(n1467), .Y(n1470) );
  MXI2X1 U2284 ( .A(n2568), .B(n1466), .S0(n1622), .Y(n1469) );
  NOR2X1 U2285 ( .A(n1599), .B(\register[1][17] ), .Y(n1468) );
  NAND2X1 U2286 ( .A(n1465), .B(n1464), .Y(n1291) );
  NOR2X1 U2287 ( .A(n1463), .B(n1462), .Y(n1465) );
  MXI2X1 U2288 ( .A(n2569), .B(n1461), .S0(n1622), .Y(n1464) );
  NOR2X1 U2289 ( .A(n1599), .B(\register[1][18] ), .Y(n1463) );
  NAND2X1 U2290 ( .A(n1460), .B(n1459), .Y(n1299) );
  NOR2X1 U2291 ( .A(n1458), .B(n1457), .Y(n1460) );
  MXI2X1 U2292 ( .A(n2570), .B(n1456), .S0(n1622), .Y(n1459) );
  NOR2X1 U2293 ( .A(n1599), .B(\register[1][19] ), .Y(n1458) );
  NAND2X1 U2294 ( .A(n1455), .B(n1454), .Y(n1307) );
  NOR2X1 U2295 ( .A(n1453), .B(n1452), .Y(n1455) );
  MXI2X1 U2296 ( .A(n2571), .B(n1451), .S0(n1622), .Y(n1454) );
  NOR2X1 U2297 ( .A(n1599), .B(\register[1][20] ), .Y(n1453) );
  NAND2X1 U2298 ( .A(n1450), .B(n1449), .Y(n1315) );
  NOR2X1 U2299 ( .A(n1448), .B(n1447), .Y(n1450) );
  MXI2X1 U2300 ( .A(n2572), .B(n1446), .S0(n1622), .Y(n1449) );
  NOR2X1 U2301 ( .A(n1600), .B(\register[1][21] ), .Y(n1448) );
  NAND2X1 U2302 ( .A(n1445), .B(n1444), .Y(n1323) );
  NOR2X1 U2303 ( .A(n1443), .B(n1442), .Y(n1445) );
  MXI2X1 U2304 ( .A(n2573), .B(n1441), .S0(n1622), .Y(n1444) );
  NOR2X1 U2305 ( .A(n1600), .B(\register[1][22] ), .Y(n1443) );
  NAND2X1 U2306 ( .A(n1440), .B(n1439), .Y(n1331) );
  NOR2X1 U2307 ( .A(n1438), .B(n1437), .Y(n1440) );
  MXI2X1 U2308 ( .A(n2574), .B(n1436), .S0(n1622), .Y(n1439) );
  NOR2X1 U2309 ( .A(n1600), .B(\register[1][23] ), .Y(n1438) );
  NAND2X1 U2310 ( .A(n1435), .B(n1434), .Y(n1339) );
  NOR2X1 U2311 ( .A(n1433), .B(n1432), .Y(n1435) );
  MXI2X1 U2312 ( .A(n2575), .B(n1431), .S0(n1622), .Y(n1434) );
  NOR2X1 U2313 ( .A(n1600), .B(\register[1][24] ), .Y(n1433) );
  NAND2X1 U2314 ( .A(n1425), .B(n1424), .Y(n1355) );
  NOR2X1 U2315 ( .A(n1423), .B(n1422), .Y(n1425) );
  MXI2X1 U2316 ( .A(n2577), .B(n1421), .S0(n1622), .Y(n1424) );
  NOR2X1 U2317 ( .A(n1594), .B(n1624), .Y(n1422) );
  NAND2X1 U2318 ( .A(n1410), .B(n1409), .Y(n1379) );
  NOR2X1 U2319 ( .A(n1408), .B(n1407), .Y(n1410) );
  MXI2X1 U2320 ( .A(n2580), .B(n1406), .S0(n1622), .Y(n1409) );
  NOR2X1 U2321 ( .A(n1578), .B(\register[1][29] ), .Y(n1408) );
  NAND2X1 U2322 ( .A(n1400), .B(n1399), .Y(n1395) );
  NOR2X1 U2323 ( .A(n1398), .B(n1397), .Y(n1400) );
  MXI2X1 U2324 ( .A(n2582), .B(n1396), .S0(n1622), .Y(n1399) );
  NOR2X1 U2325 ( .A(n1578), .B(\register[1][31] ), .Y(n1398) );
  NAND2X1 U2326 ( .A(n2105), .B(n2104), .Y(n1697) );
  NOR2X1 U2327 ( .A(n2103), .B(n2102), .Y(n2105) );
  MXI2X1 U2328 ( .A(n2551), .B(n2101), .S0(n2175), .Y(n2104) );
  NOR2X1 U2329 ( .A(n2143), .B(\register[1][0] ), .Y(n2103) );
  NAND2X1 U2330 ( .A(n1980), .B(n1979), .Y(n1897) );
  NOR2X1 U2331 ( .A(n1978), .B(n1977), .Y(n1980) );
  MXI2X1 U2332 ( .A(n2576), .B(n1976), .S0(n2175), .Y(n1979) );
  NOR2X1 U2333 ( .A(n2151), .B(\register[1][25] ), .Y(n1978) );
  NAND2X1 U2334 ( .A(n1970), .B(n1969), .Y(n1913) );
  NOR2X1 U2335 ( .A(n1968), .B(n1967), .Y(n1970) );
  MXI2X1 U2336 ( .A(n2578), .B(n1966), .S0(n2175), .Y(n1969) );
  NOR2X1 U2337 ( .A(n2129), .B(\register[1][27] ), .Y(n1968) );
  NAND2X1 U2338 ( .A(n1965), .B(n1964), .Y(n1921) );
  NOR2X1 U2339 ( .A(n1963), .B(n1962), .Y(n1965) );
  MXI2X1 U2340 ( .A(n2579), .B(n1961), .S0(n2175), .Y(n1964) );
  NOR2X1 U2341 ( .A(n2137), .B(\register[1][28] ), .Y(n1963) );
  NAND2X1 U2342 ( .A(n1955), .B(n1954), .Y(n1937) );
  NOR2X1 U2343 ( .A(n1953), .B(n1952), .Y(n1955) );
  MXI2X1 U2344 ( .A(n2581), .B(n1951), .S0(n2175), .Y(n1954) );
  NOR2X1 U2345 ( .A(n2129), .B(\register[1][30] ), .Y(n1953) );
  NAND2X1 U2346 ( .A(n1555), .B(n1554), .Y(n1147) );
  NOR2X1 U2347 ( .A(n1553), .B(n1552), .Y(n1555) );
  MXI2X1 U2348 ( .A(n2551), .B(n1551), .S0(n1623), .Y(n1554) );
  NOR2X1 U2349 ( .A(n1578), .B(\register[1][0] ), .Y(n1553) );
  NAND2X1 U2350 ( .A(n1430), .B(n1429), .Y(n1347) );
  NOR2X1 U2351 ( .A(n1428), .B(n1427), .Y(n1430) );
  MXI2X1 U2352 ( .A(n2576), .B(n1426), .S0(n1623), .Y(n1429) );
  NOR2X1 U2353 ( .A(n1600), .B(\register[1][25] ), .Y(n1428) );
  NAND2X1 U2354 ( .A(n1420), .B(n1419), .Y(n1363) );
  NOR2X1 U2355 ( .A(n1418), .B(n1417), .Y(n1420) );
  MXI2X1 U2356 ( .A(n2578), .B(n1416), .S0(n1623), .Y(n1419) );
  NOR2X1 U2357 ( .A(n1578), .B(\register[1][27] ), .Y(n1418) );
  NAND2X1 U2358 ( .A(n1415), .B(n1414), .Y(n1371) );
  NOR2X1 U2359 ( .A(n1413), .B(n1412), .Y(n1415) );
  MXI2X1 U2360 ( .A(n2579), .B(n1411), .S0(n1623), .Y(n1414) );
  NOR2X1 U2361 ( .A(n1578), .B(\register[1][28] ), .Y(n1413) );
  NAND2X1 U2362 ( .A(n1405), .B(n1404), .Y(n1387) );
  NOR2X1 U2363 ( .A(n1403), .B(n1402), .Y(n1405) );
  MXI2X1 U2364 ( .A(n2581), .B(n1401), .S0(n1623), .Y(n1404) );
  NOR2X1 U2365 ( .A(n1594), .B(\register[1][30] ), .Y(n1403) );
  MXI4X1 U2366 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n2165), .S1(n2141), .Y(
        n1696) );
  MXI4X1 U2367 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n2165), .S1(n2141), .Y(
        n1692) );
  MXI4X1 U2368 ( .A(\register[20][1] ), .B(\register[21][1] ), .C(
        \register[22][1] ), .D(\register[23][1] ), .S0(n2166), .S1(n2141), .Y(
        n1700) );
  MXI4X1 U2369 ( .A(\register[4][1] ), .B(\register[5][1] ), .C(
        \register[6][1] ), .D(\register[7][1] ), .S0(n2166), .S1(n2141), .Y(
        n1704) );
  MXI4X1 U2370 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n2166), .S1(n2141), .Y(
        n1708) );
  MXI4X1 U2371 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n2166), .S1(n2141), .Y(
        n1712) );
  MXI4X1 U2372 ( .A(\register[20][3] ), .B(\register[21][3] ), .C(
        \register[22][3] ), .D(\register[23][3] ), .S0(n2166), .S1(n2142), .Y(
        n1716) );
  MXI4X1 U2373 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n2167), .S1(n2142), .Y(
        n1720) );
  MXI4X1 U2374 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n2167), .S1(n2142), .Y(
        n1724) );
  MXI4X1 U2375 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n2167), .S1(n2142), .Y(
        n1728) );
  MXI4X1 U2376 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n2168), .S1(n2142), .Y(
        n1736) );
  MXI4X1 U2377 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n2167), .S1(n2142), .Y(
        n1732) );
  MXI4X1 U2378 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n2168), .S1(n2143), .Y(
        n1740) );
  MXI4X1 U2379 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n2168), .S1(n2143), .Y(
        n1744) );
  MXI4X1 U2380 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n2169), .S1(n2143), .Y(
        n1760) );
  MXI4X1 U2381 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n2169), .S1(n2143), .Y(
        n1756) );
  MXI4X1 U2382 ( .A(\register[4][9] ), .B(\register[5][9] ), .C(
        \register[6][9] ), .D(\register[7][9] ), .S0(n2170), .S1(n2144), .Y(
        n1768) );
  MXI4X1 U2383 ( .A(\register[20][9] ), .B(\register[21][9] ), .C(
        \register[22][9] ), .D(\register[23][9] ), .S0(n2169), .S1(n2144), .Y(
        n1764) );
  MXI4X1 U2384 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n2170), .S1(n2144), .Y(
        n1776) );
  MXI4X1 U2385 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1772) );
  MXI4X1 U2386 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n2171), .S1(n2144), .Y(
        n1784) );
  MXI4X1 U2387 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1780) );
  MXI4X1 U2388 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n2171), .S1(n2145), 
        .Y(n1788) );
  MXI4X1 U2389 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n2169), .S1(n2143), .Y(
        n1792) );
  MXI4X1 U2390 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n2171), .S1(n2145), .Y(
        n1800) );
  MXI4X1 U2391 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1796) );
  MXI4X1 U2392 ( .A(\register[20][14] ), .B(\register[21][14] ), .C(
        \register[22][14] ), .D(\register[23][14] ), .S0(n2172), .S1(n2145), 
        .Y(n1804) );
  MXI4X1 U2393 ( .A(\register[4][14] ), .B(\register[5][14] ), .C(
        \register[6][14] ), .D(\register[7][14] ), .S0(n2172), .S1(n2145), .Y(
        n1808) );
  MXI4X1 U2394 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n2172), .S1(n2145), 
        .Y(n1812) );
  MXI4X1 U2395 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n2169), .S1(n2143), .Y(
        n1816) );
  MXI4X1 U2396 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n2158), .S1(n2136), .Y(
        n1824) );
  MXI4X1 U2397 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1820) );
  MXI4X1 U2398 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n2158), .S1(n2136), .Y(
        n1832) );
  MXI4X1 U2399 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1828) );
  MXI4X1 U2400 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n2159), .S1(n2136), .Y(
        n1840) );
  MXI4X1 U2401 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n2159), .S1(n2136), 
        .Y(n1836) );
  MXI4X1 U2402 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n2159), .S1(n2137), .Y(
        n1848) );
  MXI4X1 U2403 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n2159), .S1(n2137), 
        .Y(n1844) );
  MXI4X1 U2404 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n2160), .S1(n2137), .Y(
        n1864) );
  MXI4X1 U2405 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1860) );
  MXI4X1 U2406 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n2161), .S1(n2138), .Y(
        n1872) );
  MXI4X1 U2407 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n2160), .S1(n2138), 
        .Y(n1868) );
  MXI4X1 U2408 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n2161), .S1(n2138), .Y(
        n1880) );
  MXI4X1 U2409 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1876) );
  MXI4X1 U2410 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n2162), .S1(n2138), .Y(
        n1888) );
  MXI4X1 U2411 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n2161), .S1(n2138), 
        .Y(n1884) );
  MXI4X1 U2412 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n2162), .S1(n2139), .Y(
        n1896) );
  MXI4X1 U2413 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n2162), .S1(n2139), 
        .Y(n1892) );
  MXI4X1 U2414 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n2163), .S1(n2139), .Y(
        n1904) );
  MXI4X1 U2415 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n2162), .S1(n2139), 
        .Y(n1900) );
  MXI4X1 U2416 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n2163), .S1(n2139), .Y(
        n1912) );
  MXI4X1 U2417 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1908) );
  MXI4X1 U2418 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n2164), .S1(n2140), .Y(
        n1920) );
  MXI4X1 U2419 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n2163), .S1(n2139), 
        .Y(n1916) );
  MXI4X1 U2420 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n2164), .S1(n2140), .Y(
        n1928) );
  MXI4X1 U2421 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1924) );
  MXI4X1 U2422 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n2165), .S1(n2140), .Y(
        n1936) );
  MXI4X1 U2423 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1932) );
  MXI4X1 U2424 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n2165), .S1(n2140), 
        .Y(n1940) );
  MXI4X1 U2425 ( .A(\register[4][0] ), .B(\register[5][0] ), .C(
        \register[6][0] ), .D(\register[7][0] ), .S0(n1615), .S1(n1590), .Y(
        n1146) );
  MXI4X1 U2426 ( .A(\register[20][0] ), .B(\register[21][0] ), .C(
        \register[22][0] ), .D(\register[23][0] ), .S0(n1615), .S1(n1590), .Y(
        n1142) );
  MXI4X1 U2427 ( .A(\register[20][2] ), .B(\register[21][2] ), .C(
        \register[22][2] ), .D(\register[23][2] ), .S0(n1616), .S1(n1590), .Y(
        n1158) );
  MXI4X1 U2428 ( .A(\register[4][2] ), .B(\register[5][2] ), .C(
        \register[6][2] ), .D(\register[7][2] ), .S0(n1616), .S1(n1590), .Y(
        n1162) );
  MXI4X1 U2429 ( .A(\register[4][3] ), .B(\register[5][3] ), .C(
        \register[6][3] ), .D(\register[7][3] ), .S0(n1617), .S1(n1591), .Y(
        n1170) );
  MXI4X1 U2430 ( .A(\register[20][4] ), .B(\register[21][4] ), .C(
        \register[22][4] ), .D(\register[23][4] ), .S0(n1617), .S1(n1591), .Y(
        n1174) );
  MXI4X1 U2431 ( .A(\register[4][4] ), .B(\register[5][4] ), .C(
        \register[6][4] ), .D(\register[7][4] ), .S0(n1617), .S1(n1591), .Y(
        n1178) );
  MXI4X1 U2432 ( .A(\register[4][5] ), .B(\register[5][5] ), .C(
        \register[6][5] ), .D(\register[7][5] ), .S0(n1624), .S1(n1591), .Y(
        n1186) );
  MXI4X1 U2433 ( .A(\register[20][5] ), .B(\register[21][5] ), .C(
        \register[22][5] ), .D(\register[23][5] ), .S0(n1617), .S1(n1591), .Y(
        n1182) );
  MXI4X1 U2434 ( .A(\register[20][6] ), .B(\register[21][6] ), .C(
        \register[22][6] ), .D(\register[23][6] ), .S0(n1624), .S1(n1592), .Y(
        n1190) );
  MXI4X1 U2435 ( .A(\register[4][6] ), .B(\register[5][6] ), .C(
        \register[6][6] ), .D(\register[7][6] ), .S0(n1624), .S1(n1592), .Y(
        n1194) );
  MXI4X1 U2436 ( .A(\register[20][7] ), .B(\register[21][7] ), .C(
        \register[22][7] ), .D(\register[23][7] ), .S0(n1624), .S1(n1592), .Y(
        n1198) );
  MXI4X1 U2437 ( .A(\register[20][8] ), .B(\register[21][8] ), .C(
        \register[22][8] ), .D(\register[23][8] ), .S0(n1624), .S1(n1592), .Y(
        n1206) );
  MXI4X1 U2438 ( .A(\register[4][8] ), .B(\register[5][8] ), .C(
        \register[6][8] ), .D(\register[7][8] ), .S0(n1624), .S1(n1592), .Y(
        n1210) );
  MXI4X1 U2439 ( .A(\register[4][10] ), .B(\register[5][10] ), .C(
        \register[6][10] ), .D(\register[7][10] ), .S0(n1618), .S1(n1593), .Y(
        n1226) );
  MXI4X1 U2440 ( .A(\register[20][10] ), .B(\register[21][10] ), .C(
        \register[22][10] ), .D(\register[23][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1222) );
  MXI4X1 U2441 ( .A(\register[4][11] ), .B(\register[5][11] ), .C(
        \register[6][11] ), .D(\register[7][11] ), .S0(n1619), .S1(n1593), .Y(
        n1234) );
  MXI4X1 U2442 ( .A(\register[20][11] ), .B(\register[21][11] ), .C(
        \register[22][11] ), .D(\register[23][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1230) );
  MXI4X1 U2443 ( .A(\register[20][12] ), .B(\register[21][12] ), .C(
        \register[22][12] ), .D(\register[23][12] ), .S0(n1619), .S1(n1594), 
        .Y(n1238) );
  MXI4X1 U2444 ( .A(\register[4][12] ), .B(\register[5][12] ), .C(
        \register[6][12] ), .D(\register[7][12] ), .S0(n1624), .S1(n1592), .Y(
        n1242) );
  MXI4X1 U2445 ( .A(\register[4][13] ), .B(\register[5][13] ), .C(
        \register[6][13] ), .D(\register[7][13] ), .S0(n1619), .S1(n1594), .Y(
        n1250) );
  MXI4X1 U2446 ( .A(\register[20][13] ), .B(\register[21][13] ), .C(
        \register[22][13] ), .D(\register[23][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1246) );
  MXI4X1 U2447 ( .A(\register[20][15] ), .B(\register[21][15] ), .C(
        \register[22][15] ), .D(\register[23][15] ), .S0(n1620), .S1(n1594), 
        .Y(n1262) );
  MXI4X1 U2448 ( .A(\register[4][15] ), .B(\register[5][15] ), .C(
        \register[6][15] ), .D(\register[7][15] ), .S0(n1625), .S1(n1592), .Y(
        n1266) );
  MXI4X1 U2449 ( .A(\register[4][16] ), .B(\register[5][16] ), .C(
        \register[6][16] ), .D(\register[7][16] ), .S0(n1608), .S1(n1585), .Y(
        n1274) );
  MXI4X1 U2450 ( .A(\register[20][16] ), .B(\register[21][16] ), .C(
        \register[22][16] ), .D(\register[23][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1270) );
  MXI4X1 U2451 ( .A(\register[4][17] ), .B(\register[5][17] ), .C(
        \register[6][17] ), .D(\register[7][17] ), .S0(n1608), .S1(n1585), .Y(
        n1282) );
  MXI4X1 U2452 ( .A(\register[20][17] ), .B(\register[21][17] ), .C(
        \register[22][17] ), .D(\register[23][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1278) );
  MXI4X1 U2453 ( .A(\register[4][18] ), .B(\register[5][18] ), .C(
        \register[6][18] ), .D(\register[7][18] ), .S0(n1609), .S1(n1585), .Y(
        n1290) );
  MXI4X1 U2454 ( .A(\register[20][18] ), .B(\register[21][18] ), .C(
        \register[22][18] ), .D(\register[23][18] ), .S0(n1609), .S1(n1585), 
        .Y(n1286) );
  MXI4X1 U2455 ( .A(\register[4][19] ), .B(\register[5][19] ), .C(
        \register[6][19] ), .D(\register[7][19] ), .S0(n1609), .S1(n1586), .Y(
        n1298) );
  MXI4X1 U2456 ( .A(\register[20][19] ), .B(\register[21][19] ), .C(
        \register[22][19] ), .D(\register[23][19] ), .S0(n1609), .S1(n1586), 
        .Y(n1294) );
  MXI4X1 U2457 ( .A(\register[4][20] ), .B(\register[5][20] ), .C(
        \register[6][20] ), .D(\register[7][20] ), .S0(n1610), .S1(n1586), .Y(
        n1306) );
  MXI4X1 U2458 ( .A(\register[20][20] ), .B(\register[21][20] ), .C(
        \register[22][20] ), .D(\register[23][20] ), .S0(n1610), .S1(n1586), 
        .Y(n1302) );
  MXI4X1 U2459 ( .A(\register[4][21] ), .B(\register[5][21] ), .C(
        \register[6][21] ), .D(\register[7][21] ), .S0(n1610), .S1(n1586), .Y(
        n1314) );
  MXI4X1 U2460 ( .A(\register[20][21] ), .B(\register[21][21] ), .C(
        \register[22][21] ), .D(\register[23][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1310) );
  MXI4X1 U2461 ( .A(\register[4][22] ), .B(\register[5][22] ), .C(
        \register[6][22] ), .D(\register[7][22] ), .S0(n1611), .S1(n1587), .Y(
        n1322) );
  MXI4X1 U2462 ( .A(\register[20][22] ), .B(\register[21][22] ), .C(
        \register[22][22] ), .D(\register[23][22] ), .S0(n1610), .S1(n1587), 
        .Y(n1318) );
  MXI4X1 U2463 ( .A(\register[4][23] ), .B(\register[5][23] ), .C(
        \register[6][23] ), .D(\register[7][23] ), .S0(n1611), .S1(n1587), .Y(
        n1330) );
  MXI4X1 U2464 ( .A(\register[20][23] ), .B(\register[21][23] ), .C(
        \register[22][23] ), .D(\register[23][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1326) );
  MXI4X1 U2465 ( .A(\register[4][24] ), .B(\register[5][24] ), .C(
        \register[6][24] ), .D(\register[7][24] ), .S0(n1612), .S1(n1587), .Y(
        n1338) );
  MXI4X1 U2466 ( .A(\register[20][24] ), .B(\register[21][24] ), .C(
        \register[22][24] ), .D(\register[23][24] ), .S0(n1611), .S1(n1587), 
        .Y(n1334) );
  MXI4X1 U2467 ( .A(\register[4][25] ), .B(\register[5][25] ), .C(
        \register[6][25] ), .D(\register[7][25] ), .S0(n1612), .S1(n1588), .Y(
        n1346) );
  MXI4X1 U2468 ( .A(\register[20][25] ), .B(\register[21][25] ), .C(
        \register[22][25] ), .D(\register[23][25] ), .S0(n1612), .S1(n1588), 
        .Y(n1342) );
  MXI4X1 U2469 ( .A(\register[4][26] ), .B(\register[5][26] ), .C(
        \register[6][26] ), .D(\register[7][26] ), .S0(n1613), .S1(n1588), .Y(
        n1354) );
  MXI4X1 U2470 ( .A(\register[20][26] ), .B(\register[21][26] ), .C(
        \register[22][26] ), .D(\register[23][26] ), .S0(n1612), .S1(n1588), 
        .Y(n1350) );
  MXI4X1 U2471 ( .A(\register[4][27] ), .B(\register[5][27] ), .C(
        \register[6][27] ), .D(\register[7][27] ), .S0(n1613), .S1(n1588), .Y(
        n1362) );
  MXI4X1 U2472 ( .A(\register[20][27] ), .B(\register[21][27] ), .C(
        \register[22][27] ), .D(\register[23][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1358) );
  MXI4X1 U2473 ( .A(\register[4][28] ), .B(\register[5][28] ), .C(
        \register[6][28] ), .D(\register[7][28] ), .S0(n1614), .S1(n1589), .Y(
        n1370) );
  MXI4X1 U2474 ( .A(\register[20][28] ), .B(\register[21][28] ), .C(
        \register[22][28] ), .D(\register[23][28] ), .S0(n1613), .S1(n1588), 
        .Y(n1366) );
  MXI4X1 U2475 ( .A(\register[4][29] ), .B(\register[5][29] ), .C(
        \register[6][29] ), .D(\register[7][29] ), .S0(n1614), .S1(n1589), .Y(
        n1378) );
  MXI4X1 U2476 ( .A(\register[20][29] ), .B(\register[21][29] ), .C(
        \register[22][29] ), .D(\register[23][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1374) );
  MXI4X1 U2477 ( .A(\register[4][30] ), .B(\register[5][30] ), .C(
        \register[6][30] ), .D(\register[7][30] ), .S0(n1615), .S1(n1589), .Y(
        n1386) );
  MXI4X1 U2478 ( .A(\register[20][30] ), .B(\register[21][30] ), .C(
        \register[22][30] ), .D(\register[23][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1382) );
  MXI4X1 U2479 ( .A(\register[4][31] ), .B(\register[5][31] ), .C(
        \register[6][31] ), .D(\register[7][31] ), .S0(n1620), .S1(n1595), .Y(
        n1394) );
  MXI4X1 U2480 ( .A(\register[20][31] ), .B(\register[21][31] ), .C(
        \register[22][31] ), .D(\register[23][31] ), .S0(n1615), .S1(n1589), 
        .Y(n1390) );
  MXI4X1 U2481 ( .A(\register[16][1] ), .B(\register[17][1] ), .C(
        \register[18][1] ), .D(\register[19][1] ), .S0(n2166), .S1(n2141), .Y(
        n1701) );
  MXI4X1 U2482 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n2166), .S1(n2141), .Y(
        n1709) );
  MXI4X1 U2483 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n2167), .S1(n2142), .Y(
        n1717) );
  MXI4X1 U2484 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n2167), .S1(n2142), .Y(
        n1725) );
  MXI4X1 U2485 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n2168), .S1(n2143), .Y(
        n1741) );
  MXI4X1 U2486 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n2171), .S1(n2145), 
        .Y(n1789) );
  MXI4X1 U2487 ( .A(\register[16][14] ), .B(\register[17][14] ), .C(
        \register[18][14] ), .D(\register[19][14] ), .S0(n2172), .S1(n2145), 
        .Y(n1805) );
  MXI4X1 U2488 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n2172), .S1(n2145), 
        .Y(n1813) );
  MXI4X1 U2489 ( .A(\register[16][2] ), .B(\register[17][2] ), .C(
        \register[18][2] ), .D(\register[19][2] ), .S0(n1616), .S1(n1590), .Y(
        n1159) );
  MXI4X1 U2490 ( .A(\register[16][3] ), .B(\register[17][3] ), .C(
        \register[18][3] ), .D(\register[19][3] ), .S0(n1617), .S1(n1591), .Y(
        n1167) );
  MXI4X1 U2491 ( .A(\register[16][4] ), .B(\register[17][4] ), .C(
        \register[18][4] ), .D(\register[19][4] ), .S0(n1617), .S1(n1591), .Y(
        n1175) );
  MXI4X1 U2492 ( .A(\register[16][6] ), .B(\register[17][6] ), .C(
        \register[18][6] ), .D(\register[19][6] ), .S0(n1625), .S1(n1592), .Y(
        n1191) );
  MXI4X1 U2493 ( .A(\register[16][8] ), .B(\register[17][8] ), .C(
        \register[18][8] ), .D(\register[19][8] ), .S0(n1625), .S1(n1592), .Y(
        n1207) );
  MXI4X1 U2494 ( .A(\register[16][12] ), .B(\register[17][12] ), .C(
        \register[18][12] ), .D(\register[19][12] ), .S0(n1619), .S1(n1594), 
        .Y(n1239) );
  MXI4X1 U2495 ( .A(\register[16][15] ), .B(\register[17][15] ), .C(
        \register[18][15] ), .D(\register[19][15] ), .S0(n1620), .S1(n1594), 
        .Y(n1263) );
  MXI4X1 U2496 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n2165), .S1(n2141), .Y(
        n1694) );
  MXI4X1 U2497 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n2165), .S1(n2141), .Y(
        n1690) );
  MXI4X1 U2498 ( .A(\register[28][1] ), .B(\register[29][1] ), .C(
        \register[30][1] ), .D(\register[31][1] ), .S0(n2165), .S1(n2141), .Y(
        n1698) );
  MXI4X1 U2499 ( .A(\register[12][1] ), .B(\register[13][1] ), .C(
        \register[14][1] ), .D(\register[15][1] ), .S0(n2166), .S1(n2141), .Y(
        n1702) );
  MXI4X1 U2500 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n2166), .S1(n2141), .Y(
        n1706) );
  MXI4X1 U2501 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n2166), .S1(n2141), .Y(
        n1710) );
  MXI4X1 U2502 ( .A(\register[28][3] ), .B(\register[29][3] ), .C(
        \register[30][3] ), .D(\register[31][3] ), .S0(n2166), .S1(n2142), .Y(
        n1714) );
  MXI4X1 U2503 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n2167), .S1(n2142), .Y(
        n1718) );
  MXI4X1 U2504 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n2167), .S1(n2142), .Y(
        n1722) );
  MXI4X1 U2505 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n2167), .S1(n2142), .Y(
        n1726) );
  MXI4X1 U2506 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n2168), .S1(n2142), .Y(
        n1734) );
  MXI4X1 U2507 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n2167), .S1(n2142), .Y(
        n1730) );
  MXI4X1 U2508 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n2168), .S1(n2142), .Y(
        n1738) );
  MXI4X1 U2509 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n2168), .S1(n2143), .Y(
        n1742) );
  MXI4X1 U2510 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n2169), .S1(n2143), .Y(
        n1758) );
  MXI4X1 U2511 ( .A(\register[12][9] ), .B(\register[13][9] ), .C(
        \register[14][9] ), .D(\register[15][9] ), .S0(n2169), .S1(n2144), .Y(
        n1766) );
  MXI4X1 U2512 ( .A(\register[28][9] ), .B(\register[29][9] ), .C(
        \register[30][9] ), .D(\register[31][9] ), .S0(n2169), .S1(n2143), .Y(
        n1762) );
  MXI4X1 U2513 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1774) );
  MXI4X1 U2514 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1770) );
  MXI4X1 U2515 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1782) );
  MXI4X1 U2516 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1778) );
  MXI4X1 U2517 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n2171), .S1(n2144), 
        .Y(n1786) );
  MXI4X1 U2518 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n2171), .S1(n2145), 
        .Y(n1790) );
  MXI4X1 U2519 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1798) );
  MXI4X1 U2520 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1794) );
  MXI4X1 U2521 ( .A(\register[28][14] ), .B(\register[29][14] ), .C(
        \register[30][14] ), .D(\register[31][14] ), .S0(n2171), .S1(n2145), 
        .Y(n1802) );
  MXI4X1 U2522 ( .A(\register[12][14] ), .B(\register[13][14] ), .C(
        \register[14][14] ), .D(\register[15][14] ), .S0(n2172), .S1(n2145), 
        .Y(n1806) );
  MXI4X1 U2523 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n2172), .S1(n2145), 
        .Y(n1810) );
  MXI4X1 U2524 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1822) );
  MXI4X1 U2525 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1818) );
  MXI4X1 U2526 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1830) );
  MXI4X1 U2527 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1826) );
  MXI4X1 U2528 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n2159), .S1(n2136), 
        .Y(n1838) );
  MXI4X1 U2529 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n2158), .S1(n2136), 
        .Y(n1834) );
  MXI4X1 U2530 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n2159), .S1(n2137), 
        .Y(n1846) );
  MXI4X1 U2531 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n2159), .S1(n2136), 
        .Y(n1842) );
  MXI4X1 U2532 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1862) );
  MXI4X1 U2533 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1858) );
  MXI4X1 U2534 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n2161), .S1(n2138), 
        .Y(n1870) );
  MXI4X1 U2535 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n2160), .S1(n2137), 
        .Y(n1866) );
  MXI4X1 U2536 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1878) );
  MXI4X1 U2537 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1874) );
  MXI4X1 U2538 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n2162), .S1(n2138), 
        .Y(n1886) );
  MXI4X1 U2539 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n2161), .S1(n2138), 
        .Y(n1882) );
  MXI4X1 U2540 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n2162), .S1(n2139), 
        .Y(n1894) );
  MXI4X1 U2541 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n2162), .S1(n2138), 
        .Y(n1890) );
  MXI4X1 U2542 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n2163), .S1(n2139), 
        .Y(n1902) );
  MXI4X1 U2543 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n2162), .S1(n2139), 
        .Y(n1898) );
  MXI4X1 U2544 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1910) );
  MXI4X1 U2545 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1906) );
  MXI4X1 U2546 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n2163), .S1(n2140), 
        .Y(n1918) );
  MXI4X1 U2547 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n2163), .S1(n2139), 
        .Y(n1914) );
  MXI4X1 U2548 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1926) );
  MXI4X1 U2549 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1922) );
  MXI4X1 U2550 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1934) );
  MXI4X1 U2551 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1930) );
  MXI4X1 U2552 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n2165), .S1(n2141), 
        .Y(n1942) );
  MXI4X1 U2553 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n2165), .S1(n2140), 
        .Y(n1938) );
  MXI4X1 U2554 ( .A(\register[12][0] ), .B(\register[13][0] ), .C(
        \register[14][0] ), .D(\register[15][0] ), .S0(n1615), .S1(n1590), .Y(
        n1144) );
  MXI4X1 U2555 ( .A(\register[28][0] ), .B(\register[29][0] ), .C(
        \register[30][0] ), .D(\register[31][0] ), .S0(n1615), .S1(n1590), .Y(
        n1140) );
  MXI4X1 U2556 ( .A(\register[28][2] ), .B(\register[29][2] ), .C(
        \register[30][2] ), .D(\register[31][2] ), .S0(n1616), .S1(n1590), .Y(
        n1156) );
  MXI4X1 U2557 ( .A(\register[12][2] ), .B(\register[13][2] ), .C(
        \register[14][2] ), .D(\register[15][2] ), .S0(n1616), .S1(n1590), .Y(
        n1160) );
  MXI4X1 U2558 ( .A(\register[12][3] ), .B(\register[13][3] ), .C(
        \register[14][3] ), .D(\register[15][3] ), .S0(n1617), .S1(n1591), .Y(
        n1168) );
  MXI4X1 U2559 ( .A(\register[28][4] ), .B(\register[29][4] ), .C(
        \register[30][4] ), .D(\register[31][4] ), .S0(n1617), .S1(n1591), .Y(
        n1172) );
  MXI4X1 U2560 ( .A(\register[12][4] ), .B(\register[13][4] ), .C(
        \register[14][4] ), .D(\register[15][4] ), .S0(n1617), .S1(n1591), .Y(
        n1176) );
  MXI4X1 U2561 ( .A(\register[12][5] ), .B(\register[13][5] ), .C(
        \register[14][5] ), .D(\register[15][5] ), .S0(n1624), .S1(n1591), .Y(
        n1184) );
  MXI4X1 U2562 ( .A(\register[28][5] ), .B(\register[29][5] ), .C(
        \register[30][5] ), .D(\register[31][5] ), .S0(n1617), .S1(n1591), .Y(
        n1180) );
  MXI4X1 U2563 ( .A(\register[28][6] ), .B(\register[29][6] ), .C(
        \register[30][6] ), .D(\register[31][6] ), .S0(n1624), .S1(n1591), .Y(
        n1188) );
  MXI4X1 U2564 ( .A(\register[12][6] ), .B(\register[13][6] ), .C(
        \register[14][6] ), .D(\register[15][6] ), .S0(n1624), .S1(n1592), .Y(
        n1192) );
  MXI4X1 U2565 ( .A(\register[12][7] ), .B(\register[13][7] ), .C(
        \register[14][7] ), .D(\register[15][7] ), .S0(n1624), .S1(n1592), .Y(
        n1200) );
  MXI4X1 U2566 ( .A(\register[28][7] ), .B(\register[29][7] ), .C(
        \register[30][7] ), .D(\register[31][7] ), .S0(n1624), .S1(n1592), .Y(
        n1196) );
  MXI4X1 U2567 ( .A(\register[28][8] ), .B(\register[29][8] ), .C(
        \register[30][8] ), .D(\register[31][8] ), .S0(n1620), .S1(n1595), .Y(
        n1204) );
  MXI4X1 U2568 ( .A(\register[12][8] ), .B(\register[13][8] ), .C(
        \register[14][8] ), .D(\register[15][8] ), .S0(n1624), .S1(n1592), .Y(
        n1208) );
  MXI4X1 U2569 ( .A(\register[12][10] ), .B(\register[13][10] ), .C(
        \register[14][10] ), .D(\register[15][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1224) );
  MXI4X1 U2570 ( .A(\register[28][10] ), .B(\register[29][10] ), .C(
        \register[30][10] ), .D(\register[31][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1220) );
  MXI4X1 U2571 ( .A(\register[12][11] ), .B(\register[13][11] ), .C(
        \register[14][11] ), .D(\register[15][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1232) );
  MXI4X1 U2572 ( .A(\register[28][11] ), .B(\register[29][11] ), .C(
        \register[30][11] ), .D(\register[31][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1228) );
  MXI4X1 U2573 ( .A(\register[28][12] ), .B(\register[29][12] ), .C(
        \register[30][12] ), .D(\register[31][12] ), .S0(n1619), .S1(n1593), 
        .Y(n1236) );
  MXI4X1 U2574 ( .A(\register[12][12] ), .B(\register[13][12] ), .C(
        \register[14][12] ), .D(\register[15][12] ), .S0(n1619), .S1(n1594), 
        .Y(n1240) );
  MXI4X1 U2575 ( .A(\register[12][13] ), .B(\register[13][13] ), .C(
        \register[14][13] ), .D(\register[15][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1248) );
  MXI4X1 U2576 ( .A(\register[28][13] ), .B(\register[29][13] ), .C(
        \register[30][13] ), .D(\register[31][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1244) );
  MXI4X1 U2577 ( .A(\register[28][15] ), .B(\register[29][15] ), .C(
        \register[30][15] ), .D(\register[31][15] ), .S0(n1620), .S1(n1594), 
        .Y(n1260) );
  MXI4X1 U2578 ( .A(\register[12][15] ), .B(\register[13][15] ), .C(
        \register[14][15] ), .D(\register[15][15] ), .S0(n1620), .S1(n1595), 
        .Y(n1264) );
  MXI4X1 U2579 ( .A(\register[12][16] ), .B(\register[13][16] ), .C(
        \register[14][16] ), .D(\register[15][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1272) );
  MXI4X1 U2580 ( .A(\register[28][16] ), .B(\register[29][16] ), .C(
        \register[30][16] ), .D(\register[31][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1268) );
  MXI4X1 U2581 ( .A(\register[12][17] ), .B(\register[13][17] ), .C(
        \register[14][17] ), .D(\register[15][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1280) );
  MXI4X1 U2582 ( .A(\register[28][17] ), .B(\register[29][17] ), .C(
        \register[30][17] ), .D(\register[31][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1276) );
  MXI4X1 U2583 ( .A(\register[12][18] ), .B(\register[13][18] ), .C(
        \register[14][18] ), .D(\register[15][18] ), .S0(n1609), .S1(n1585), 
        .Y(n1288) );
  MXI4X1 U2584 ( .A(\register[28][18] ), .B(\register[29][18] ), .C(
        \register[30][18] ), .D(\register[31][18] ), .S0(n1608), .S1(n1585), 
        .Y(n1284) );
  MXI4X1 U2585 ( .A(\register[12][19] ), .B(\register[13][19] ), .C(
        \register[14][19] ), .D(\register[15][19] ), .S0(n1609), .S1(n1586), 
        .Y(n1296) );
  MXI4X1 U2586 ( .A(\register[28][19] ), .B(\register[29][19] ), .C(
        \register[30][19] ), .D(\register[31][19] ), .S0(n1609), .S1(n1585), 
        .Y(n1292) );
  MXI4X1 U2587 ( .A(\register[12][20] ), .B(\register[13][20] ), .C(
        \register[14][20] ), .D(\register[15][20] ), .S0(n1610), .S1(n1586), 
        .Y(n1304) );
  MXI4X1 U2588 ( .A(\register[28][20] ), .B(\register[29][20] ), .C(
        \register[30][20] ), .D(\register[31][20] ), .S0(n1609), .S1(n1586), 
        .Y(n1300) );
  MXI4X1 U2589 ( .A(\register[12][21] ), .B(\register[13][21] ), .C(
        \register[14][21] ), .D(\register[15][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1312) );
  MXI4X1 U2590 ( .A(\register[28][21] ), .B(\register[29][21] ), .C(
        \register[30][21] ), .D(\register[31][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1308) );
  MXI4X1 U2591 ( .A(\register[12][22] ), .B(\register[13][22] ), .C(
        \register[14][22] ), .D(\register[15][22] ), .S0(n1611), .S1(n1587), 
        .Y(n1320) );
  MXI4X1 U2592 ( .A(\register[28][22] ), .B(\register[29][22] ), .C(
        \register[30][22] ), .D(\register[31][22] ), .S0(n1610), .S1(n1586), 
        .Y(n1316) );
  MXI4X1 U2593 ( .A(\register[12][23] ), .B(\register[13][23] ), .C(
        \register[14][23] ), .D(\register[15][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1328) );
  MXI4X1 U2594 ( .A(\register[28][23] ), .B(\register[29][23] ), .C(
        \register[30][23] ), .D(\register[31][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1324) );
  MXI4X1 U2595 ( .A(\register[12][24] ), .B(\register[13][24] ), .C(
        \register[14][24] ), .D(\register[15][24] ), .S0(n1612), .S1(n1587), 
        .Y(n1336) );
  MXI4X1 U2596 ( .A(\register[28][24] ), .B(\register[29][24] ), .C(
        \register[30][24] ), .D(\register[31][24] ), .S0(n1611), .S1(n1587), 
        .Y(n1332) );
  MXI4X1 U2597 ( .A(\register[12][25] ), .B(\register[13][25] ), .C(
        \register[14][25] ), .D(\register[15][25] ), .S0(n1612), .S1(n1588), 
        .Y(n1344) );
  MXI4X1 U2598 ( .A(\register[28][25] ), .B(\register[29][25] ), .C(
        \register[30][25] ), .D(\register[31][25] ), .S0(n1612), .S1(n1587), 
        .Y(n1340) );
  MXI4X1 U2599 ( .A(\register[12][26] ), .B(\register[13][26] ), .C(
        \register[14][26] ), .D(\register[15][26] ), .S0(n1613), .S1(n1588), 
        .Y(n1352) );
  MXI4X1 U2600 ( .A(\register[28][26] ), .B(\register[29][26] ), .C(
        \register[30][26] ), .D(\register[31][26] ), .S0(n1612), .S1(n1588), 
        .Y(n1348) );
  MXI4X1 U2601 ( .A(\register[12][27] ), .B(\register[13][27] ), .C(
        \register[14][27] ), .D(\register[15][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1360) );
  MXI4X1 U2602 ( .A(\register[28][27] ), .B(\register[29][27] ), .C(
        \register[30][27] ), .D(\register[31][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1356) );
  MXI4X1 U2603 ( .A(\register[12][28] ), .B(\register[13][28] ), .C(
        \register[14][28] ), .D(\register[15][28] ), .S0(n1613), .S1(n1589), 
        .Y(n1368) );
  MXI4X1 U2604 ( .A(\register[28][28] ), .B(\register[29][28] ), .C(
        \register[30][28] ), .D(\register[31][28] ), .S0(n1613), .S1(n1588), 
        .Y(n1364) );
  MXI4X1 U2605 ( .A(\register[12][29] ), .B(\register[13][29] ), .C(
        \register[14][29] ), .D(\register[15][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1376) );
  MXI4X1 U2606 ( .A(\register[28][29] ), .B(\register[29][29] ), .C(
        \register[30][29] ), .D(\register[31][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1372) );
  MXI4X1 U2607 ( .A(\register[12][30] ), .B(\register[13][30] ), .C(
        \register[14][30] ), .D(\register[15][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1384) );
  MXI4X1 U2608 ( .A(\register[28][30] ), .B(\register[29][30] ), .C(
        \register[30][30] ), .D(\register[31][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1380) );
  MXI4X1 U2609 ( .A(\register[12][31] ), .B(\register[13][31] ), .C(
        \register[14][31] ), .D(\register[15][31] ), .S0(n1615), .S1(n1590), 
        .Y(n1392) );
  MXI4X1 U2610 ( .A(\register[28][31] ), .B(\register[29][31] ), .C(
        \register[30][31] ), .D(\register[31][31] ), .S0(n1615), .S1(n1589), 
        .Y(n1388) );
  MXI4X1 U2611 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n2165), .S1(n2141), .Y(
        n1695) );
  MXI4X1 U2612 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n2165), .S1(n2141), .Y(
        n1691) );
  MXI4X1 U2613 ( .A(\register[24][1] ), .B(\register[25][1] ), .C(
        \register[26][1] ), .D(\register[27][1] ), .S0(n2165), .S1(n2141), .Y(
        n1699) );
  MXI4X1 U2614 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n2166), .S1(n2141), .Y(
        n1707) );
  MXI4X1 U2615 ( .A(\register[24][3] ), .B(\register[25][3] ), .C(
        \register[26][3] ), .D(\register[27][3] ), .S0(n2166), .S1(n2142), .Y(
        n1715) );
  MXI4X1 U2616 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n2167), .S1(n2142), .Y(
        n1723) );
  MXI4X1 U2617 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n2168), .S1(n2142), .Y(
        n1735) );
  MXI4X1 U2618 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n2167), .S1(n2142), .Y(
        n1731) );
  MXI4X1 U2619 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n2168), .S1(n2143), .Y(
        n1739) );
  MXI4X1 U2620 ( .A(\register[8][8] ), .B(\register[9][8] ), .C(
        \register[10][8] ), .D(\register[11][8] ), .S0(n2169), .S1(n2143), .Y(
        n1759) );
  MXI4X1 U2621 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n2169), .S1(n2143), .Y(
        n1755) );
  MXI4X1 U2622 ( .A(\register[8][9] ), .B(\register[9][9] ), .C(
        \register[10][9] ), .D(\register[11][9] ), .S0(n2170), .S1(n2144), .Y(
        n1767) );
  MXI4X1 U2623 ( .A(\register[24][9] ), .B(\register[25][9] ), .C(
        \register[26][9] ), .D(\register[27][9] ), .S0(n2169), .S1(n2144), .Y(
        n1763) );
  MXI4X1 U2624 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1775) );
  MXI4X1 U2625 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n2170), .S1(n2144), 
        .Y(n1771) );
  MXI4X1 U2626 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1783) );
  MXI4X1 U2627 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n2170), .S1(n2144), 
        .Y(n1779) );
  MXI4X1 U2628 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n2171), .S1(n2144), 
        .Y(n1787) );
  MXI4X1 U2629 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1799) );
  MXI4X1 U2630 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n2171), .S1(n2145), 
        .Y(n1795) );
  MXI4X1 U2631 ( .A(\register[24][14] ), .B(\register[25][14] ), .C(
        \register[26][14] ), .D(\register[27][14] ), .S0(n2172), .S1(n2145), 
        .Y(n1803) );
  MXI4X1 U2632 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n2172), .S1(n2145), 
        .Y(n1811) );
  MXI4X1 U2633 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1823) );
  MXI4X1 U2634 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n2158), .S1(n2136), 
        .Y(n1819) );
  MXI4X1 U2635 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1831) );
  MXI4X1 U2636 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n2158), .S1(n2136), 
        .Y(n1827) );
  MXI4X1 U2637 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n2159), .S1(n2136), 
        .Y(n1839) );
  MXI4X1 U2638 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n2159), .S1(n2136), 
        .Y(n1835) );
  MXI4X1 U2639 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n2159), .S1(n2137), 
        .Y(n1847) );
  MXI4X1 U2640 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n2159), .S1(n2137), 
        .Y(n1843) );
  MXI4X1 U2641 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1863) );
  MXI4X1 U2642 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n2160), .S1(n2137), 
        .Y(n1859) );
  MXI4X1 U2643 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n2161), .S1(n2138), 
        .Y(n1871) );
  MXI4X1 U2644 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n2160), .S1(n2137), 
        .Y(n1867) );
  MXI4X1 U2645 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1879) );
  MXI4X1 U2646 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n2161), .S1(n2138), 
        .Y(n1875) );
  MXI4X1 U2647 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n2162), .S1(n2138), 
        .Y(n1887) );
  MXI4X1 U2648 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n2161), .S1(n2138), 
        .Y(n1883) );
  MXI4X1 U2649 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n2162), .S1(n2139), 
        .Y(n1895) );
  MXI4X1 U2650 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n2162), .S1(n2138), 
        .Y(n1891) );
  MXI4X1 U2651 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n2163), .S1(n2139), 
        .Y(n1903) );
  MXI4X1 U2652 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n2162), .S1(n2139), 
        .Y(n1899) );
  MXI4X1 U2653 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1911) );
  MXI4X1 U2654 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n2163), .S1(n2139), 
        .Y(n1907) );
  MXI4X1 U2655 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n2164), .S1(n2140), 
        .Y(n1919) );
  MXI4X1 U2656 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n2163), .S1(n2139), 
        .Y(n1915) );
  MXI4X1 U2657 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1927) );
  MXI4X1 U2658 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n2164), .S1(n2140), 
        .Y(n1923) );
  MXI4X1 U2659 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1935) );
  MXI4X1 U2660 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n2164), .S1(n2140), 
        .Y(n1931) );
  MXI4X1 U2661 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n2161), .S1(n2138), 
        .Y(n1943) );
  MXI4X1 U2662 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n2165), .S1(n2140), 
        .Y(n1939) );
  MXI4X1 U2663 ( .A(\register[8][0] ), .B(\register[9][0] ), .C(
        \register[10][0] ), .D(\register[11][0] ), .S0(n1615), .S1(n1590), .Y(
        n1145) );
  MXI4X1 U2664 ( .A(\register[24][0] ), .B(\register[25][0] ), .C(
        \register[26][0] ), .D(\register[27][0] ), .S0(n1615), .S1(n1590), .Y(
        n1141) );
  MXI4X1 U2665 ( .A(\register[24][2] ), .B(\register[25][2] ), .C(
        \register[26][2] ), .D(\register[27][2] ), .S0(n1616), .S1(n1590), .Y(
        n1157) );
  MXI4X1 U2666 ( .A(\register[24][4] ), .B(\register[25][4] ), .C(
        \register[26][4] ), .D(\register[27][4] ), .S0(n1617), .S1(n1591), .Y(
        n1173) );
  MXI4X1 U2667 ( .A(\register[8][5] ), .B(\register[9][5] ), .C(
        \register[10][5] ), .D(\register[11][5] ), .S0(n1605), .S1(n1591), .Y(
        n1185) );
  MXI4X1 U2668 ( .A(\register[24][5] ), .B(\register[25][5] ), .C(
        \register[26][5] ), .D(\register[27][5] ), .S0(n1617), .S1(n1591), .Y(
        n1181) );
  MXI4X1 U2669 ( .A(\register[24][6] ), .B(\register[25][6] ), .C(
        \register[26][6] ), .D(\register[27][6] ), .S0(n1624), .S1(n1592), .Y(
        n1189) );
  MXI4X1 U2670 ( .A(\register[24][7] ), .B(\register[25][7] ), .C(
        \register[26][7] ), .D(\register[27][7] ), .S0(n1624), .S1(n1592), .Y(
        n1197) );
  MXI4X1 U2671 ( .A(\register[24][8] ), .B(\register[25][8] ), .C(
        \register[26][8] ), .D(\register[27][8] ), .S0(n1624), .S1(n1592), .Y(
        n1205) );
  MXI4X1 U2672 ( .A(\register[8][10] ), .B(\register[9][10] ), .C(
        \register[10][10] ), .D(\register[11][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1225) );
  MXI4X1 U2673 ( .A(\register[24][10] ), .B(\register[25][10] ), .C(
        \register[26][10] ), .D(\register[27][10] ), .S0(n1618), .S1(n1593), 
        .Y(n1221) );
  MXI4X1 U2674 ( .A(\register[8][11] ), .B(\register[9][11] ), .C(
        \register[10][11] ), .D(\register[11][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1233) );
  MXI4X1 U2675 ( .A(\register[24][11] ), .B(\register[25][11] ), .C(
        \register[26][11] ), .D(\register[27][11] ), .S0(n1618), .S1(n1593), 
        .Y(n1229) );
  MXI4X1 U2676 ( .A(\register[24][12] ), .B(\register[25][12] ), .C(
        \register[26][12] ), .D(\register[27][12] ), .S0(n1619), .S1(n1593), 
        .Y(n1237) );
  MXI4X1 U2677 ( .A(\register[8][13] ), .B(\register[9][13] ), .C(
        \register[10][13] ), .D(\register[11][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1249) );
  MXI4X1 U2678 ( .A(\register[24][13] ), .B(\register[25][13] ), .C(
        \register[26][13] ), .D(\register[27][13] ), .S0(n1619), .S1(n1594), 
        .Y(n1245) );
  MXI4X1 U2679 ( .A(\register[24][15] ), .B(\register[25][15] ), .C(
        \register[26][15] ), .D(\register[27][15] ), .S0(n1620), .S1(n1594), 
        .Y(n1261) );
  MXI4X1 U2680 ( .A(\register[8][16] ), .B(\register[9][16] ), .C(
        \register[10][16] ), .D(\register[11][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1273) );
  MXI4X1 U2681 ( .A(\register[24][16] ), .B(\register[25][16] ), .C(
        \register[26][16] ), .D(\register[27][16] ), .S0(n1608), .S1(n1585), 
        .Y(n1269) );
  MXI4X1 U2682 ( .A(\register[8][17] ), .B(\register[9][17] ), .C(
        \register[10][17] ), .D(\register[11][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1281) );
  MXI4X1 U2683 ( .A(\register[24][17] ), .B(\register[25][17] ), .C(
        \register[26][17] ), .D(\register[27][17] ), .S0(n1608), .S1(n1585), 
        .Y(n1277) );
  MXI4X1 U2684 ( .A(\register[8][18] ), .B(\register[9][18] ), .C(
        \register[10][18] ), .D(\register[11][18] ), .S0(n1609), .S1(n1585), 
        .Y(n1289) );
  MXI4X1 U2685 ( .A(\register[24][18] ), .B(\register[25][18] ), .C(
        \register[26][18] ), .D(\register[27][18] ), .S0(n1609), .S1(n1585), 
        .Y(n1285) );
  MXI4X1 U2686 ( .A(\register[8][19] ), .B(\register[9][19] ), .C(
        \register[10][19] ), .D(\register[11][19] ), .S0(n1609), .S1(n1586), 
        .Y(n1297) );
  MXI4X1 U2687 ( .A(\register[24][19] ), .B(\register[25][19] ), .C(
        \register[26][19] ), .D(\register[27][19] ), .S0(n1609), .S1(n1586), 
        .Y(n1293) );
  MXI4X1 U2688 ( .A(\register[8][20] ), .B(\register[9][20] ), .C(
        \register[10][20] ), .D(\register[11][20] ), .S0(n1610), .S1(n1586), 
        .Y(n1305) );
  MXI4X1 U2689 ( .A(\register[24][20] ), .B(\register[25][20] ), .C(
        \register[26][20] ), .D(\register[27][20] ), .S0(n1609), .S1(n1586), 
        .Y(n1301) );
  MXI4X1 U2690 ( .A(\register[8][21] ), .B(\register[9][21] ), .C(
        \register[10][21] ), .D(\register[11][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1313) );
  MXI4X1 U2691 ( .A(\register[24][21] ), .B(\register[25][21] ), .C(
        \register[26][21] ), .D(\register[27][21] ), .S0(n1610), .S1(n1586), 
        .Y(n1309) );
  MXI4X1 U2692 ( .A(\register[8][22] ), .B(\register[9][22] ), .C(
        \register[10][22] ), .D(\register[11][22] ), .S0(n1611), .S1(n1587), 
        .Y(n1321) );
  MXI4X1 U2693 ( .A(\register[24][22] ), .B(\register[25][22] ), .C(
        \register[26][22] ), .D(\register[27][22] ), .S0(n1610), .S1(n1586), 
        .Y(n1317) );
  MXI4X1 U2694 ( .A(\register[8][23] ), .B(\register[9][23] ), .C(
        \register[10][23] ), .D(\register[11][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1329) );
  MXI4X1 U2695 ( .A(\register[24][23] ), .B(\register[25][23] ), .C(
        \register[26][23] ), .D(\register[27][23] ), .S0(n1611), .S1(n1587), 
        .Y(n1325) );
  MXI4X1 U2696 ( .A(\register[8][24] ), .B(\register[9][24] ), .C(
        \register[10][24] ), .D(\register[11][24] ), .S0(n1612), .S1(n1587), 
        .Y(n1337) );
  MXI4X1 U2697 ( .A(\register[24][24] ), .B(\register[25][24] ), .C(
        \register[26][24] ), .D(\register[27][24] ), .S0(n1611), .S1(n1587), 
        .Y(n1333) );
  MXI4X1 U2698 ( .A(\register[8][25] ), .B(\register[9][25] ), .C(
        \register[10][25] ), .D(\register[11][25] ), .S0(n1612), .S1(n1588), 
        .Y(n1345) );
  MXI4X1 U2699 ( .A(\register[24][25] ), .B(\register[25][25] ), .C(
        \register[26][25] ), .D(\register[27][25] ), .S0(n1612), .S1(n1587), 
        .Y(n1341) );
  MXI4X1 U2700 ( .A(\register[8][26] ), .B(\register[9][26] ), .C(
        \register[10][26] ), .D(\register[11][26] ), .S0(n1613), .S1(n1588), 
        .Y(n1353) );
  MXI4X1 U2701 ( .A(\register[24][26] ), .B(\register[25][26] ), .C(
        \register[26][26] ), .D(\register[27][26] ), .S0(n1612), .S1(n1588), 
        .Y(n1349) );
  MXI4X1 U2702 ( .A(\register[8][27] ), .B(\register[9][27] ), .C(
        \register[10][27] ), .D(\register[11][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1361) );
  MXI4X1 U2703 ( .A(\register[24][27] ), .B(\register[25][27] ), .C(
        \register[26][27] ), .D(\register[27][27] ), .S0(n1613), .S1(n1588), 
        .Y(n1357) );
  MXI4X1 U2704 ( .A(\register[8][28] ), .B(\register[9][28] ), .C(
        \register[10][28] ), .D(\register[11][28] ), .S0(n1614), .S1(n1589), 
        .Y(n1369) );
  MXI4X1 U2705 ( .A(\register[24][28] ), .B(\register[25][28] ), .C(
        \register[26][28] ), .D(\register[27][28] ), .S0(n1613), .S1(n1588), 
        .Y(n1365) );
  MXI4X1 U2706 ( .A(\register[8][29] ), .B(\register[9][29] ), .C(
        \register[10][29] ), .D(\register[11][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1377) );
  MXI4X1 U2707 ( .A(\register[24][29] ), .B(\register[25][29] ), .C(
        \register[26][29] ), .D(\register[27][29] ), .S0(n1614), .S1(n1589), 
        .Y(n1373) );
  MXI4X1 U2708 ( .A(\register[8][30] ), .B(\register[9][30] ), .C(
        \register[10][30] ), .D(\register[11][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1385) );
  MXI4X1 U2709 ( .A(\register[24][30] ), .B(\register[25][30] ), .C(
        \register[26][30] ), .D(\register[27][30] ), .S0(n1614), .S1(n1589), 
        .Y(n1381) );
  MXI4X1 U2710 ( .A(\register[8][31] ), .B(\register[9][31] ), .C(
        \register[10][31] ), .D(\register[11][31] ), .S0(n1611), .S1(n1587), 
        .Y(n1393) );
  MXI4X1 U2711 ( .A(\register[24][31] ), .B(\register[25][31] ), .C(
        \register[26][31] ), .D(\register[27][31] ), .S0(n1615), .S1(n1589), 
        .Y(n1389) );
  XNOR2XL U2712 ( .A(n2544), .B(wsel[0]), .Y(n49) );
  XNOR2XL U2713 ( .A(n2546), .B(wsel[0]), .Y(n58) );
  NOR3X1 U2714 ( .A(n2619), .B(wsel[1]), .C(n2617), .Y(n75) );
  XNOR2XL U2715 ( .A(n2545), .B(wsel[1]), .Y(n48) );
  XNOR2XL U2716 ( .A(n2547), .B(wsel[1]), .Y(n57) );
  XNOR2XL U2717 ( .A(n2548), .B(wsel[2]), .Y(n59) );
  XNOR2XL U2718 ( .A(N19), .B(wsel[2]), .Y(n50) );
endmodule


module extender ( shamt_i, immed_i, ExtOp_i, ExtOut_o );
  input [4:0] shamt_i;
  input [15:0] immed_i;
  output [31:0] ExtOut_o;
  input ExtOp_i;
  wire   n2, n1, n3, n20;

  CLKAND2X8 U1 ( .A(shamt_i[4]), .B(ExtOp_i), .Y(n1) );
  INVX12 U2 ( .A(n1), .Y(n2) );
  CLKINVX8 U3 ( .A(ExtOp_i), .Y(n20) );
  OAI2BB1X2 U4 ( .A0N(immed_i[15]), .A1N(n20), .B0(n2), .Y(ExtOut_o[30]) );
  INVX1 U5 ( .A(n3), .Y(ExtOut_o[18]) );
  OAI2BB1XL U6 ( .A0N(immed_i[6]), .A1N(n20), .B0(n2), .Y(ExtOut_o[6]) );
  OAI2BB1XL U7 ( .A0N(immed_i[7]), .A1N(n20), .B0(n2), .Y(ExtOut_o[7]) );
  OAI2BB1XL U8 ( .A0N(immed_i[8]), .A1N(n20), .B0(n2), .Y(ExtOut_o[8]) );
  OAI2BB1XL U9 ( .A0N(immed_i[9]), .A1N(n20), .B0(n2), .Y(ExtOut_o[9]) );
  OAI2BB1XL U10 ( .A0N(immed_i[10]), .A1N(n20), .B0(n2), .Y(ExtOut_o[10]) );
  OAI2BB1XL U11 ( .A0N(immed_i[11]), .A1N(n20), .B0(n2), .Y(ExtOut_o[11]) );
  OAI2BB1XL U12 ( .A0N(immed_i[12]), .A1N(n20), .B0(n2), .Y(ExtOut_o[12]) );
  OAI2BB1XL U13 ( .A0N(immed_i[14]), .A1N(n20), .B0(n2), .Y(ExtOut_o[14]) );
  INVXL U14 ( .A(n3), .Y(ExtOut_o[15]) );
  INVXL U15 ( .A(n3), .Y(ExtOut_o[16]) );
  INVXL U16 ( .A(n3), .Y(ExtOut_o[17]) );
  INVXL U17 ( .A(n3), .Y(ExtOut_o[19]) );
  INVXL U18 ( .A(n3), .Y(ExtOut_o[20]) );
  OAI2BB1XL U19 ( .A0N(immed_i[4]), .A1N(n20), .B0(n2), .Y(ExtOut_o[4]) );
  OAI2BB1XL U20 ( .A0N(immed_i[5]), .A1N(n20), .B0(n2), .Y(ExtOut_o[5]) );
  OAI2BB1XL U21 ( .A0N(immed_i[13]), .A1N(n20), .B0(n2), .Y(ExtOut_o[13]) );
  INVX3 U22 ( .A(ExtOut_o[30]), .Y(n3) );
  AO22X1 U23 ( .A0(shamt_i[0]), .A1(ExtOp_i), .B0(immed_i[0]), .B1(n20), .Y(
        ExtOut_o[0]) );
  AO22X1 U24 ( .A0(shamt_i[1]), .A1(ExtOp_i), .B0(immed_i[1]), .B1(n20), .Y(
        ExtOut_o[1]) );
  AO22X1 U25 ( .A0(shamt_i[2]), .A1(ExtOp_i), .B0(immed_i[2]), .B1(n20), .Y(
        ExtOut_o[2]) );
  AO22X1 U26 ( .A0(shamt_i[3]), .A1(ExtOp_i), .B0(immed_i[3]), .B1(n20), .Y(
        ExtOut_o[3]) );
  INVXL U27 ( .A(n3), .Y(ExtOut_o[21]) );
  INVXL U28 ( .A(n3), .Y(ExtOut_o[22]) );
  INVXL U29 ( .A(n3), .Y(ExtOut_o[23]) );
  INVXL U30 ( .A(n3), .Y(ExtOut_o[24]) );
  INVXL U31 ( .A(n3), .Y(ExtOut_o[25]) );
  INVXL U32 ( .A(n3), .Y(ExtOut_o[26]) );
  INVXL U33 ( .A(n3), .Y(ExtOut_o[27]) );
  INVXL U34 ( .A(n3), .Y(ExtOut_o[28]) );
  INVXL U35 ( .A(n3), .Y(ExtOut_o[29]) );
  INVXL U36 ( .A(n3), .Y(ExtOut_o[31]) );
endmodule


module MUX_5_3to1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [4:0] data0_i;
  input [4:0] data1_i;
  input [4:0] data2_i;
  input [1:0] select_i;
  output [4:0] data_o;
  wire   n6, n7, n8, n9, n10, n11, n12, n13;

  NOR2BX1 U2 ( .AN(select_i[1]), .B(select_i[0]), .Y(n8) );
  NOR2BX1 U3 ( .AN(select_i[0]), .B(select_i[1]), .Y(n9) );
  NOR2X1 U4 ( .A(select_i[0]), .B(select_i[1]), .Y(n7) );
  CLKINVX1 U5 ( .A(n13), .Y(data_o[0]) );
  AOI222XL U6 ( .A0(data0_i[0]), .A1(n7), .B0(data2_i[0]), .B1(n8), .C0(
        data1_i[0]), .C1(n9), .Y(n13) );
  CLKINVX1 U7 ( .A(n12), .Y(data_o[1]) );
  AOI222XL U8 ( .A0(data0_i[1]), .A1(n7), .B0(data2_i[1]), .B1(n8), .C0(
        data1_i[1]), .C1(n9), .Y(n12) );
  CLKINVX1 U9 ( .A(n11), .Y(data_o[2]) );
  AOI222XL U10 ( .A0(data0_i[2]), .A1(n7), .B0(data2_i[2]), .B1(n8), .C0(
        data1_i[2]), .C1(n9), .Y(n11) );
  CLKINVX1 U11 ( .A(n10), .Y(data_o[3]) );
  AOI222XL U12 ( .A0(data0_i[3]), .A1(n7), .B0(data2_i[3]), .B1(n8), .C0(
        data1_i[3]), .C1(n9), .Y(n10) );
  CLKINVX1 U13 ( .A(n6), .Y(data_o[4]) );
  AOI222XL U14 ( .A0(data0_i[4]), .A1(n7), .B0(data2_i[4]), .B1(n8), .C0(
        data1_i[4]), .C1(n9), .Y(n6) );
endmodule


module MUX_32_3to1_0 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  INVX12 U2 ( .A(select_i[1]), .Y(n32) );
  AO22X4 U3 ( .A0(data2_i[10]), .A1(n4), .B0(data1_i[10]), .B1(n8), .Y(n42) );
  BUFX20 U4 ( .A(n20), .Y(n4) );
  NAND2X2 U5 ( .A(data2_i[0]), .B(n11), .Y(n35) );
  AND2X8 U6 ( .A(n32), .B(n31), .Y(n18) );
  NAND3X6 U7 ( .A(n35), .B(n34), .C(n33), .Y(data_o[0]) );
  BUFX20 U8 ( .A(n20), .Y(n1) );
  AO22X2 U9 ( .A0(data2_i[26]), .A1(n11), .B0(data1_i[26]), .B1(n7), .Y(n48)
         );
  AO22X4 U10 ( .A0(data2_i[12]), .A1(n11), .B0(data1_i[12]), .B1(n7), .Y(n2)
         );
  CLKINVX20 U11 ( .A(n2), .Y(n24) );
  AO22X2 U12 ( .A0(data2_i[1]), .A1(n1), .B0(data1_i[1]), .B1(n8), .Y(n36) );
  AOI22X1 U13 ( .A0(data2_i[11]), .A1(n11), .B0(data1_i[11]), .B1(n7), .Y(n26)
         );
  AO21X4 U14 ( .A0(data0_i[8]), .A1(n10), .B0(n3), .Y(data_o[8]) );
  AO22X4 U15 ( .A0(data2_i[8]), .A1(n11), .B0(data1_i[8]), .B1(n6), .Y(n3) );
  AND2X8 U16 ( .A(select_i[1]), .B(n31), .Y(n20) );
  AO22X4 U17 ( .A0(data2_i[2]), .A1(n1), .B0(data1_i[2]), .B1(n6), .Y(n37) );
  AO22X4 U18 ( .A0(data2_i[13]), .A1(n1), .B0(data1_i[13]), .B1(n6), .Y(n15)
         );
  OAI2BB1X4 U19 ( .A0N(data0_i[29]), .A1N(n10), .B0(n29), .Y(data_o[29]) );
  AOI22X2 U20 ( .A0(data2_i[29]), .A1(n11), .B0(data1_i[29]), .B1(n6), .Y(n29)
         );
  CLKINVX16 U21 ( .A(n19), .Y(n5) );
  INVX16 U22 ( .A(n5), .Y(n6) );
  INVX20 U23 ( .A(n5), .Y(n7) );
  INVX16 U24 ( .A(n5), .Y(n8) );
  AND2X8 U25 ( .A(select_i[0]), .B(n32), .Y(n19) );
  AO22X4 U26 ( .A0(data2_i[4]), .A1(n1), .B0(data1_i[4]), .B1(n7), .Y(n38) );
  AO22X2 U27 ( .A0(data2_i[21]), .A1(n4), .B0(data1_i[21]), .B1(n7), .Y(n46)
         );
  INVX4 U28 ( .A(select_i[0]), .Y(n31) );
  AO22X4 U29 ( .A0(data2_i[6]), .A1(n1), .B0(data1_i[6]), .B1(n7), .Y(n40) );
  AO22X4 U30 ( .A0(data2_i[9]), .A1(n11), .B0(data1_i[9]), .B1(n6), .Y(n41) );
  AO22X2 U31 ( .A0(data2_i[25]), .A1(n4), .B0(data1_i[25]), .B1(n8), .Y(n47)
         );
  AOI22X4 U32 ( .A0(data2_i[3]), .A1(n4), .B0(data1_i[3]), .B1(n8), .Y(n30) );
  AO22X4 U33 ( .A0(data2_i[5]), .A1(n4), .B0(data1_i[5]), .B1(n7), .Y(n39) );
  AO22X2 U34 ( .A0(data2_i[27]), .A1(n4), .B0(data1_i[27]), .B1(n7), .Y(n49)
         );
  OAI2BB1X4 U35 ( .A0N(data0_i[23]), .A1N(n10), .B0(n22), .Y(data_o[23]) );
  AOI22X2 U36 ( .A0(data2_i[23]), .A1(n11), .B0(data1_i[23]), .B1(n6), .Y(n22)
         );
  OAI2BB1X4 U37 ( .A0N(data0_i[11]), .A1N(n10), .B0(n26), .Y(data_o[11]) );
  OAI2BB1X4 U38 ( .A0N(data0_i[24]), .A1N(n10), .B0(n21), .Y(data_o[24]) );
  AOI22X2 U39 ( .A0(data2_i[24]), .A1(n1), .B0(data1_i[24]), .B1(n8), .Y(n21)
         );
  OAI2BB1X4 U40 ( .A0N(data0_i[12]), .A1N(n10), .B0(n24), .Y(data_o[12]) );
  AO22X4 U41 ( .A0(data2_i[20]), .A1(n4), .B0(data1_i[20]), .B1(n7), .Y(n45)
         );
  AO21X4 U42 ( .A0(data0_i[26]), .A1(n10), .B0(n48), .Y(data_o[26]) );
  AOI22X2 U43 ( .A0(data2_i[14]), .A1(n1), .B0(data1_i[14]), .B1(n7), .Y(n23)
         );
  AOI22X1 U44 ( .A0(data2_i[30]), .A1(n1), .B0(data1_i[30]), .B1(n8), .Y(n28)
         );
  AO21X4 U45 ( .A0(data0_i[1]), .A1(n10), .B0(n36), .Y(data_o[1]) );
  AOI22X1 U46 ( .A0(data2_i[22]), .A1(n11), .B0(data1_i[22]), .B1(n6), .Y(n25)
         );
  OAI2BB1X2 U47 ( .A0N(data0_i[30]), .A1N(n10), .B0(n28), .Y(data_o[30]) );
  AOI22X1 U48 ( .A0(data2_i[17]), .A1(n1), .B0(data1_i[17]), .B1(n6), .Y(n27)
         );
  AO21X4 U49 ( .A0(data0_i[13]), .A1(n10), .B0(n15), .Y(data_o[13]) );
  AO21X4 U50 ( .A0(data0_i[2]), .A1(n10), .B0(n37), .Y(data_o[2]) );
  OAI2BB1X2 U51 ( .A0N(data0_i[18]), .A1N(n10), .B0(n13), .Y(data_o[18]) );
  AOI22X2 U52 ( .A0(data2_i[18]), .A1(n11), .B0(data1_i[18]), .B1(n8), .Y(n13)
         );
  AO21X4 U53 ( .A0(data0_i[21]), .A1(n10), .B0(n46), .Y(data_o[21]) );
  AO21X4 U54 ( .A0(data0_i[25]), .A1(n10), .B0(n47), .Y(data_o[25]) );
  OAI2BB1X2 U55 ( .A0N(data0_i[22]), .A1N(n10), .B0(n25), .Y(data_o[22]) );
  AO21X4 U56 ( .A0(data0_i[20]), .A1(n10), .B0(n45), .Y(data_o[20]) );
  AO21X4 U57 ( .A0(data0_i[6]), .A1(n10), .B0(n40), .Y(data_o[6]) );
  AO21X4 U58 ( .A0(data0_i[5]), .A1(n10), .B0(n39), .Y(data_o[5]) );
  AO21X4 U59 ( .A0(data0_i[4]), .A1(n10), .B0(n38), .Y(data_o[4]) );
  AO21X4 U60 ( .A0(data0_i[31]), .A1(n10), .B0(n16), .Y(data_o[31]) );
  AO22X4 U61 ( .A0(data2_i[31]), .A1(n1), .B0(data1_i[31]), .B1(n7), .Y(n16)
         );
  CLKINVX20 U62 ( .A(n9), .Y(n10) );
  INVX16 U63 ( .A(n18), .Y(n9) );
  OAI2BB1X4 U64 ( .A0N(data0_i[3]), .A1N(n10), .B0(n30), .Y(data_o[3]) );
  AO21X4 U65 ( .A0(data0_i[19]), .A1(n10), .B0(n44), .Y(data_o[19]) );
  AO22X4 U66 ( .A0(data2_i[19]), .A1(n1), .B0(data1_i[19]), .B1(n6), .Y(n44)
         );
  AO21X4 U67 ( .A0(data0_i[28]), .A1(n10), .B0(n17), .Y(data_o[28]) );
  AO22X4 U68 ( .A0(data2_i[28]), .A1(n1), .B0(data1_i[28]), .B1(n6), .Y(n17)
         );
  AO21X4 U69 ( .A0(data0_i[7]), .A1(n10), .B0(n14), .Y(data_o[7]) );
  AO22X4 U70 ( .A0(data2_i[7]), .A1(n11), .B0(data1_i[7]), .B1(n8), .Y(n14) );
  AO21X4 U71 ( .A0(data0_i[10]), .A1(n10), .B0(n42), .Y(data_o[10]) );
  BUFX20 U72 ( .A(n20), .Y(n11) );
  NAND2X2 U73 ( .A(data0_i[0]), .B(n10), .Y(n33) );
  AO21X4 U74 ( .A0(data0_i[16]), .A1(n10), .B0(n43), .Y(data_o[16]) );
  AO21X4 U75 ( .A0(data0_i[9]), .A1(n10), .B0(n41), .Y(data_o[9]) );
  AO21X4 U76 ( .A0(data0_i[15]), .A1(n10), .B0(n12), .Y(data_o[15]) );
  OAI2BB1X2 U77 ( .A0N(data0_i[14]), .A1N(n10), .B0(n23), .Y(data_o[14]) );
  AO21X4 U78 ( .A0(data0_i[27]), .A1(n10), .B0(n49), .Y(data_o[27]) );
  AO22X1 U79 ( .A0(data2_i[15]), .A1(n11), .B0(data1_i[15]), .B1(n6), .Y(n12)
         );
  OAI2BB1X2 U80 ( .A0N(data0_i[17]), .A1N(n10), .B0(n27), .Y(data_o[17]) );
  NAND2X2 U81 ( .A(data1_i[0]), .B(n8), .Y(n34) );
  AO22X4 U82 ( .A0(data2_i[16]), .A1(n1), .B0(data1_i[16]), .B1(n8), .Y(n43)
         );
endmodule


module MUX_32_3to1_2 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  AND2X2 U2 ( .A(data2_i[25]), .B(n36), .Y(n39) );
  BUFX20 U3 ( .A(n26), .Y(n5) );
  BUFX4 U4 ( .A(n52), .Y(n9) );
  OR3X6 U5 ( .A(n39), .B(n40), .C(n41), .Y(data_o[25]) );
  OAI2BB1X4 U6 ( .A0N(data0_i[12]), .A1N(n11), .B0(n1), .Y(data_o[12]) );
  AOI22X2 U7 ( .A0(data2_i[12]), .A1(n36), .B0(data1_i[12]), .B1(n24), .Y(n1)
         );
  CLKINVX20 U8 ( .A(n27), .Y(n11) );
  NAND2X2 U9 ( .A(data1_i[30]), .B(n24), .Y(n15) );
  CLKAND2X8 U10 ( .A(data0_i[30]), .B(n28), .Y(n25) );
  NAND2X2 U11 ( .A(data2_i[30]), .B(n36), .Y(n14) );
  OAI2BB2X4 U12 ( .B0(n17), .B1(n13), .A0N(data1_i[8]), .A1N(n24), .Y(n34) );
  CLKINVX1 U13 ( .A(data2_i[8]), .Y(n17) );
  AO21X4 U14 ( .A0(data0_i[8]), .A1(n11), .B0(n34), .Y(data_o[8]) );
  INVX3 U15 ( .A(data2_i[19]), .Y(n23) );
  INVX2 U16 ( .A(data2_i[15]), .Y(n6) );
  INVX6 U17 ( .A(select_i[1]), .Y(n52) );
  INVX12 U18 ( .A(n36), .Y(n13) );
  CLKINVX16 U19 ( .A(n35), .Y(n27) );
  OAI2BB1X4 U20 ( .A0N(data0_i[5]), .A1N(n11), .B0(n2), .Y(data_o[5]) );
  AOI22X2 U21 ( .A0(data2_i[5]), .A1(n36), .B0(data1_i[5]), .B1(n24), .Y(n2)
         );
  CLKAND2X12 U22 ( .A(data0_i[25]), .B(n11), .Y(n41) );
  AOI2BB1X4 U23 ( .A0N(n3), .A1N(n27), .B0(n59), .Y(n4) );
  CLKINVX1 U24 ( .A(data0_i[24]), .Y(n3) );
  INVX6 U25 ( .A(n4), .Y(data_o[24]) );
  CLKAND2X2 U26 ( .A(data1_i[25]), .B(n26), .Y(n40) );
  AOI22X2 U27 ( .A0(data2_i[1]), .A1(n36), .B0(data1_i[1]), .B1(n24), .Y(n50)
         );
  OAI2BB1X4 U28 ( .A0N(data0_i[2]), .A1N(n28), .B0(n48), .Y(data_o[2]) );
  INVX2 U29 ( .A(select_i[0]), .Y(n51) );
  OAI2BB1X4 U30 ( .A0N(data0_i[23]), .A1N(n28), .B0(n45), .Y(data_o[23]) );
  AOI2BB2X4 U31 ( .B0(data1_i[15]), .B1(n5), .A0N(n6), .A1N(n13), .Y(n43) );
  OAI2BB1X4 U32 ( .A0N(data0_i[22]), .A1N(n11), .B0(n44), .Y(data_o[22]) );
  OAI2BB1X4 U33 ( .A0N(data0_i[3]), .A1N(n28), .B0(n7), .Y(data_o[3]) );
  AOI22X2 U34 ( .A0(data2_i[3]), .A1(n36), .B0(data1_i[3]), .B1(n24), .Y(n7)
         );
  OAI2BB1X4 U35 ( .A0N(data0_i[28]), .A1N(n11), .B0(n8), .Y(data_o[28]) );
  AOI22X2 U36 ( .A0(data2_i[28]), .A1(n12), .B0(data1_i[28]), .B1(n26), .Y(n8)
         );
  AOI22X2 U37 ( .A0(data2_i[29]), .A1(n36), .B0(data1_i[29]), .B1(n24), .Y(n42) );
  OAI2BB1X4 U38 ( .A0N(data0_i[11]), .A1N(n28), .B0(n10), .Y(data_o[11]) );
  AOI22X2 U39 ( .A0(data2_i[11]), .A1(n36), .B0(data1_i[11]), .B1(n24), .Y(n10) );
  INVX16 U40 ( .A(n20), .Y(n12) );
  INVX16 U41 ( .A(n20), .Y(n36) );
  AOI2BB2X4 U42 ( .B0(data1_i[19]), .B1(n5), .A0N(n23), .A1N(n13), .Y(n47) );
  OAI2BB1X4 U43 ( .A0N(data0_i[15]), .A1N(n28), .B0(n43), .Y(data_o[15]) );
  CLKINVX8 U44 ( .A(n54), .Y(n19) );
  NAND2X4 U45 ( .A(n14), .B(n15), .Y(n31) );
  AOI22X2 U46 ( .A0(data2_i[27]), .A1(n36), .B0(data1_i[27]), .B1(n24), .Y(n46) );
  CLKAND2X12 U47 ( .A(select_i[0]), .B(n52), .Y(n37) );
  AOI22X4 U48 ( .A0(data2_i[14]), .A1(n36), .B0(data1_i[14]), .B1(n5), .Y(n16)
         );
  AO22X4 U49 ( .A0(data2_i[9]), .A1(n12), .B0(data1_i[9]), .B1(n26), .Y(n33)
         );
  AO22X4 U50 ( .A0(data2_i[31]), .A1(n12), .B0(data1_i[31]), .B1(n26), .Y(n61)
         );
  NAND2X2 U51 ( .A(data0_i[4]), .B(n11), .Y(n18) );
  NAND2X8 U52 ( .A(n18), .B(n19), .Y(data_o[4]) );
  OR2X8 U53 ( .A(select_i[0]), .B(n52), .Y(n20) );
  CLKAND2X12 U54 ( .A(n9), .B(n51), .Y(n35) );
  AOI22X2 U55 ( .A0(data2_i[13]), .A1(n36), .B0(data1_i[13]), .B1(n24), .Y(n49) );
  NAND2X2 U56 ( .A(data0_i[26]), .B(n28), .Y(n21) );
  INVX6 U57 ( .A(n60), .Y(n22) );
  NAND2X8 U58 ( .A(n21), .B(n22), .Y(data_o[26]) );
  OAI2BB1X4 U59 ( .A0N(data0_i[13]), .A1N(n11), .B0(n49), .Y(data_o[13]) );
  OR2X8 U60 ( .A(n25), .B(n31), .Y(data_o[30]) );
  AO22X4 U61 ( .A0(data2_i[21]), .A1(n12), .B0(data1_i[21]), .B1(n26), .Y(n58)
         );
  AO22X4 U62 ( .A0(data2_i[7]), .A1(n12), .B0(data1_i[7]), .B1(n26), .Y(n56)
         );
  OAI2BB1X4 U63 ( .A0N(data0_i[19]), .A1N(n11), .B0(n47), .Y(data_o[19]) );
  AO22X4 U64 ( .A0(data2_i[18]), .A1(n12), .B0(data1_i[18]), .B1(n26), .Y(n30)
         );
  BUFX20 U65 ( .A(n37), .Y(n24) );
  OAI2BB1X4 U66 ( .A0N(data0_i[17]), .A1N(n28), .B0(n38), .Y(data_o[17]) );
  AOI22X2 U67 ( .A0(data2_i[17]), .A1(n36), .B0(data1_i[17]), .B1(n24), .Y(n38) );
  AO22X4 U68 ( .A0(data2_i[16]), .A1(n12), .B0(data1_i[16]), .B1(n26), .Y(n57)
         );
  AO22X4 U69 ( .A0(data2_i[20]), .A1(n12), .B0(data1_i[20]), .B1(n26), .Y(n29)
         );
  AOI22X2 U70 ( .A0(data2_i[2]), .A1(n12), .B0(data1_i[2]), .B1(n24), .Y(n48)
         );
  AOI22X2 U71 ( .A0(data2_i[23]), .A1(n36), .B0(data1_i[23]), .B1(n24), .Y(n45) );
  AO22X4 U72 ( .A0(data2_i[4]), .A1(n36), .B0(data1_i[4]), .B1(n24), .Y(n54)
         );
  AOI22X2 U73 ( .A0(data2_i[22]), .A1(n36), .B0(data1_i[22]), .B1(n24), .Y(n44) );
  AO22X4 U74 ( .A0(data2_i[6]), .A1(n12), .B0(data1_i[6]), .B1(n26), .Y(n55)
         );
  AO22X4 U75 ( .A0(data2_i[10]), .A1(n12), .B0(data1_i[10]), .B1(n26), .Y(n32)
         );
  OAI2BB1X4 U76 ( .A0N(data0_i[29]), .A1N(n28), .B0(n42), .Y(data_o[29]) );
  BUFX20 U77 ( .A(n37), .Y(n26) );
  AO22X4 U78 ( .A0(data2_i[24]), .A1(n12), .B0(data1_i[24]), .B1(n26), .Y(n59)
         );
  AO21X4 U79 ( .A0(data0_i[20]), .A1(n28), .B0(n29), .Y(data_o[20]) );
  AO22X4 U80 ( .A0(data2_i[26]), .A1(n36), .B0(data1_i[26]), .B1(n24), .Y(n60)
         );
  AO22X4 U81 ( .A0(data2_i[0]), .A1(n12), .B0(data1_i[0]), .B1(n26), .Y(n53)
         );
  INVX20 U82 ( .A(n27), .Y(n28) );
  OAI2BB1X4 U83 ( .A0N(data0_i[27]), .A1N(n11), .B0(n46), .Y(data_o[27]) );
  OAI2BB1X4 U84 ( .A0N(data0_i[1]), .A1N(n28), .B0(n50), .Y(data_o[1]) );
  AO21X4 U85 ( .A0(data0_i[18]), .A1(n11), .B0(n30), .Y(data_o[18]) );
  AO21X4 U86 ( .A0(data0_i[10]), .A1(n28), .B0(n32), .Y(data_o[10]) );
  AO21X4 U87 ( .A0(data0_i[9]), .A1(n28), .B0(n33), .Y(data_o[9]) );
  OAI2BB1X4 U88 ( .A0N(data0_i[14]), .A1N(n11), .B0(n16), .Y(data_o[14]) );
  AO21X4 U89 ( .A0(data0_i[0]), .A1(n11), .B0(n53), .Y(data_o[0]) );
  AO21X4 U90 ( .A0(data0_i[6]), .A1(n11), .B0(n55), .Y(data_o[6]) );
  AO21X4 U91 ( .A0(data0_i[7]), .A1(n11), .B0(n56), .Y(data_o[7]) );
  AO21X4 U92 ( .A0(data0_i[16]), .A1(n28), .B0(n57), .Y(data_o[16]) );
  AO21X4 U93 ( .A0(data0_i[21]), .A1(n11), .B0(n58), .Y(data_o[21]) );
  AO21X4 U94 ( .A0(data0_i[31]), .A1(n28), .B0(n61), .Y(data_o[31]) );
endmodule


module MUX_32_3to1_1 ( data0_i, data1_i, data2_i, select_i, data_o );
  input [31:0] data0_i;
  input [31:0] data1_i;
  input [31:0] data2_i;
  input [1:0] select_i;
  output [31:0] data_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  NAND2X6 U2 ( .A(n11), .B(data1_i[0]), .Y(n59) );
  CLKBUFX12 U3 ( .A(n44), .Y(n58) );
  NAND2X6 U4 ( .A(n6), .B(data2_i[1]), .Y(n13) );
  AO22X2 U5 ( .A0(data2_i[30]), .A1(n34), .B0(data1_i[30]), .B1(n35), .Y(n39)
         );
  AND2X4 U6 ( .A(data2_i[8]), .B(n34), .Y(n24) );
  AO22X4 U7 ( .A0(data2_i[28]), .A1(n6), .B0(data1_i[28]), .B1(n35), .Y(n74)
         );
  CLKAND2X8 U8 ( .A(data1_i[16]), .B(n35), .Y(n23) );
  CLKAND2X6 U9 ( .A(data1_i[10]), .B(n35), .Y(n31) );
  CLKAND2X4 U10 ( .A(data1_i[8]), .B(n35), .Y(n25) );
  INVX12 U11 ( .A(n19), .Y(n2) );
  AO22X2 U12 ( .A0(data2_i[21]), .A1(n6), .B0(n35), .B1(data1_i[21]), .Y(n70)
         );
  NAND2X4 U13 ( .A(data2_i[26]), .B(n6), .Y(n26) );
  AOI22X2 U14 ( .A0(n34), .A1(data2_i[2]), .B0(data0_i[2]), .B1(n44), .Y(n16)
         );
  CLKAND2X4 U15 ( .A(data2_i[16]), .B(n34), .Y(n22) );
  AND2X6 U16 ( .A(n34), .B(data2_i[10]), .Y(n30) );
  MX2X2 U17 ( .A(data0_i[0]), .B(data2_i[0]), .S0(select_i[1]), .Y(n10) );
  OAI2BB1X4 U18 ( .A0N(data1_i[2]), .A1N(n35), .B0(n16), .Y(data_o[2]) );
  NAND2X4 U19 ( .A(n6), .B(data2_i[5]), .Y(n68) );
  NAND2X6 U20 ( .A(data0_i[4]), .B(n57), .Y(n64) );
  NAND2X4 U21 ( .A(data0_i[5]), .B(n57), .Y(n67) );
  NAND2X2 U22 ( .A(n26), .B(n27), .Y(n73) );
  AND2X2 U23 ( .A(data0_i[28]), .B(n3), .Y(n28) );
  NAND2X2 U24 ( .A(n8), .B(n9), .Y(n40) );
  INVX4 U25 ( .A(data2_i[17]), .Y(n18) );
  INVX4 U26 ( .A(data2_i[15]), .Y(n4) );
  INVX6 U27 ( .A(data2_i[22]), .Y(n7) );
  NOR2X4 U28 ( .A(n22), .B(n23), .Y(n55) );
  BUFX20 U29 ( .A(n35), .Y(n5) );
  OAI2BB1X4 U30 ( .A0N(data0_i[8]), .A1N(n3), .B0(n48), .Y(data_o[8]) );
  NAND2X8 U31 ( .A(n60), .B(n56), .Y(n17) );
  INVX12 U32 ( .A(n6), .Y(n19) );
  INVX12 U33 ( .A(select_i[1]), .Y(n60) );
  NAND2X6 U34 ( .A(n59), .B(n33), .Y(data_o[0]) );
  NOR2X6 U35 ( .A(n24), .B(n25), .Y(n48) );
  AOI22X4 U36 ( .A0(n2), .A1(data2_i[9]), .B0(n5), .B1(data1_i[9]), .Y(n50) );
  OAI2BB1X4 U37 ( .A0N(data1_i[1]), .A1N(n5), .B0(n1), .Y(data_o[1]) );
  CLKAND2X12 U38 ( .A(n13), .B(n14), .Y(n1) );
  OR2X6 U39 ( .A(n28), .B(n74), .Y(data_o[28]) );
  NAND2X2 U40 ( .A(n35), .B(data1_i[26]), .Y(n27) );
  AOI22X4 U41 ( .A0(data2_i[11]), .A1(n34), .B0(data1_i[11]), .B1(n35), .Y(n45) );
  OAI2BB1X4 U42 ( .A0N(data0_i[13]), .A1N(n57), .B0(n46), .Y(data_o[13]) );
  AO22X4 U43 ( .A0(data2_i[31]), .A1(n2), .B0(data1_i[31]), .B1(n5), .Y(n75)
         );
  NAND2X2 U44 ( .A(data2_i[20]), .B(n6), .Y(n8) );
  AOI22X2 U45 ( .A0(data2_i[13]), .A1(n34), .B0(data1_i[13]), .B1(n35), .Y(n46) );
  BUFX12 U46 ( .A(n44), .Y(n3) );
  BUFX20 U47 ( .A(n44), .Y(n57) );
  NAND3X6 U48 ( .A(n64), .B(n65), .C(n63), .Y(data_o[4]) );
  INVX20 U49 ( .A(n20), .Y(n6) );
  INVX16 U50 ( .A(n20), .Y(n34) );
  AND2X4 U51 ( .A(n56), .B(n60), .Y(n11) );
  AND2X8 U52 ( .A(n32), .B(n60), .Y(n44) );
  AOI2BB2X4 U53 ( .B0(data1_i[15]), .B1(n5), .A0N(n4), .A1N(n19), .Y(n53) );
  NAND2X8 U54 ( .A(n67), .B(n12), .Y(data_o[5]) );
  CLKAND2X12 U55 ( .A(n66), .B(n68), .Y(n12) );
  CLKINVX12 U56 ( .A(n60), .Y(n21) );
  NAND2X2 U57 ( .A(data1_i[4]), .B(n35), .Y(n63) );
  NAND2X2 U58 ( .A(n32), .B(n10), .Y(n33) );
  OAI2BB2X4 U59 ( .B0(n7), .B1(n19), .A0N(data1_i[22]), .A1N(n35), .Y(n37) );
  NAND2X2 U60 ( .A(data1_i[20]), .B(n35), .Y(n9) );
  AOI22X4 U61 ( .A0(data2_i[3]), .A1(n21), .B0(data0_i[3]), .B1(n60), .Y(n62)
         );
  AO22X4 U62 ( .A0(data2_i[27]), .A1(n6), .B0(data1_i[27]), .B1(n35), .Y(n36)
         );
  CLKAND2X3 U63 ( .A(data0_i[31]), .B(n3), .Y(n29) );
  OAI2BB1X4 U64 ( .A0N(data0_i[11]), .A1N(n57), .B0(n45), .Y(data_o[11]) );
  CLKINVX1 U65 ( .A(n32), .Y(n15) );
  OAI2BB1X4 U66 ( .A0N(data0_i[9]), .A1N(n3), .B0(n50), .Y(data_o[9]) );
  OAI21X4 U67 ( .A0(n15), .A1(n62), .B0(n61), .Y(data_o[3]) );
  AOI22X2 U68 ( .A0(n6), .A1(data2_i[6]), .B0(n35), .B1(data1_i[6]), .Y(n54)
         );
  OR2X8 U69 ( .A(n29), .B(n75), .Y(data_o[31]) );
  NAND2X2 U70 ( .A(n44), .B(data0_i[1]), .Y(n14) );
  OAI2BB1X4 U71 ( .A0N(data0_i[15]), .A1N(n58), .B0(n53), .Y(data_o[15]) );
  AOI22X2 U72 ( .A0(data2_i[18]), .A1(n34), .B0(data1_i[18]), .B1(n35), .Y(n49) );
  NAND2X2 U73 ( .A(n11), .B(data1_i[5]), .Y(n66) );
  OAI2BB1X4 U74 ( .A0N(data0_i[12]), .A1N(n57), .B0(n47), .Y(data_o[12]) );
  INVX20 U75 ( .A(n56), .Y(n32) );
  NAND2X8 U76 ( .A(n32), .B(n21), .Y(n20) );
  AO22X4 U77 ( .A0(data2_i[7]), .A1(n6), .B0(data1_i[7]), .B1(n35), .Y(n43) );
  AOI2BB2X4 U78 ( .B0(data1_i[17]), .B1(n5), .A0N(n19), .A1N(n18), .Y(n51) );
  AO22X2 U79 ( .A0(data2_i[29]), .A1(n34), .B0(data1_i[29]), .B1(n35), .Y(n42)
         );
  OAI2BB1X4 U80 ( .A0N(data0_i[17]), .A1N(n58), .B0(n51), .Y(data_o[17]) );
  OAI2BB1X4 U81 ( .A0N(data0_i[6]), .A1N(n57), .B0(n54), .Y(data_o[6]) );
  AO22X4 U82 ( .A0(data2_i[19]), .A1(n34), .B0(data1_i[19]), .B1(n35), .Y(n38)
         );
  AO21X4 U83 ( .A0(data0_i[27]), .A1(n3), .B0(n36), .Y(data_o[27]) );
  NOR2X6 U84 ( .A(n30), .B(n31), .Y(n52) );
  AO22X4 U85 ( .A0(data2_i[24]), .A1(n6), .B0(data1_i[24]), .B1(n35), .Y(n71)
         );
  AO21X4 U86 ( .A0(data0_i[19]), .A1(n58), .B0(n38), .Y(data_o[19]) );
  AOI22X2 U87 ( .A0(data2_i[12]), .A1(n34), .B0(data1_i[12]), .B1(n35), .Y(n47) );
  NAND3BX2 U88 ( .AN(n21), .B(n56), .C(data1_i[3]), .Y(n61) );
  OAI2BB1X4 U89 ( .A0N(data0_i[18]), .A1N(n57), .B0(n49), .Y(data_o[18]) );
  AO22X4 U90 ( .A0(data2_i[23]), .A1(n6), .B0(data1_i[23]), .B1(n35), .Y(n41)
         );
  NAND2X2 U91 ( .A(data2_i[4]), .B(n34), .Y(n65) );
  AO22X4 U92 ( .A0(data2_i[25]), .A1(n34), .B0(data1_i[25]), .B1(n35), .Y(n72)
         );
  AO22X4 U93 ( .A0(data2_i[14]), .A1(n34), .B0(data1_i[14]), .B1(n35), .Y(n69)
         );
  INVX20 U94 ( .A(n17), .Y(n35) );
  OAI2BB1X4 U95 ( .A0N(data0_i[16]), .A1N(n58), .B0(n55), .Y(data_o[16]) );
  OAI2BB1X4 U96 ( .A0N(data0_i[10]), .A1N(n3), .B0(n52), .Y(data_o[10]) );
  AO21X4 U97 ( .A0(data0_i[14]), .A1(n58), .B0(n69), .Y(data_o[14]) );
  AO21X4 U98 ( .A0(data0_i[23]), .A1(n57), .B0(n41), .Y(data_o[23]) );
  AO21X4 U99 ( .A0(data0_i[30]), .A1(n58), .B0(n39), .Y(data_o[30]) );
  AO21X4 U100 ( .A0(data0_i[22]), .A1(n58), .B0(n37), .Y(data_o[22]) );
  AO21X4 U101 ( .A0(data0_i[21]), .A1(n58), .B0(n70), .Y(data_o[21]) );
  AO21X4 U102 ( .A0(data0_i[29]), .A1(n58), .B0(n42), .Y(data_o[29]) );
  AO21X4 U103 ( .A0(data0_i[20]), .A1(n57), .B0(n40), .Y(data_o[20]) );
  AO21X4 U104 ( .A0(data0_i[7]), .A1(n3), .B0(n43), .Y(data_o[7]) );
  BUFX20 U105 ( .A(select_i[0]), .Y(n56) );
  AO21X4 U106 ( .A0(data0_i[24]), .A1(n57), .B0(n71), .Y(data_o[24]) );
  AO21X4 U107 ( .A0(data0_i[25]), .A1(n58), .B0(n72), .Y(data_o[25]) );
  AO21X4 U108 ( .A0(data0_i[26]), .A1(n58), .B0(n73), .Y(data_o[26]) );
endmodule


module forwarding ( Rs_regD, Rt_regD, RegWrite_regE, wsel_regE, RegWrite_regM, 
        wsel_regM, FU_Asel, FU_Bsel );
  input [4:0] Rs_regD;
  input [4:0] Rt_regD;
  input [4:0] wsel_regE;
  input [4:0] wsel_regM;
  output [1:0] FU_Asel;
  output [1:0] FU_Bsel;
  input RegWrite_regE, RegWrite_regM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66;

  AND2X6 U2 ( .A(n51), .B(n32), .Y(n8) );
  NAND3X8 U3 ( .A(n50), .B(n48), .C(n49), .Y(n54) );
  BUFX8 U4 ( .A(n13), .Y(n6) );
  AND2X8 U5 ( .A(n23), .B(n22), .Y(n50) );
  INVX16 U6 ( .A(wsel_regE[4]), .Y(n13) );
  CLKINVX4 U7 ( .A(wsel_regM[2]), .Y(n60) );
  NAND2X4 U8 ( .A(n14), .B(n15), .Y(n23) );
  NAND2X4 U9 ( .A(n63), .B(n62), .Y(n64) );
  NAND2X4 U10 ( .A(n60), .B(n16), .Y(n17) );
  XOR2X1 U11 ( .A(Rs_regD[0]), .B(wsel_regM[0]), .Y(n65) );
  NAND2X6 U12 ( .A(n52), .B(RegWrite_regE), .Y(n53) );
  INVX12 U13 ( .A(wsel_regM[4]), .Y(n18) );
  INVX4 U14 ( .A(wsel_regE[3]), .Y(n33) );
  INVX12 U15 ( .A(wsel_regE[1]), .Y(n47) );
  NAND4X4 U16 ( .A(n18), .B(n56), .C(n55), .D(n24), .Y(n29) );
  OR2X8 U17 ( .A(n64), .B(n65), .Y(n1) );
  NAND3X8 U18 ( .A(n34), .B(n33), .C(n7), .Y(n36) );
  INVX16 U19 ( .A(wsel_regM[3]), .Y(n56) );
  NAND2X2 U20 ( .A(Rs_regD[2]), .B(wsel_regM[2]), .Y(n2) );
  NAND2X4 U21 ( .A(n11), .B(n10), .Y(n25) );
  NAND2X4 U22 ( .A(n13), .B(n12), .Y(n15) );
  NAND3X4 U23 ( .A(n36), .B(n35), .C(n37), .Y(n3) );
  NAND3X6 U24 ( .A(n36), .B(n35), .C(n37), .Y(n43) );
  NOR3X8 U25 ( .A(FU_Asel[1]), .B(n1), .C(n66), .Y(FU_Asel[0]) );
  NAND4X6 U26 ( .A(RegWrite_regM), .B(n59), .C(n58), .D(n57), .Y(n66) );
  AND2X6 U27 ( .A(n4), .B(n5), .Y(n28) );
  XNOR2X4 U28 ( .A(Rt_regD[1]), .B(wsel_regM[1]), .Y(n4) );
  XNOR2X4 U29 ( .A(Rt_regD[0]), .B(wsel_regM[0]), .Y(n5) );
  INVX8 U30 ( .A(wsel_regE[0]), .Y(n51) );
  XNOR2X4 U31 ( .A(wsel_regE[0]), .B(Rt_regD[0]), .Y(n38) );
  NOR2X4 U32 ( .A(wsel_regE[1]), .B(wsel_regE[2]), .Y(n7) );
  INVX12 U33 ( .A(wsel_regE[2]), .Y(n32) );
  NOR2X6 U34 ( .A(wsel_regM[2]), .B(wsel_regM[1]), .Y(n24) );
  INVX4 U35 ( .A(Rt_regD[3]), .Y(n9) );
  INVX8 U36 ( .A(Rs_regD[4]), .Y(n12) );
  NAND4X4 U37 ( .A(n8), .B(n33), .C(n6), .D(n47), .Y(n48) );
  XNOR2X4 U38 ( .A(n47), .B(Rs_regD[1]), .Y(n45) );
  XOR2X4 U39 ( .A(n32), .B(Rs_regD[2]), .Y(n22) );
  XOR2X4 U40 ( .A(n18), .B(Rs_regD[4]), .Y(n57) );
  NAND2X2 U41 ( .A(wsel_regE[4]), .B(Rs_regD[4]), .Y(n14) );
  NAND4X8 U42 ( .A(n39), .B(n40), .C(n38), .D(RegWrite_regE), .Y(n44) );
  CLKINVX6 U43 ( .A(Rt_regD[4]), .Y(n19) );
  CLKINVX3 U44 ( .A(Rs_regD[2]), .Y(n16) );
  NAND2X6 U45 ( .A(n56), .B(n9), .Y(n11) );
  XOR2X4 U46 ( .A(n32), .B(Rt_regD[2]), .Y(n37) );
  CLKINVX3 U47 ( .A(wsel_regM[1]), .Y(n61) );
  NAND4X8 U48 ( .A(n28), .B(n30), .C(n31), .D(n29), .Y(n42) );
  NOR2X8 U49 ( .A(n46), .B(n45), .Y(n49) );
  NOR2X8 U50 ( .A(n44), .B(n43), .Y(n41) );
  XOR2X4 U51 ( .A(wsel_regE[3]), .B(Rs_regD[3]), .Y(n46) );
  NAND2X6 U52 ( .A(n19), .B(n18), .Y(n21) );
  NAND2X6 U53 ( .A(n21), .B(n20), .Y(n27) );
  NAND2X4 U54 ( .A(wsel_regM[4]), .B(Rt_regD[4]), .Y(n20) );
  XNOR2X4 U55 ( .A(wsel_regM[2]), .B(Rt_regD[2]), .Y(n26) );
  NAND2X4 U56 ( .A(n17), .B(n2), .Y(n63) );
  NOR2X4 U57 ( .A(wsel_regE[0]), .B(wsel_regE[4]), .Y(n34) );
  NAND4X4 U58 ( .A(n18), .B(n55), .C(n56), .D(n24), .Y(n59) );
  XOR2X4 U59 ( .A(n56), .B(Rs_regD[3]), .Y(n58) );
  XNOR2X4 U60 ( .A(Rt_regD[3]), .B(wsel_regE[3]), .Y(n35) );
  NOR2X8 U61 ( .A(n54), .B(n53), .Y(FU_Asel[1]) );
  AND2X8 U62 ( .A(n26), .B(n27), .Y(n30) );
  XOR2X4 U63 ( .A(n61), .B(Rs_regD[1]), .Y(n62) );
  INVX6 U64 ( .A(wsel_regM[0]), .Y(n55) );
  NAND2X2 U65 ( .A(Rt_regD[3]), .B(wsel_regM[3]), .Y(n10) );
  AND2X8 U66 ( .A(n25), .B(RegWrite_regM), .Y(n31) );
  NOR2X8 U67 ( .A(n3), .B(n44), .Y(FU_Bsel[1]) );
  XOR2X4 U68 ( .A(n51), .B(Rs_regD[0]), .Y(n52) );
  NOR2X8 U69 ( .A(n42), .B(n41), .Y(FU_Bsel[0]) );
  XOR2X4 U70 ( .A(n47), .B(Rt_regD[1]), .Y(n40) );
  XOR2X4 U71 ( .A(n13), .B(Rt_regD[4]), .Y(n39) );
endmodule


module hazard_detection ( Branch_EX, equal, branchpred_his, JumpReg_regD, 
        MemRead_regD, Rt_regD, Rs, Rt, ICACHE_stall, DCACHE_stall, 
        stall_lw_use, stallcache, flush, pred_cond, stall_muldiv );
  input [4:0] Rt_regD;
  input [4:0] Rs;
  input [4:0] Rt;
  input Branch_EX, equal, branchpred_his, JumpReg_regD, MemRead_regD,
         ICACHE_stall, DCACHE_stall, stall_muldiv;
  output stall_lw_use, stallcache, flush, pred_cond;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;

  INVX2 U2 ( .A(Rt_regD[3]), .Y(n9) );
  XOR2X4 U3 ( .A(equal), .B(n3), .Y(n1) );
  INVX4 U4 ( .A(Rt_regD[2]), .Y(n8) );
  CLKINVX1 U5 ( .A(branchpred_his), .Y(n3) );
  AO21X4 U6 ( .A0(n20), .A1(n2), .B0(JumpReg_regD), .Y(flush) );
  NOR2XL U7 ( .A(n4), .B(n1), .Y(n2) );
  OR3X6 U8 ( .A(DCACHE_stall), .B(ICACHE_stall), .C(stall_muldiv), .Y(
        stallcache) );
  NOR2X8 U9 ( .A(n20), .B(JumpReg_regD), .Y(stall_lw_use) );
  XOR2XL U10 ( .A(Rt[1]), .B(Rt_regD[1]), .Y(n14) );
  XOR2XL U11 ( .A(Rt[4]), .B(Rt_regD[4]), .Y(n13) );
  XOR2XL U12 ( .A(Rs[1]), .B(Rt_regD[1]), .Y(n17) );
  XOR2XL U13 ( .A(Rs[4]), .B(Rt_regD[4]), .Y(n16) );
  XOR2X1 U14 ( .A(n9), .B(Rt[3]), .Y(n10) );
  XOR2X1 U15 ( .A(n8), .B(Rt[2]), .Y(n11) );
  XOR2XL U16 ( .A(Rt[0]), .B(Rt_regD[0]), .Y(n12) );
  XOR2X1 U17 ( .A(n9), .B(Rs[3]), .Y(n5) );
  XOR2X1 U18 ( .A(n8), .B(Rs[2]), .Y(n6) );
  XOR2XL U19 ( .A(Rs[0]), .B(Rt_regD[0]), .Y(n7) );
  NOR2X8 U20 ( .A(n1), .B(n4), .Y(pred_cond) );
  CLKINVX6 U21 ( .A(Branch_EX), .Y(n4) );
  NAND3BX2 U22 ( .AN(n7), .B(n6), .C(n5), .Y(n18) );
  NAND3BX2 U23 ( .AN(n12), .B(n11), .C(n10), .Y(n15) );
  OAI33X2 U24 ( .A0(n18), .A1(n17), .A2(n16), .B0(n15), .B1(n14), .B2(n13), 
        .Y(n19) );
  NAND2X2 U25 ( .A(MemRead_regD), .B(n19), .Y(n20) );
endmodule


module branch_prediction ( clk, rst_n, branch, equal, predict, branchpred_his
 );
  input clk, rst_n, branch, equal;
  output predict, branchpred_his;
  wire   n9, n10, n1, n2, n3, n4, n6, n7, n8;
  wire   [1:0] state;

  DFFRX1 branchpred_reg_reg ( .D(predict), .CK(clk), .RN(rst_n), .Q(
        branchpred_his) );
  DFFRX1 \state_reg[1]  ( .D(n9), .CK(clk), .RN(rst_n), .Q(state[1]), .QN(
        predict) );
  DFFSX1 \state_reg[0]  ( .D(n10), .CK(clk), .SN(rst_n), .Q(state[0]), .QN(n8)
         );
  INVXL U3 ( .A(equal), .Y(n3) );
  OAI2BB1X1 U4 ( .A0N(n2), .A1N(branch), .B0(n1), .Y(n10) );
  NAND2X1 U5 ( .A(state[0]), .B(n4), .Y(n1) );
  OAI32XL U6 ( .A0(equal), .A1(n8), .A2(n7), .B0(n6), .B1(predict), .Y(n9) );
  INVXL U7 ( .A(branch), .Y(n7) );
  AND3XL U8 ( .A(equal), .B(branch), .C(n8), .Y(n6) );
  OAI21XL U9 ( .A0(predict), .A1(equal), .B0(branch), .Y(n4) );
  AO22X1 U10 ( .A0(state[1]), .A1(n8), .B0(n8), .B1(n3), .Y(n2) );
endmodule


module precontrolDec ( instruction_next, Jump_IF, Branch_IF );
  input [31:0] instruction_next;
  output Jump_IF, Branch_IF;
  wire   n1, n2, n3;

  AND3X8 U1 ( .A(instruction_next[27]), .B(n3), .C(n2), .Y(Jump_IF) );
  INVX6 U2 ( .A(n1), .Y(n3) );
  INVX6 U3 ( .A(instruction_next[28]), .Y(n2) );
  OR3X8 U4 ( .A(instruction_next[30]), .B(instruction_next[31]), .C(
        instruction_next[29]), .Y(n1) );
  NOR4X4 U5 ( .A(instruction_next[27]), .B(instruction_next[26]), .C(n1), .D(
        n2), .Y(Branch_IF) );
endmodule


module nextPCcalculator_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n7, n9, n10, n11, n13, n14, n15, n16, n19, n20, n21, n22,
         n23, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n41, n43, n44, n45, n46, n47, n49, n50, n51, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n69, n70, n72, n73,
         n75, n76, n77, n79, n80, n83, n85, n87, n88, n90, n92, n94, n96, n97,
         n98, n99, n100, n101, n102, n103, n106, n108, n109, n110, n111, n116,
         n117, n118, n119, n120, n122, n123, n124, n125, n126, n127, n128,
         n129, n132, n133, n134, n135, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n152, n153, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n166, n167, n168, n171, n173, n174,
         n179, n180, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n193, n194, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n210, n212, n214, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n351, n352, n353, n354, n357,
         n358, n359;
  assign n23 = A[30];
  assign n29 = A[29];
  assign n33 = A[28];
  assign n39 = A[27];
  assign n43 = A[26];
  assign n51 = A[25];
  assign n55 = A[24];
  assign n61 = A[23];
  assign n65 = A[22];
  assign n73 = A[21];
  assign n77 = A[20];
  assign n83 = A[19];
  assign n87 = A[18];

  OAI21X4 U181 ( .A0(n159), .A1(n187), .B0(n160), .Y(n158) );
  NOR2X8 U188 ( .A(B[9]), .B(A[9]), .Y(n163) );
  AOI21X4 U222 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  NOR2X8 U233 ( .A(B[4]), .B(A[4]), .Y(n193) );
  NOR2X2 U250 ( .A(n123), .B(n116), .Y(n317) );
  NOR2X8 U251 ( .A(A[14]), .B(B[14]), .Y(n123) );
  NAND2X6 U252 ( .A(A[12]), .B(B[12]), .Y(n142) );
  NOR2X6 U253 ( .A(B[12]), .B(A[12]), .Y(n141) );
  NAND2X6 U254 ( .A(A[4]), .B(B[4]), .Y(n194) );
  CLKINVX2 U255 ( .A(n142), .Y(n140) );
  NAND2X4 U256 ( .A(n146), .B(n132), .Y(n126) );
  OAI21X2 U257 ( .A0(n157), .A1(n126), .B0(n345), .Y(n125) );
  XOR2X4 U258 ( .A(n319), .B(n318), .Y(SUM[16]) );
  CLKINVX20 U259 ( .A(n342), .Y(n318) );
  OA21X4 U260 ( .A0(n108), .A1(n157), .B0(n109), .Y(n319) );
  NAND2X2 U261 ( .A(n69), .B(n65), .Y(n64) );
  INVX8 U262 ( .A(n69), .Y(n70) );
  NOR2X8 U263 ( .A(n80), .B(n72), .Y(n69) );
  XOR2X4 U264 ( .A(n35), .B(n320), .Y(SUM[28]) );
  CLKINVX20 U265 ( .A(n34), .Y(n320) );
  NOR2BX4 U266 ( .AN(n321), .B(n1), .Y(n41) );
  CLKAND2X8 U267 ( .A(n47), .B(n43), .Y(n321) );
  OA21X4 U268 ( .A0(n116), .A1(n124), .B0(n117), .Y(n322) );
  NAND2X8 U269 ( .A(B[14]), .B(A[14]), .Y(n124) );
  NAND2X4 U270 ( .A(B[15]), .B(A[15]), .Y(n117) );
  AOI21X4 U271 ( .A0(n129), .A1(n101), .B0(n102), .Y(n100) );
  AOI21X4 U272 ( .A0(n129), .A1(n317), .B0(n359), .Y(n109) );
  NOR2X4 U273 ( .A(n1), .B(n20), .Y(n19) );
  NOR2X2 U274 ( .A(n1), .B(n36), .Y(n35) );
  NOR2X2 U275 ( .A(n1), .B(n58), .Y(n57) );
  CLKINVX2 U276 ( .A(n116), .Y(n203) );
  INVXL U277 ( .A(n134), .Y(n205) );
  INVX3 U278 ( .A(n140), .Y(n323) );
  BUFX4 U279 ( .A(A[0]), .Y(SUM[0]) );
  BUFX4 U280 ( .A(A[1]), .Y(SUM[1]) );
  NAND2X2 U281 ( .A(n212), .B(n185), .Y(n13) );
  OAI2BB1X4 U282 ( .A0N(n173), .A1N(n186), .B0(n324), .Y(n349) );
  OA21X4 U283 ( .A0(n179), .A1(n185), .B0(n180), .Y(n324) );
  AOI21X2 U284 ( .A0(n334), .A1(n206), .B0(n140), .Y(n138) );
  CLKINVX1 U285 ( .A(n145), .Y(n334) );
  XOR2X4 U286 ( .A(n57), .B(n325), .Y(SUM[24]) );
  CLKINVX20 U287 ( .A(n56), .Y(n325) );
  BUFX3 U288 ( .A(n5), .Y(n326) );
  XOR2X1 U289 ( .A(n338), .B(n16), .Y(SUM[3]) );
  XOR2X4 U290 ( .A(n157), .B(n9), .Y(SUM[10]) );
  XNOR2X4 U291 ( .A(n143), .B(n7), .Y(SUM[12]) );
  XOR2X4 U292 ( .A(n327), .B(n14), .Y(SUM[5]) );
  OA21X4 U293 ( .A0(n344), .A1(n193), .B0(n358), .Y(n327) );
  XOR2X2 U294 ( .A(n344), .B(n15), .Y(SUM[4]) );
  NOR2BX4 U295 ( .AN(n87), .B(n1), .Y(n85) );
  OAI21X4 U296 ( .A0(n119), .A1(n157), .B0(n120), .Y(n118) );
  CLKINVX3 U297 ( .A(n129), .Y(n345) );
  INVX6 U298 ( .A(n210), .Y(n328) );
  INVX8 U299 ( .A(n168), .Y(n210) );
  XOR2X4 U300 ( .A(n330), .B(n329), .Y(SUM[11]) );
  NAND2X2 U301 ( .A(n207), .B(n153), .Y(n329) );
  OA21X4 U302 ( .A0(n157), .A1(n155), .B0(n156), .Y(n330) );
  XNOR2X4 U303 ( .A(n331), .B(n6), .Y(SUM[13]) );
  OAI21X4 U304 ( .A0(n157), .A1(n137), .B0(n138), .Y(n331) );
  OR2XL U305 ( .A(n346), .B(A[7]), .Y(n337) );
  NOR2X6 U306 ( .A(n155), .B(n152), .Y(n146) );
  NOR2X6 U307 ( .A(n46), .B(n38), .Y(n37) );
  INVX3 U308 ( .A(n357), .Y(n358) );
  AND2X4 U309 ( .A(n201), .B(n97), .Y(n343) );
  NAND2X1 U310 ( .A(n340), .B(n164), .Y(n10) );
  CLKINVX1 U311 ( .A(n44), .Y(n336) );
  CLKINVX1 U312 ( .A(n66), .Y(n335) );
  INVX2 U313 ( .A(n187), .Y(n186) );
  NAND2X6 U314 ( .A(n77), .B(n73), .Y(n72) );
  NAND2BX4 U315 ( .AN(n80), .B(n77), .Y(n76) );
  INVX4 U316 ( .A(n37), .Y(n36) );
  NAND2X2 U317 ( .A(n37), .B(n33), .Y(n32) );
  OA21X2 U318 ( .A0(n179), .A1(n185), .B0(n180), .Y(n332) );
  NOR2BX1 U319 ( .AN(n173), .B(n328), .Y(n166) );
  NOR2X8 U320 ( .A(n103), .B(n96), .Y(n94) );
  OAI2BB1X4 U321 ( .A0N(n111), .A1N(n94), .B0(n333), .Y(n339) );
  OA21X4 U322 ( .A0(n96), .A1(n106), .B0(n97), .Y(n333) );
  NAND2X6 U323 ( .A(n346), .B(A[7]), .Y(n180) );
  NAND2X8 U324 ( .A(n110), .B(n94), .Y(n92) );
  OR2XL U325 ( .A(A[9]), .B(B[9]), .Y(n340) );
  NAND2X4 U326 ( .A(B[13]), .B(A[13]), .Y(n135) );
  NOR2X8 U327 ( .A(B[13]), .B(A[13]), .Y(n134) );
  NAND2X6 U328 ( .A(n161), .B(n173), .Y(n159) );
  XNOR2X2 U329 ( .A(n186), .B(n13), .Y(SUM[6]) );
  NOR2X8 U330 ( .A(n141), .B(n134), .Y(n132) );
  AOI21X4 U331 ( .A0(n174), .A1(n161), .B0(n162), .Y(n160) );
  CLKINVX4 U332 ( .A(n147), .Y(n145) );
  XOR2X4 U333 ( .A(n67), .B(n335), .Y(SUM[22]) );
  XOR2X4 U334 ( .A(n45), .B(n336), .Y(SUM[26]) );
  NAND2BXL U335 ( .AN(n197), .B(n198), .Y(n16) );
  BUFX16 U336 ( .A(B[7]), .Y(n346) );
  NOR2X8 U337 ( .A(B[3]), .B(A[3]), .Y(n197) );
  NOR2X6 U338 ( .A(B[10]), .B(A[10]), .Y(n155) );
  XOR2X4 U339 ( .A(n79), .B(n77), .Y(SUM[20]) );
  XOR2X2 U340 ( .A(n1), .B(n88), .Y(SUM[18]) );
  INVX2 U341 ( .A(n351), .Y(n338) );
  INVX1 U342 ( .A(n200), .Y(n351) );
  NAND2X6 U343 ( .A(B[2]), .B(A[2]), .Y(n200) );
  AOI2BB1X4 U344 ( .A0N(n127), .A1N(n92), .B0(n339), .Y(n348) );
  INVXL U345 ( .A(n185), .Y(n183) );
  NOR2X2 U346 ( .A(n1), .B(n26), .Y(n25) );
  NOR2X2 U347 ( .A(n1), .B(n80), .Y(n79) );
  INVX6 U348 ( .A(n126), .Y(n128) );
  NOR2X2 U349 ( .A(n1), .B(n76), .Y(n75) );
  OA21X1 U350 ( .A0(n200), .A1(n197), .B0(n198), .Y(n344) );
  NAND2X1 U351 ( .A(n128), .B(n317), .Y(n108) );
  NAND2BXL U352 ( .AN(n155), .B(n156), .Y(n9) );
  AOI21X4 U353 ( .A0(n129), .A1(n204), .B0(n122), .Y(n120) );
  INVX4 U354 ( .A(n127), .Y(n129) );
  NOR2X8 U355 ( .A(B[17]), .B(A[17]), .Y(n96) );
  NOR2X4 U356 ( .A(n126), .B(n92), .Y(n90) );
  XOR2X4 U357 ( .A(n118), .B(n341), .Y(SUM[15]) );
  CLKAND2X8 U358 ( .A(n203), .B(n117), .Y(n341) );
  CLKAND2X8 U359 ( .A(n202), .B(n106), .Y(n342) );
  XOR2X4 U360 ( .A(n98), .B(n343), .Y(SUM[17]) );
  NOR2X8 U361 ( .A(B[11]), .B(A[11]), .Y(n152) );
  NAND2X1 U362 ( .A(n59), .B(n55), .Y(n54) );
  INVX4 U363 ( .A(n59), .Y(n58) );
  NOR2X8 U364 ( .A(n70), .B(n60), .Y(n59) );
  INVX16 U365 ( .A(n347), .Y(n1) );
  INVX6 U366 ( .A(n141), .Y(n206) );
  OAI21X4 U367 ( .A0(n157), .A1(n144), .B0(n145), .Y(n143) );
  XOR2X4 U368 ( .A(n53), .B(n51), .Y(SUM[25]) );
  NOR2X2 U369 ( .A(n46), .B(n22), .Y(n21) );
  AND2X1 U370 ( .A(n337), .B(n180), .Y(n353) );
  NAND2X6 U371 ( .A(B[10]), .B(A[10]), .Y(n156) );
  XOR2X4 U372 ( .A(n63), .B(n61), .Y(SUM[23]) );
  INVX3 U373 ( .A(n21), .Y(n20) );
  NOR2X8 U374 ( .A(n184), .B(n179), .Y(n173) );
  NOR2X6 U375 ( .A(n193), .B(n190), .Y(n188) );
  XOR2X4 U376 ( .A(n85), .B(n83), .Y(SUM[19]) );
  INVX4 U377 ( .A(n46), .Y(n47) );
  NAND2X2 U378 ( .A(n101), .B(n128), .Y(n99) );
  NOR2X2 U379 ( .A(n1), .B(n70), .Y(n67) );
  OAI21X2 U380 ( .A0(n322), .A1(n103), .B0(n106), .Y(n102) );
  NAND2X6 U381 ( .A(B[16]), .B(A[16]), .Y(n106) );
  NOR2X8 U382 ( .A(n346), .B(A[7]), .Y(n179) );
  NAND2X8 U383 ( .A(A[6]), .B(B[6]), .Y(n185) );
  OAI21X4 U384 ( .A0(n171), .A1(n163), .B0(n164), .Y(n162) );
  NOR2X8 U385 ( .A(n168), .B(n163), .Y(n161) );
  NOR2X8 U386 ( .A(n38), .B(n28), .Y(n27) );
  NAND2X4 U387 ( .A(n33), .B(n29), .Y(n28) );
  XOR2X4 U388 ( .A(n19), .B(A[31]), .Y(SUM[31]) );
  NOR2X8 U389 ( .A(B[16]), .B(A[16]), .Y(n103) );
  NOR2BX4 U390 ( .AN(n110), .B(n103), .Y(n101) );
  INVX6 U391 ( .A(n123), .Y(n204) );
  XNOR2X4 U392 ( .A(n125), .B(n326), .Y(SUM[14]) );
  NOR2X8 U393 ( .A(B[8]), .B(A[8]), .Y(n168) );
  NOR2X2 U394 ( .A(n1), .B(n32), .Y(n31) );
  XOR2X4 U395 ( .A(n31), .B(n29), .Y(SUM[29]) );
  INVX8 U396 ( .A(n158), .Y(n157) );
  XOR2X4 U397 ( .A(n25), .B(n23), .Y(SUM[30]) );
  NAND2X6 U398 ( .A(n43), .B(n39), .Y(n38) );
  AO21X4 U399 ( .A0(n186), .A1(n166), .B0(n167), .Y(n354) );
  XNOR2X4 U400 ( .A(n349), .B(n11), .Y(SUM[8]) );
  AO21X4 U401 ( .A0(n186), .A1(n212), .B0(n183), .Y(n352) );
  OAI21X4 U402 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X8 U403 ( .A(B[5]), .B(A[5]), .Y(n190) );
  OAI21X2 U404 ( .A0(n332), .A1(n328), .B0(n171), .Y(n167) );
  NOR2X8 U405 ( .A(A[15]), .B(B[15]), .Y(n116) );
  XNOR2X4 U406 ( .A(n354), .B(n10), .Y(SUM[9]) );
  XOR2X4 U407 ( .A(n41), .B(n39), .Y(SUM[27]) );
  NOR2X2 U408 ( .A(n1), .B(n46), .Y(n45) );
  NAND2X2 U409 ( .A(B[17]), .B(A[17]), .Y(n97) );
  OAI21X2 U410 ( .A0(n99), .A1(n157), .B0(n100), .Y(n98) );
  NOR2X8 U411 ( .A(n123), .B(n116), .Y(n110) );
  NOR2X2 U412 ( .A(n1), .B(n54), .Y(n53) );
  NAND2X6 U413 ( .A(B[8]), .B(A[8]), .Y(n171) );
  NAND2X4 U414 ( .A(n65), .B(n61), .Y(n60) );
  XOR2X4 U415 ( .A(n75), .B(n73), .Y(SUM[21]) );
  NAND2X4 U416 ( .A(B[11]), .B(A[11]), .Y(n153) );
  OAI21X4 U417 ( .A0(n134), .A1(n142), .B0(n135), .Y(n133) );
  NOR2X2 U418 ( .A(n1), .B(n64), .Y(n63) );
  NAND2X6 U419 ( .A(n69), .B(n49), .Y(n46) );
  NAND2X4 U420 ( .A(B[9]), .B(A[9]), .Y(n164) );
  NAND2X4 U421 ( .A(B[3]), .B(A[3]), .Y(n198) );
  NOR2X4 U422 ( .A(A[6]), .B(B[6]), .Y(n184) );
  NAND2X6 U423 ( .A(n87), .B(n83), .Y(n80) );
  AOI21X4 U424 ( .A0(n132), .A1(n147), .B0(n133), .Y(n127) );
  NAND2X1 U425 ( .A(n128), .B(n204), .Y(n119) );
  NAND2XL U426 ( .A(n205), .B(n135), .Y(n6) );
  OAI21X4 U427 ( .A0(n152), .A1(n156), .B0(n153), .Y(n147) );
  OAI2BB1X4 U428 ( .A0N(n158), .A1N(n90), .B0(n348), .Y(n347) );
  NAND2XL U429 ( .A(n206), .B(n323), .Y(n7) );
  OAI21X4 U430 ( .A0(n116), .A1(n124), .B0(n117), .Y(n111) );
  NAND2X2 U431 ( .A(n214), .B(n358), .Y(n15) );
  OAI21X4 U432 ( .A0(n179), .A1(n185), .B0(n180), .Y(n174) );
  OAI21X4 U433 ( .A0(n197), .A1(n200), .B0(n198), .Y(n196) );
  INVXL U434 ( .A(n152), .Y(n207) );
  NAND2XL U435 ( .A(n204), .B(n124), .Y(n5) );
  INVXL U436 ( .A(n124), .Y(n122) );
  NAND2BXL U437 ( .AN(n190), .B(n191), .Y(n14) );
  NOR2X2 U438 ( .A(n60), .B(n50), .Y(n49) );
  NAND2X1 U439 ( .A(n146), .B(n206), .Y(n137) );
  CLKINVX1 U440 ( .A(n146), .Y(n144) );
  NAND2X1 U441 ( .A(n210), .B(n171), .Y(n11) );
  CLKINVX1 U442 ( .A(n96), .Y(n201) );
  CLKINVX1 U443 ( .A(n103), .Y(n202) );
  NOR2X1 U444 ( .A(n199), .B(n351), .Y(SUM[2]) );
  CLKINVX1 U445 ( .A(n184), .Y(n212) );
  NAND2X1 U446 ( .A(n47), .B(n27), .Y(n26) );
  XOR2X4 U447 ( .A(n352), .B(n353), .Y(SUM[7]) );
  INVXL U448 ( .A(n193), .Y(n214) );
  CLKINVX1 U449 ( .A(n194), .Y(n357) );
  NAND2X1 U450 ( .A(n55), .B(n51), .Y(n50) );
  CLKINVX1 U451 ( .A(n87), .Y(n88) );
  CLKINVX1 U452 ( .A(n65), .Y(n66) );
  CLKINVX1 U453 ( .A(n55), .Y(n56) );
  NAND2X1 U454 ( .A(n27), .B(n23), .Y(n22) );
  CLKINVX1 U455 ( .A(n33), .Y(n34) );
  CLKINVX1 U456 ( .A(n43), .Y(n44) );
  CLKBUFX2 U457 ( .A(n111), .Y(n359) );
  NOR2XL U458 ( .A(A[2]), .B(B[2]), .Y(n199) );
  NAND2X4 U459 ( .A(B[5]), .B(A[5]), .Y(n191) );
endmodule


module nextPCcalculator ( PCcur, PCplus4, PCplus4_regD, targetAddr, 
        branchOffset_I, branchOffset_regD, JumpRegAddr, PCsrc, PCnext );
  input [31:0] PCcur;
  input [31:0] PCplus4;
  input [31:0] PCplus4_regD;
  input [25:0] targetAddr;
  input [15:0] branchOffset_I;
  input [15:0] branchOffset_regD;
  input [31:0] JumpRegAddr;
  input [2:0] PCsrc;
  output [31:0] PCnext;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179;
  wire   [31:0] PCplus4_actual;
  wire   [17:2] branchOffset_actual;
  wire   [31:0] ADDresult;

  nextPCcalculator_DW01_add_1 add_1660 ( .A(PCplus4_actual), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        branchOffset_actual, 1'b0, 1'b0}), .CI(1'b0), .SUM(ADDresult) );
  MX2X8 U4 ( .A(PCplus4_regD[3]), .B(PCplus4[3]), .S0(n41), .Y(
        PCplus4_actual[3]) );
  MX2X6 U5 ( .A(PCplus4_regD[5]), .B(PCplus4[5]), .S0(n41), .Y(
        PCplus4_actual[5]) );
  MX2X6 U6 ( .A(PCplus4_regD[7]), .B(PCplus4[7]), .S0(n1), .Y(
        PCplus4_actual[7]) );
  AOI222X4 U7 ( .A0(PCplus4_regD[16]), .A1(n152), .B0(targetAddr[14]), .B1(n31), .C0(JumpRegAddr[16]), .C1(n39), .Y(n110) );
  NAND3BX2 U8 ( .AN(n53), .B(n13), .C(n52), .Y(n158) );
  CLKINVX1 U9 ( .A(PCsrc[0]), .Y(n42) );
  INVX12 U10 ( .A(n10), .Y(n1) );
  INVX12 U11 ( .A(n10), .Y(n41) );
  INVX3 U12 ( .A(n166), .Y(n20) );
  NAND3X4 U13 ( .A(n165), .B(n164), .C(n163), .Y(n166) );
  NAND2X2 U14 ( .A(n178), .B(ADDresult[10]), .Y(n85) );
  MX2X6 U15 ( .A(PCplus4_regD[17]), .B(PCplus4[17]), .S0(n30), .Y(
        PCplus4_actual[17]) );
  CLKMX2X4 U16 ( .A(PCplus4_regD[6]), .B(PCplus4[6]), .S0(n1), .Y(
        PCplus4_actual[6]) );
  MX2XL U17 ( .A(PCplus4_regD[0]), .B(PCplus4[0]), .S0(n30), .Y(
        PCplus4_actual[0]) );
  MX2X8 U18 ( .A(PCplus4_regD[13]), .B(PCplus4[13]), .S0(n12), .Y(
        PCplus4_actual[13]) );
  INVX4 U19 ( .A(n53), .Y(n27) );
  MX2X8 U20 ( .A(branchOffset_regD[10]), .B(branchOffset_I[10]), .S0(n12), .Y(
        branchOffset_actual[12]) );
  MX2X8 U21 ( .A(branchOffset_regD[3]), .B(branchOffset_I[3]), .S0(n1), .Y(
        branchOffset_actual[5]) );
  CLKINVX1 U22 ( .A(n9), .Y(n14) );
  INVX16 U23 ( .A(n116), .Y(n178) );
  CLKINVX8 U24 ( .A(n43), .Y(n173) );
  BUFX20 U25 ( .A(n173), .Y(n38) );
  AOI22X1 U26 ( .A0(n174), .A1(PCplus4[31]), .B0(JumpRegAddr[31]), .B1(n38), 
        .Y(n175) );
  AOI222X1 U27 ( .A0(PCplus4_regD[27]), .A1(n152), .B0(targetAddr[25]), .B1(
        n32), .C0(JumpRegAddr[27]), .C1(n38), .Y(n155) );
  AOI222X2 U28 ( .A0(PCplus4_regD[1]), .A1(n152), .B0(ADDresult[1]), .B1(n178), 
        .C0(JumpRegAddr[1]), .C1(n38), .Y(n50) );
  AOI2BB2X1 U29 ( .B0(PCcur[0]), .B1(n36), .A0N(n33), .A1N(n45), .Y(n46) );
  NAND2X2 U30 ( .A(n50), .B(n49), .Y(PCnext[1]) );
  NAND3BX4 U31 ( .AN(n87), .B(n85), .C(n86), .Y(PCnext[10]) );
  AOI222X1 U32 ( .A0(JumpRegAddr[3]), .A1(n38), .B0(targetAddr[1]), .B1(n32), 
        .C0(ADDresult[3]), .C1(n178), .Y(n58) );
  NAND2X2 U33 ( .A(n158), .B(n33), .Y(n174) );
  INVX8 U34 ( .A(ADDresult[12]), .Y(n95) );
  INVX6 U35 ( .A(ADDresult[14]), .Y(n103) );
  AOI2BB2X4 U36 ( .B0(n25), .B1(n17), .A0N(ADDresult[28]), .A1N(n162), .Y(
        PCnext[28]) );
  INVX6 U37 ( .A(ADDresult[13]), .Y(n99) );
  INVX8 U38 ( .A(n157), .Y(n35) );
  INVX20 U39 ( .A(n29), .Y(n152) );
  MX2X6 U40 ( .A(PCplus4_regD[15]), .B(PCplus4[15]), .S0(n12), .Y(
        PCplus4_actual[15]) );
  AOI2BB2X4 U41 ( .B0(n25), .B1(n26), .A0N(ADDresult[24]), .A1N(n142), .Y(
        PCnext[24]) );
  AOI222XL U42 ( .A0(PCplus4_regD[21]), .A1(n152), .B0(targetAddr[19]), .B1(
        n31), .C0(JumpRegAddr[21]), .C1(n39), .Y(n131) );
  MX2X8 U43 ( .A(branchOffset_regD[14]), .B(branchOffset_I[14]), .S0(n30), .Y(
        branchOffset_actual[16]) );
  MX2X8 U44 ( .A(PCplus4_regD[16]), .B(PCplus4[16]), .S0(n30), .Y(
        PCplus4_actual[16]) );
  NAND3X8 U45 ( .A(n9), .B(n11), .C(n53), .Y(n10) );
  INVX6 U46 ( .A(n42), .Y(n13) );
  NAND2X6 U47 ( .A(branchOffset_regD[4]), .B(n6), .Y(n7) );
  AOI2BB2X2 U48 ( .B0(PCcur[8]), .B1(n37), .A0N(n29), .A1N(n77), .Y(n79) );
  AOI2BB2XL U49 ( .B0(PCcur[1]), .B1(n37), .A0N(n34), .A1N(n48), .Y(n49) );
  AND2X2 U50 ( .A(n131), .B(n130), .Y(n5) );
  AOI2BB2XL U51 ( .B0(PCcur[21]), .B1(n36), .A0N(n34), .A1N(n129), .Y(n130) );
  AND2X2 U52 ( .A(n138), .B(n137), .Y(n2) );
  AOI2BB2XL U53 ( .B0(PCcur[16]), .B1(n37), .A0N(n34), .A1N(n108), .Y(n109) );
  AOI2BB2XL U54 ( .B0(PCcur[18]), .B1(n37), .A0N(n34), .A1N(n117), .Y(n118) );
  AOI2BB2XL U55 ( .B0(PCcur[19]), .B1(n36), .A0N(n34), .A1N(n121), .Y(n122) );
  AOI2BB2X1 U56 ( .B0(PCcur[5]), .B1(n37), .A0N(n29), .A1N(n65), .Y(n67) );
  NAND2X4 U57 ( .A(n15), .B(n28), .Y(n116) );
  INVX6 U58 ( .A(n14), .Y(n15) );
  NAND3BX4 U59 ( .AN(n13), .B(n28), .C(n52), .Y(n157) );
  NAND3BX4 U60 ( .AN(n27), .B(n13), .C(n52), .Y(n44) );
  MX2X8 U61 ( .A(branchOffset_regD[1]), .B(branchOffset_I[1]), .S0(n41), .Y(
        branchOffset_actual[3]) );
  CLKMX2X8 U62 ( .A(PCplus4_regD[20]), .B(PCplus4[20]), .S0(n12), .Y(
        PCplus4_actual[20]) );
  BUFX12 U63 ( .A(PCsrc[2]), .Y(n9) );
  CLKINVX6 U64 ( .A(n12), .Y(n6) );
  NAND2X4 U65 ( .A(branchOffset_I[4]), .B(n12), .Y(n8) );
  NAND2X8 U66 ( .A(n7), .B(n8), .Y(branchOffset_actual[6]) );
  AOI222X1 U67 ( .A0(PCplus4_regD[0]), .A1(n152), .B0(ADDresult[0]), .B1(n178), 
        .C0(JumpRegAddr[0]), .C1(n38), .Y(n47) );
  CLKMX2X4 U68 ( .A(PCplus4_regD[14]), .B(PCplus4[14]), .S0(n12), .Y(
        PCplus4_actual[14]) );
  INVX8 U69 ( .A(PCsrc[1]), .Y(n53) );
  AOI222X1 U70 ( .A0(PCplus4_regD[17]), .A1(n152), .B0(targetAddr[15]), .B1(
        n31), .C0(JumpRegAddr[17]), .C1(n39), .Y(n114) );
  BUFX20 U71 ( .A(n173), .Y(n39) );
  CLKINVX8 U72 ( .A(PCsrc[0]), .Y(n11) );
  MX2X8 U73 ( .A(PCplus4_regD[12]), .B(PCplus4[12]), .S0(n12), .Y(
        PCplus4_actual[12]) );
  AND3X8 U74 ( .A(n9), .B(n11), .C(n53), .Y(n40) );
  OAI2BB1X4 U75 ( .A0N(ADDresult[21]), .A1N(n178), .B0(n5), .Y(PCnext[21]) );
  OAI2BB1X4 U76 ( .A0N(ADDresult[23]), .A1N(n178), .B0(n2), .Y(PCnext[23]) );
  CLKMX2X4 U77 ( .A(PCplus4_regD[11]), .B(PCplus4[11]), .S0(n1), .Y(
        PCplus4_actual[11]) );
  CLKMX2X4 U78 ( .A(branchOffset_regD[9]), .B(branchOffset_I[9]), .S0(n1), .Y(
        branchOffset_actual[11]) );
  INVX8 U79 ( .A(n15), .Y(n52) );
  NAND3BX2 U80 ( .AN(n28), .B(n15), .C(n42), .Y(n43) );
  OAI211X1 U81 ( .A0(n33), .A1(n64), .B0(n63), .C0(n62), .Y(PCnext[4]) );
  INVX6 U82 ( .A(ADDresult[11]), .Y(n91) );
  INVX6 U83 ( .A(n27), .Y(n28) );
  MX2X8 U84 ( .A(branchOffset_regD[2]), .B(branchOffset_I[2]), .S0(n41), .Y(
        branchOffset_actual[4]) );
  AOI22X1 U85 ( .A0(n174), .A1(PCplus4[29]), .B0(JumpRegAddr[29]), .B1(n38), 
        .Y(n163) );
  AOI222X1 U86 ( .A0(JumpRegAddr[4]), .A1(n38), .B0(targetAddr[2]), .B1(n32), 
        .C0(ADDresult[4]), .C1(n178), .Y(n62) );
  MX2X8 U87 ( .A(PCplus4_regD[4]), .B(PCplus4[4]), .S0(n41), .Y(
        PCplus4_actual[4]) );
  MX2X8 U88 ( .A(branchOffset_regD[13]), .B(branchOffset_I[13]), .S0(n12), .Y(
        branchOffset_actual[15]) );
  AOI2BB2X1 U89 ( .B0(PCcur[2]), .B1(n37), .A0N(n29), .A1N(n51), .Y(n55) );
  OAI211X2 U90 ( .A0(n33), .A1(n56), .B0(n54), .C0(n55), .Y(PCnext[2]) );
  INVX4 U91 ( .A(n44), .Y(n171) );
  OAI211X2 U92 ( .A0(n103), .A1(n116), .B0(n102), .C0(n101), .Y(PCnext[14]) );
  NAND2X2 U93 ( .A(n47), .B(n46), .Y(PCnext[0]) );
  NAND3BX4 U94 ( .AN(n13), .B(n27), .C(n52), .Y(n172) );
  BUFX20 U95 ( .A(n172), .Y(n29) );
  NAND2BX4 U96 ( .AN(n29), .B(PCplus4_regD[29]), .Y(n164) );
  NAND2BX4 U97 ( .AN(n29), .B(PCplus4_regD[30]), .Y(n168) );
  NAND2BX4 U98 ( .AN(n29), .B(PCplus4_regD[28]), .Y(n160) );
  NAND2BX4 U99 ( .AN(n29), .B(PCplus4_regD[31]), .Y(n176) );
  AOI2BB2X1 U100 ( .B0(PCcur[6]), .B1(n37), .A0N(n29), .A1N(n69), .Y(n71) );
  OA22X4 U101 ( .A0(n178), .A1(n156), .B0(ADDresult[27]), .B1(n156), .Y(
        PCnext[27]) );
  INVX6 U102 ( .A(n178), .Y(n25) );
  NAND2X2 U103 ( .A(n155), .B(n154), .Y(n156) );
  OA22X4 U104 ( .A0(n178), .A1(n124), .B0(ADDresult[19]), .B1(n124), .Y(
        PCnext[19]) );
  NAND2X4 U105 ( .A(n123), .B(n122), .Y(n124) );
  AOI2BB2X4 U106 ( .B0(PCcur[25]), .B1(n36), .A0N(n34), .A1N(n143), .Y(n144)
         );
  AOI2BB2X4 U107 ( .B0(PCcur[22]), .B1(n36), .A0N(n34), .A1N(n132), .Y(n133)
         );
  AOI2BB2X4 U108 ( .B0(PCcur[20]), .B1(n36), .A0N(n34), .A1N(n125), .Y(n126)
         );
  INVX20 U109 ( .A(n35), .Y(n34) );
  AOI222X2 U110 ( .A0(JumpRegAddr[5]), .A1(n38), .B0(targetAddr[3]), .B1(n32), 
        .C0(ADDresult[5]), .C1(n178), .Y(n66) );
  AOI222X4 U111 ( .A0(JumpRegAddr[2]), .A1(n38), .B0(targetAddr[0]), .B1(n31), 
        .C0(ADDresult[2]), .C1(n178), .Y(n54) );
  CLKMX2X6 U112 ( .A(branchOffset_regD[7]), .B(branchOffset_I[7]), .S0(n12), 
        .Y(branchOffset_actual[9]) );
  BUFX20 U113 ( .A(n171), .Y(n36) );
  CLKMX2X4 U114 ( .A(branchOffset_regD[5]), .B(branchOffset_I[5]), .S0(n1), 
        .Y(branchOffset_actual[7]) );
  CLKMX2X4 U115 ( .A(branchOffset_regD[0]), .B(branchOffset_I[0]), .S0(n41), 
        .Y(branchOffset_actual[2]) );
  CLKMX2X4 U116 ( .A(PCplus4_regD[2]), .B(PCplus4[2]), .S0(n41), .Y(
        PCplus4_actual[2]) );
  AOI2BB2X4 U117 ( .B0(n25), .B1(n20), .A0N(ADDresult[29]), .A1N(n166), .Y(
        PCnext[29]) );
  AOI2BB2X4 U118 ( .B0(n25), .B1(n19), .A0N(ADDresult[26]), .A1N(n150), .Y(
        PCnext[26]) );
  INVX6 U119 ( .A(ADDresult[16]), .Y(n111) );
  INVX6 U120 ( .A(ADDresult[17]), .Y(n115) );
  INVX8 U121 ( .A(n158), .Y(n151) );
  NAND3X2 U122 ( .A(n177), .B(n176), .C(n175), .Y(n179) );
  CLKBUFX20 U123 ( .A(n40), .Y(n12) );
  NAND2X1 U124 ( .A(n149), .B(n148), .Y(n150) );
  AOI222X4 U125 ( .A0(PCplus4_regD[26]), .A1(n152), .B0(targetAddr[24]), .B1(
        n31), .C0(JumpRegAddr[26]), .C1(n39), .Y(n149) );
  CLKINVX1 U126 ( .A(n150), .Y(n19) );
  INVX3 U127 ( .A(n179), .Y(n18) );
  AOI222X4 U128 ( .A0(PCplus4_regD[23]), .A1(n152), .B0(targetAddr[21]), .B1(
        n31), .C0(JumpRegAddr[23]), .C1(n39), .Y(n138) );
  INVX6 U129 ( .A(ADDresult[15]), .Y(n107) );
  OA22X4 U130 ( .A0(ADDresult[18]), .A1(n120), .B0(n178), .B1(n120), .Y(
        PCnext[18]) );
  AOI2BB2X4 U131 ( .B0(n25), .B1(n23), .A0N(ADDresult[20]), .A1N(n128), .Y(
        PCnext[20]) );
  AOI2BB2X4 U132 ( .B0(n25), .B1(n22), .A0N(ADDresult[25]), .A1N(n146), .Y(
        PCnext[25]) );
  CLKMX2X4 U133 ( .A(PCplus4_regD[10]), .B(PCplus4[10]), .S0(n1), .Y(
        PCplus4_actual[10]) );
  CLKMX2X6 U134 ( .A(branchOffset_regD[12]), .B(branchOffset_I[12]), .S0(n30), 
        .Y(branchOffset_actual[14]) );
  AOI222X4 U135 ( .A0(PCplus4_regD[25]), .A1(n152), .B0(targetAddr[23]), .B1(
        n31), .C0(JumpRegAddr[25]), .C1(n39), .Y(n145) );
  AOI222X4 U136 ( .A0(PCplus4_regD[22]), .A1(n152), .B0(targetAddr[20]), .B1(
        n31), .C0(JumpRegAddr[22]), .C1(n39), .Y(n134) );
  OAI211X2 U137 ( .A0(n33), .A1(n84), .B0(n83), .C0(n82), .Y(PCnext[9]) );
  CLKMX2X6 U138 ( .A(PCplus4_regD[9]), .B(PCplus4[9]), .S0(n12), .Y(
        PCplus4_actual[9]) );
  BUFX20 U139 ( .A(n171), .Y(n37) );
  AOI2BB2X4 U140 ( .B0(n25), .B1(n24), .A0N(ADDresult[22]), .A1N(n135), .Y(
        PCnext[22]) );
  OA21X2 U141 ( .A0(n33), .A1(n80), .B0(n79), .Y(n16) );
  AOI2BB2X1 U142 ( .B0(PCcur[23]), .B1(n37), .A0N(n33), .A1N(n136), .Y(n137)
         );
  AOI222X1 U143 ( .A0(PCplus4_regD[24]), .A1(n152), .B0(targetAddr[22]), .B1(
        n31), .C0(JumpRegAddr[24]), .C1(n39), .Y(n141) );
  BUFX20 U144 ( .A(n151), .Y(n31) );
  CLKMX2X6 U145 ( .A(branchOffset_regD[6]), .B(branchOffset_I[6]), .S0(n12), 
        .Y(branchOffset_actual[8]) );
  CLKINVX2 U146 ( .A(n142), .Y(n26) );
  CLKMX2X6 U147 ( .A(branchOffset_regD[11]), .B(branchOffset_I[11]), .S0(n30), 
        .Y(branchOffset_actual[13]) );
  AOI222X4 U148 ( .A0(PCplus4_regD[19]), .A1(n152), .B0(targetAddr[17]), .B1(
        n31), .C0(JumpRegAddr[19]), .C1(n39), .Y(n123) );
  CLKMX2X6 U149 ( .A(PCplus4_regD[26]), .B(PCplus4[26]), .S0(n30), .Y(
        PCplus4_actual[26]) );
  NAND2X2 U150 ( .A(n141), .B(n140), .Y(n142) );
  AOI222X4 U151 ( .A0(PCplus4_regD[20]), .A1(n152), .B0(targetAddr[18]), .B1(
        n31), .C0(JumpRegAddr[20]), .C1(n39), .Y(n127) );
  AOI2BB2X4 U152 ( .B0(n25), .B1(n21), .A0N(ADDresult[30]), .A1N(n170), .Y(
        PCnext[30]) );
  MX2X6 U153 ( .A(branchOffset_regD[15]), .B(branchOffset_I[15]), .S0(n30), 
        .Y(branchOffset_actual[17]) );
  NAND2X2 U154 ( .A(n78), .B(n16), .Y(PCnext[8]) );
  AOI222X2 U155 ( .A0(JumpRegAddr[8]), .A1(n38), .B0(targetAddr[6]), .B1(n32), 
        .C0(ADDresult[8]), .C1(n178), .Y(n78) );
  CLKMX2X4 U156 ( .A(branchOffset_regD[8]), .B(branchOffset_I[8]), .S0(n1), 
        .Y(branchOffset_actual[10]) );
  CLKMX2X6 U157 ( .A(PCplus4_regD[8]), .B(PCplus4[8]), .S0(n12), .Y(
        PCplus4_actual[8]) );
  AOI222X4 U158 ( .A0(PCplus4_regD[18]), .A1(n152), .B0(targetAddr[16]), .B1(
        n31), .C0(JumpRegAddr[18]), .C1(n39), .Y(n119) );
  INVX20 U159 ( .A(n35), .Y(n33) );
  BUFX20 U160 ( .A(n151), .Y(n32) );
  CLKBUFX20 U161 ( .A(n40), .Y(n30) );
  AOI2BB2X4 U162 ( .B0(n25), .B1(n18), .A0N(ADDresult[31]), .A1N(n179), .Y(
        PCnext[31]) );
  AOI22X1 U163 ( .A0(n174), .A1(PCplus4[28]), .B0(JumpRegAddr[28]), .B1(n38), 
        .Y(n159) );
  CLKMX2X8 U164 ( .A(PCplus4_regD[28]), .B(PCplus4[28]), .S0(n30), .Y(
        PCplus4_actual[28]) );
  AOI22X1 U165 ( .A0(n174), .A1(PCplus4[30]), .B0(JumpRegAddr[30]), .B1(n38), 
        .Y(n167) );
  CLKMX2X8 U166 ( .A(PCplus4_regD[19]), .B(PCplus4[19]), .S0(n30), .Y(
        PCplus4_actual[19]) );
  AOI2BB2XL U167 ( .B0(PCcur[4]), .B1(n37), .A0N(n29), .A1N(n61), .Y(n63) );
  AOI2BB2XL U168 ( .B0(PCcur[3]), .B1(n37), .A0N(n29), .A1N(n57), .Y(n59) );
  OAI211X2 U169 ( .A0(n116), .A1(n95), .B0(n94), .C0(n93), .Y(PCnext[12]) );
  INVXL U170 ( .A(PCplus4[18]), .Y(n117) );
  INVXL U171 ( .A(PCplus4[17]), .Y(n112) );
  INVXL U172 ( .A(PCplus4[15]), .Y(n104) );
  INVXL U173 ( .A(PCplus4[16]), .Y(n108) );
  INVXL U174 ( .A(PCplus4[14]), .Y(n100) );
  INVXL U175 ( .A(PCplus4[12]), .Y(n92) );
  INVX1 U176 ( .A(PCplus4[13]), .Y(n96) );
  INVXL U177 ( .A(PCplus4[11]), .Y(n88) );
  AOI222XL U178 ( .A0(PCplus4_regD[12]), .A1(n152), .B0(targetAddr[10]), .B1(
        n32), .C0(JumpRegAddr[12]), .C1(n39), .Y(n94) );
  AOI222XL U179 ( .A0(PCplus4_regD[15]), .A1(n152), .B0(targetAddr[13]), .B1(
        n32), .C0(JumpRegAddr[15]), .C1(n39), .Y(n106) );
  AOI222XL U180 ( .A0(PCplus4_regD[11]), .A1(n152), .B0(targetAddr[9]), .B1(
        n32), .C0(JumpRegAddr[11]), .C1(n39), .Y(n90) );
  AOI222XL U181 ( .A0(PCplus4_regD[14]), .A1(n152), .B0(targetAddr[12]), .B1(
        n32), .C0(JumpRegAddr[14]), .C1(n39), .Y(n102) );
  CLKMX2X4 U182 ( .A(PCplus4_regD[24]), .B(PCplus4[24]), .S0(n30), .Y(
        PCplus4_actual[24]) );
  CLKMX2X4 U183 ( .A(PCplus4_regD[22]), .B(PCplus4[22]), .S0(n30), .Y(
        PCplus4_actual[22]) );
  CLKMX2X4 U184 ( .A(PCplus4_regD[21]), .B(PCplus4[21]), .S0(n30), .Y(
        PCplus4_actual[21]) );
  CLKMX2X4 U185 ( .A(PCplus4_regD[25]), .B(PCplus4[25]), .S0(n30), .Y(
        PCplus4_actual[25]) );
  CLKMX2X4 U186 ( .A(PCplus4_regD[23]), .B(PCplus4[23]), .S0(n30), .Y(
        PCplus4_actual[23]) );
  CLKMX2X4 U187 ( .A(PCplus4_regD[30]), .B(PCplus4[30]), .S0(n30), .Y(
        PCplus4_actual[30]) );
  CLKMX2X4 U188 ( .A(PCplus4_regD[29]), .B(PCplus4[29]), .S0(n30), .Y(
        PCplus4_actual[29]) );
  CLKMX2X4 U189 ( .A(PCplus4_regD[18]), .B(PCplus4[18]), .S0(n30), .Y(
        PCplus4_actual[18]) );
  AOI222XL U190 ( .A0(PCplus4_regD[13]), .A1(n152), .B0(targetAddr[11]), .B1(
        n32), .C0(JumpRegAddr[13]), .C1(n39), .Y(n98) );
  INVXL U191 ( .A(PCplus4[3]), .Y(n60) );
  AOI2BB2XL U192 ( .B0(PCcur[24]), .B1(n36), .A0N(n33), .A1N(n139), .Y(n140)
         );
  INVXL U193 ( .A(PCplus4[24]), .Y(n139) );
  INVXL U194 ( .A(PCplus4[22]), .Y(n132) );
  INVXL U195 ( .A(PCplus4[19]), .Y(n121) );
  INVXL U196 ( .A(PCplus4[21]), .Y(n129) );
  INVXL U197 ( .A(PCplus4[25]), .Y(n143) );
  INVXL U198 ( .A(PCplus4[23]), .Y(n136) );
  INVXL U199 ( .A(PCplus4[2]), .Y(n56) );
  MX2XL U200 ( .A(PCplus4_regD[31]), .B(PCplus4[31]), .S0(n30), .Y(
        PCplus4_actual[31]) );
  CLKMX2X4 U201 ( .A(PCplus4_regD[27]), .B(PCplus4[27]), .S0(n30), .Y(
        PCplus4_actual[27]) );
  INVXL U202 ( .A(PCplus4_regD[8]), .Y(n77) );
  NAND2XL U203 ( .A(PCcur[29]), .B(n36), .Y(n165) );
  NAND2XL U204 ( .A(PCcur[30]), .B(n36), .Y(n169) );
  INVXL U205 ( .A(PCplus4_regD[2]), .Y(n51) );
  INVXL U206 ( .A(PCplus4_regD[3]), .Y(n57) );
  INVXL U207 ( .A(PCplus4_regD[4]), .Y(n61) );
  INVXL U208 ( .A(PCplus4_regD[5]), .Y(n65) );
  INVXL U209 ( .A(PCplus4_regD[9]), .Y(n81) );
  INVXL U210 ( .A(PCplus4_regD[7]), .Y(n73) );
  INVXL U211 ( .A(PCplus4_regD[6]), .Y(n69) );
  CLKINVX1 U212 ( .A(n135), .Y(n24) );
  NAND2X1 U213 ( .A(n134), .B(n133), .Y(n135) );
  CLKINVX1 U214 ( .A(n128), .Y(n23) );
  NAND2X1 U215 ( .A(n127), .B(n126), .Y(n128) );
  CLKINVX1 U216 ( .A(n146), .Y(n22) );
  NAND2X1 U217 ( .A(n145), .B(n144), .Y(n146) );
  INVX1 U218 ( .A(n162), .Y(n17) );
  NAND3X1 U219 ( .A(n161), .B(n160), .C(n159), .Y(n162) );
  INVX1 U220 ( .A(n170), .Y(n21) );
  NAND3X1 U221 ( .A(n169), .B(n168), .C(n167), .Y(n170) );
  CLKINVX1 U222 ( .A(PCplus4[1]), .Y(n48) );
  AOI2BB2XL U223 ( .B0(PCcur[14]), .B1(n37), .A0N(n34), .A1N(n100), .Y(n101)
         );
  AOI2BB2XL U224 ( .B0(PCcur[15]), .B1(n37), .A0N(n34), .A1N(n104), .Y(n105)
         );
  AOI2BB2XL U225 ( .B0(PCcur[13]), .B1(n37), .A0N(n34), .A1N(n96), .Y(n97) );
  AOI2BB2XL U226 ( .B0(PCcur[17]), .B1(n37), .A0N(n34), .A1N(n112), .Y(n113)
         );
  AOI2BB2XL U227 ( .B0(PCcur[11]), .B1(n37), .A0N(n34), .A1N(n88), .Y(n89) );
  INVXL U228 ( .A(PCplus4[20]), .Y(n125) );
  AOI2BB2X1 U229 ( .B0(PCcur[27]), .B1(n36), .A0N(n33), .A1N(n153), .Y(n154)
         );
  INVX1 U230 ( .A(PCplus4[27]), .Y(n153) );
  AOI2BB2X1 U231 ( .B0(PCcur[26]), .B1(n36), .A0N(n33), .A1N(n147), .Y(n148)
         );
  INVX1 U232 ( .A(PCplus4[26]), .Y(n147) );
  CLKINVX1 U233 ( .A(PCplus4[7]), .Y(n76) );
  CLKINVX1 U234 ( .A(PCplus4[9]), .Y(n84) );
  INVXL U235 ( .A(PCplus4[4]), .Y(n64) );
  INVXL U236 ( .A(PCplus4[5]), .Y(n68) );
  CLKINVX1 U237 ( .A(PCplus4[6]), .Y(n72) );
  MX2XL U238 ( .A(PCplus4_regD[1]), .B(PCplus4[1]), .S0(n30), .Y(
        PCplus4_actual[1]) );
  AO22X1 U239 ( .A0(targetAddr[8]), .A1(n32), .B0(JumpRegAddr[10]), .B1(n38), 
        .Y(n87) );
  AOI222XL U240 ( .A0(PCplus4[10]), .A1(n35), .B0(PCplus4_regD[10]), .B1(n152), 
        .C0(PCcur[10]), .C1(n36), .Y(n86) );
  CLKINVX1 U241 ( .A(PCplus4[0]), .Y(n45) );
  NAND2X1 U242 ( .A(n119), .B(n118), .Y(n120) );
  AOI2BB2XL U243 ( .B0(PCcur[12]), .B1(n37), .A0N(n34), .A1N(n92), .Y(n93) );
  CLKINVX1 U244 ( .A(PCplus4[8]), .Y(n80) );
  NAND2X1 U245 ( .A(PCcur[31]), .B(n36), .Y(n177) );
  NAND2X1 U246 ( .A(PCcur[28]), .B(n36), .Y(n161) );
  OAI211X2 U247 ( .A0(n33), .A1(n60), .B0(n59), .C0(n58), .Y(PCnext[3]) );
  OAI211X2 U248 ( .A0(n33), .A1(n68), .B0(n67), .C0(n66), .Y(PCnext[5]) );
  AOI222X2 U249 ( .A0(JumpRegAddr[6]), .A1(n38), .B0(targetAddr[4]), .B1(n32), 
        .C0(ADDresult[6]), .C1(n178), .Y(n70) );
  OAI211X2 U250 ( .A0(n33), .A1(n72), .B0(n71), .C0(n70), .Y(PCnext[6]) );
  AOI2BB2X2 U251 ( .B0(PCcur[7]), .B1(n37), .A0N(n29), .A1N(n73), .Y(n75) );
  AOI222X2 U252 ( .A0(JumpRegAddr[7]), .A1(n38), .B0(targetAddr[5]), .B1(n32), 
        .C0(ADDresult[7]), .C1(n178), .Y(n74) );
  OAI211X2 U253 ( .A0(n33), .A1(n76), .B0(n75), .C0(n74), .Y(PCnext[7]) );
  AOI2BB2X2 U254 ( .B0(PCcur[9]), .B1(n37), .A0N(n29), .A1N(n81), .Y(n83) );
  AOI222X2 U255 ( .A0(JumpRegAddr[9]), .A1(n38), .B0(targetAddr[7]), .B1(n32), 
        .C0(ADDresult[9]), .C1(n178), .Y(n82) );
  OAI211X2 U256 ( .A0(n91), .A1(n116), .B0(n90), .C0(n89), .Y(PCnext[11]) );
  OAI211X2 U257 ( .A0(n99), .A1(n116), .B0(n98), .C0(n97), .Y(PCnext[13]) );
  OAI211X2 U258 ( .A0(n107), .A1(n116), .B0(n106), .C0(n105), .Y(PCnext[15])
         );
  OAI211X2 U259 ( .A0(n111), .A1(n116), .B0(n110), .C0(n109), .Y(PCnext[16])
         );
  OAI211X2 U260 ( .A0(n115), .A1(n116), .B0(n114), .C0(n113), .Y(PCnext[17])
         );
endmodule


module PCsrcLogic ( pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, 
        predict, stallcache, stall_lw_use, PCsrc );
  output [2:0] PCsrc;
  input pred_cond, Branch_EX, Branch_IF, equal, Jump, JumpReg, predict,
         stallcache, stall_lw_use;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INVX4 U3 ( .A(equal), .Y(n9) );
  AND2X6 U4 ( .A(pred_cond), .B(Branch_EX), .Y(n2) );
  INVX3 U5 ( .A(JumpReg), .Y(n3) );
  OAI2BB1X4 U6 ( .A0N(n7), .A1N(n8), .B0(n1), .Y(PCsrc[0]) );
  CLKINVX1 U7 ( .A(n12), .Y(n1) );
  AND2X8 U8 ( .A(pred_cond), .B(Branch_EX), .Y(n6) );
  AND3X8 U9 ( .A(Branch_IF), .B(predict), .C(n10), .Y(n11) );
  INVX8 U10 ( .A(Jump), .Y(n10) );
  AOI21X4 U11 ( .A0(n4), .A1(n3), .B0(n12), .Y(PCsrc[1]) );
  MXI2X4 U12 ( .A(Jump), .B(n9), .S0(n2), .Y(n4) );
  AOI21X4 U13 ( .A0(n5), .A1(n3), .B0(n12), .Y(PCsrc[2]) );
  MXI2X4 U14 ( .A(n11), .B(equal), .S0(n6), .Y(n5) );
  OR2X8 U15 ( .A(stallcache), .B(stall_lw_use), .Y(n12) );
  MXI2X4 U16 ( .A(n10), .B(n9), .S0(n6), .Y(n8) );
  INVXL U17 ( .A(JumpReg), .Y(n7) );
endmodule


module ALU_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ALU_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n10, n11, n12, n14, n16, n19, n20, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n89, n91, n92, n93, n94, n99, n100, n102, n103, n105, n106, n107,
         n108, n109, n110, n113, n114, n115, n116, n117, n118, n120, n121,
         n122, n123, n124, n127, n128, n129, n130, n131, n132, n137, n138,
         n139, n140, n141, n143, n145, n146, n147, n148, n149, n150, n153,
         n154, n155, n156, n157, n158, n159, n161, n162, n163, n164, n165,
         n167, n168, n173, n174, n175, n176, n177, n179, n181, n182, n183,
         n184, n185, n186, n187, n188, n190, n191, n192, n195, n196, n197,
         n198, n199, n200, n202, n205, n206, n208, n209, n211, n212, n213,
         n214, n215, n216, n217, n221, n222, n223, n224, n225, n226, n227,
         n229, n230, n231, n232, n233, n235, n236, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n255, n256,
         n257, n260, n261, n262, n263, n265, n269, n273, n274, n276, n277,
         n278, n279, n280, n282, n283, n285, n286, n287, n288, n289, n292,
         n293, n294, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n309, n310, n311, n312, n313, n315, n317, n318, n319,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484;

  AOI21X4 U57 ( .A0(n94), .A1(n77), .B0(n78), .Y(n5) );
  AOI21X4 U107 ( .A0(n132), .A1(n115), .B0(n116), .Y(n114) );
  AOI21X4 U157 ( .A0(n168), .A1(n153), .B0(n154), .Y(n148) );
  AOI21X4 U199 ( .A0(n183), .A1(n200), .B0(n184), .Y(n182) );
  AOI21X4 U290 ( .A0(n263), .A1(n250), .B0(n251), .Y(n249) );
  AOI21X4 U329 ( .A0(n277), .A1(n285), .B0(n278), .Y(n276) );
  OAI21X2 U357 ( .A0(n434), .A1(n57), .B0(n58), .Y(n56) );
  INVX12 U358 ( .A(n480), .Y(n483) );
  CLKINVX6 U359 ( .A(n76), .Y(n434) );
  AOI2BB1X4 U360 ( .A0N(n246), .A1N(n188), .B0(n425), .Y(n424) );
  CLKINVX20 U361 ( .A(n424), .Y(n187) );
  AO21X4 U362 ( .A0(n428), .A1(n190), .B0(n191), .Y(n425) );
  INVX3 U363 ( .A(n150), .Y(n426) );
  NAND2X8 U364 ( .A(B[21]), .B(A[21]), .Y(n138) );
  NOR2X8 U365 ( .A(B[5]), .B(A[5]), .Y(n452) );
  AND2XL U366 ( .A(B[4]), .B(A[4]), .Y(n458) );
  NOR2X8 U367 ( .A(B[13]), .B(A[13]), .Y(n205) );
  OR2XL U368 ( .A(B[13]), .B(A[13]), .Y(n427) );
  NAND2X4 U369 ( .A(B[6]), .B(A[6]), .Y(n260) );
  NAND2X4 U370 ( .A(B[20]), .B(A[20]), .Y(n145) );
  NOR2X6 U371 ( .A(B[28]), .B(A[28]), .Y(n68) );
  NOR2X1 U372 ( .A(n484), .B(A[0]), .Y(n288) );
  NAND2X6 U373 ( .A(n484), .B(A[0]), .Y(n289) );
  CLKINVX3 U374 ( .A(n124), .Y(n299) );
  OAI21X1 U375 ( .A0(n435), .A1(n124), .B0(n127), .Y(n123) );
  NOR2BX2 U376 ( .AN(n131), .B(n124), .Y(n122) );
  OAI21X2 U377 ( .A0(n434), .A1(n46), .B0(n47), .Y(n45) );
  NAND2X2 U378 ( .A(B[30]), .B(A[30]), .Y(n51) );
  NAND2X2 U379 ( .A(n262), .B(n250), .Y(n248) );
  OR2X6 U380 ( .A(n205), .B(n213), .Y(n466) );
  NAND2X8 U381 ( .A(B[12]), .B(A[12]), .Y(n213) );
  NOR2X6 U382 ( .A(B[1]), .B(A[1]), .Y(n286) );
  NOR2X6 U383 ( .A(n212), .B(n205), .Y(n199) );
  NOR2X8 U384 ( .A(n117), .B(n124), .Y(n115) );
  NAND2X6 U385 ( .A(n471), .B(n426), .Y(n146) );
  NOR2X8 U386 ( .A(n185), .B(n192), .Y(n183) );
  NOR2X8 U387 ( .A(B[10]), .B(A[10]), .Y(n230) );
  NAND2X4 U388 ( .A(B[9]), .B(A[9]), .Y(n242) );
  INVX20 U389 ( .A(n477), .Y(n2) );
  NOR2X6 U390 ( .A(n230), .B(n223), .Y(n221) );
  AOI21X2 U391 ( .A0(n236), .A1(n221), .B0(n222), .Y(n216) );
  NAND2X4 U392 ( .A(n115), .B(n131), .Y(n113) );
  INVX1 U393 ( .A(n200), .Y(n202) );
  OR2X4 U394 ( .A(n246), .B(n233), .Y(n467) );
  AOI21X1 U395 ( .A0(n428), .A1(n309), .B0(n211), .Y(n209) );
  NOR2X6 U396 ( .A(B[15]), .B(A[15]), .Y(n185) );
  NAND2X2 U397 ( .A(n465), .B(n429), .Y(n67) );
  AND2X1 U398 ( .A(n300), .B(n138), .Y(n453) );
  XOR2X1 U399 ( .A(n473), .B(n474), .Y(SUM[5]) );
  NAND2X2 U400 ( .A(n454), .B(n269), .Y(n474) );
  NAND2X2 U401 ( .A(n312), .B(n242), .Y(n29) );
  INVX4 U402 ( .A(n5), .Y(n76) );
  INVX6 U403 ( .A(n430), .Y(n301) );
  NAND2X2 U404 ( .A(n293), .B(n429), .Y(n10) );
  CLKINVX1 U405 ( .A(n443), .Y(n130) );
  CLKAND2X3 U406 ( .A(n292), .B(n62), .Y(n445) );
  AO21X4 U407 ( .A0(n438), .A1(n221), .B0(n222), .Y(n428) );
  NAND2X6 U408 ( .A(B[28]), .B(A[28]), .Y(n429) );
  NOR2X8 U409 ( .A(B[20]), .B(A[20]), .Y(n430) );
  AND2X4 U410 ( .A(n301), .B(n145), .Y(n431) );
  CLKAND2X8 U411 ( .A(n304), .B(n174), .Y(n432) );
  NOR2X8 U412 ( .A(n468), .B(n105), .Y(n103) );
  OAI21XL U413 ( .A0(n202), .A1(n192), .B0(n195), .Y(n191) );
  NOR2X4 U414 ( .A(A[12]), .B(B[12]), .Y(n212) );
  NOR2X8 U415 ( .A(B[6]), .B(A[6]), .Y(n257) );
  NAND2X2 U416 ( .A(n4), .B(n84), .Y(n82) );
  NAND2X2 U417 ( .A(n4), .B(n93), .Y(n91) );
  INVX3 U418 ( .A(n4), .Y(n109) );
  NAND2X8 U419 ( .A(B[8]), .B(A[8]), .Y(n245) );
  NAND2X6 U420 ( .A(n455), .B(n103), .Y(n451) );
  INVX12 U421 ( .A(n444), .Y(n86) );
  NAND2X4 U422 ( .A(n4), .B(n66), .Y(n64) );
  OR2X2 U423 ( .A(n2), .B(n53), .Y(n463) );
  NAND2XL U424 ( .A(n427), .B(n206), .Y(n25) );
  NAND2X2 U425 ( .A(n4), .B(n55), .Y(n53) );
  NOR2X6 U426 ( .A(n252), .B(n257), .Y(n250) );
  NOR2X6 U427 ( .A(n79), .B(n86), .Y(n77) );
  INVX1 U428 ( .A(n68), .Y(n293) );
  OR2X2 U429 ( .A(n5), .B(n68), .Y(n465) );
  NOR2X8 U430 ( .A(n68), .B(n61), .Y(n59) );
  AOI21X1 U431 ( .A0(n428), .A1(n199), .B0(n200), .Y(n198) );
  NAND2X8 U432 ( .A(n466), .B(n206), .Y(n200) );
  NAND2X4 U433 ( .A(B[24]), .B(A[24]), .Y(n107) );
  NOR2X6 U434 ( .A(n137), .B(n430), .Y(n131) );
  NAND2X2 U435 ( .A(n190), .B(n217), .Y(n188) );
  OR2X8 U436 ( .A(n452), .B(n274), .Y(n464) );
  AOI21X2 U437 ( .A0(n483), .A1(n55), .B0(n56), .Y(n54) );
  INVX2 U438 ( .A(n483), .Y(n110) );
  INVXL U439 ( .A(n137), .Y(n300) );
  OAI21X2 U440 ( .A0(n246), .A1(n226), .B0(n227), .Y(n225) );
  AOI21X1 U441 ( .A0(n438), .A1(n311), .B0(n229), .Y(n227) );
  OR2X6 U442 ( .A(n2), .B(n165), .Y(n433) );
  NAND2X4 U443 ( .A(n433), .B(n436), .Y(n164) );
  INVX3 U444 ( .A(n148), .Y(n150) );
  NOR2X6 U445 ( .A(B[3]), .B(A[3]), .Y(n279) );
  NOR2X4 U446 ( .A(n215), .B(n181), .Y(n179) );
  OA21X2 U447 ( .A0(n145), .A1(n137), .B0(n138), .Y(n435) );
  OA21X2 U448 ( .A0(n286), .A1(n289), .B0(n287), .Y(n441) );
  OA21X4 U449 ( .A0(n173), .A1(n177), .B0(n174), .Y(n436) );
  NAND2X8 U450 ( .A(B[16]), .B(A[16]), .Y(n177) );
  NAND2X8 U451 ( .A(B[10]), .B(A[10]), .Y(n231) );
  NAND2X4 U452 ( .A(B[11]), .B(A[11]), .Y(n224) );
  OA21X2 U453 ( .A0(n99), .A1(n107), .B0(n100), .Y(n437) );
  NAND2X8 U454 ( .A(n93), .B(n77), .Y(n6) );
  INVX4 U455 ( .A(n282), .Y(n319) );
  NOR2X4 U456 ( .A(n282), .B(n279), .Y(n277) );
  NOR2X6 U457 ( .A(B[2]), .B(A[2]), .Y(n282) );
  NAND2X6 U458 ( .A(n199), .B(n183), .Y(n181) );
  NAND2X8 U459 ( .A(n221), .B(n235), .Y(n215) );
  OAI21X2 U460 ( .A0(n241), .A1(n245), .B0(n242), .Y(n438) );
  OAI21X2 U461 ( .A0(n279), .A1(n283), .B0(n280), .Y(n439) );
  OR2XL U462 ( .A(B[14]), .B(A[14]), .Y(n440) );
  NOR2X6 U463 ( .A(n155), .B(n162), .Y(n153) );
  NOR2X4 U464 ( .A(B[4]), .B(A[4]), .Y(n273) );
  NOR2X8 U465 ( .A(n244), .B(n241), .Y(n235) );
  NOR2X4 U466 ( .A(B[8]), .B(A[8]), .Y(n244) );
  NOR2X8 U467 ( .A(B[7]), .B(A[7]), .Y(n252) );
  XNOR2X4 U468 ( .A(n52), .B(n8), .Y(SUM[30]) );
  OAI21X1 U469 ( .A0(n2), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X2 U470 ( .A0(n2), .A1(n64), .B0(n65), .Y(n63) );
  INVX2 U471 ( .A(n60), .Y(n58) );
  XNOR2X4 U472 ( .A(n442), .B(n12), .Y(SUM[26]) );
  OAI21X2 U473 ( .A0(n2), .A1(n91), .B0(n92), .Y(n442) );
  NOR2X8 U474 ( .A(B[25]), .B(A[25]), .Y(n99) );
  OAI2BB1X4 U475 ( .A0N(n150), .A1N(n131), .B0(n435), .Y(n443) );
  NAND2X4 U476 ( .A(B[3]), .B(A[3]), .Y(n280) );
  NAND2X1 U477 ( .A(n318), .B(n280), .Y(n35) );
  OR2X8 U478 ( .A(B[26]), .B(A[26]), .Y(n444) );
  NAND2X6 U479 ( .A(B[2]), .B(A[2]), .Y(n283) );
  NOR2X6 U480 ( .A(n273), .B(n452), .Y(n262) );
  XOR2X4 U481 ( .A(n63), .B(n445), .Y(SUM[29]) );
  NAND2X4 U482 ( .A(n446), .B(n253), .Y(n31) );
  NAND2X4 U483 ( .A(B[7]), .B(A[7]), .Y(n253) );
  OR2X4 U484 ( .A(B[7]), .B(A[7]), .Y(n446) );
  OR2X2 U485 ( .A(B[30]), .B(A[30]), .Y(n481) );
  OR2X4 U486 ( .A(n2), .B(n176), .Y(n469) );
  NAND2X4 U487 ( .A(n470), .B(n43), .Y(n41) );
  NAND2X1 U488 ( .A(n149), .B(n301), .Y(n140) );
  XOR2X4 U489 ( .A(n451), .B(n447), .Y(SUM[25]) );
  CLKAND2X8 U490 ( .A(n296), .B(n100), .Y(n447) );
  XOR2X4 U491 ( .A(n479), .B(n448), .Y(SUM[23]) );
  NAND2X2 U492 ( .A(n298), .B(n118), .Y(n448) );
  XOR2X4 U493 ( .A(n146), .B(n431), .Y(SUM[20]) );
  XNOR2X4 U494 ( .A(n462), .B(n34), .Y(SUM[4]) );
  NOR2X6 U495 ( .A(B[16]), .B(A[16]), .Y(n176) );
  XOR2X2 U496 ( .A(n441), .B(n36), .Y(SUM[2]) );
  NAND2X4 U497 ( .A(B[1]), .B(A[1]), .Y(n287) );
  INVXL U498 ( .A(n428), .Y(n449) );
  AOI21X4 U499 ( .A0(n483), .A1(n84), .B0(n85), .Y(n83) );
  BUFX3 U500 ( .A(B[0]), .Y(n484) );
  XOR2X4 U501 ( .A(n472), .B(n35), .Y(SUM[3]) );
  OA21X4 U502 ( .A0(n441), .A1(n460), .B0(n283), .Y(n472) );
  NAND2X6 U503 ( .A(B[14]), .B(A[14]), .Y(n195) );
  NAND2X4 U504 ( .A(B[15]), .B(A[15]), .Y(n186) );
  CLKBUFX2 U505 ( .A(n263), .Y(n450) );
  OA21X4 U506 ( .A0(n246), .A1(n208), .B0(n209), .Y(n475) );
  OAI21X2 U507 ( .A0(n185), .A1(n195), .B0(n186), .Y(n184) );
  NAND2X2 U508 ( .A(n306), .B(n186), .Y(n23) );
  OR2X1 U509 ( .A(B[5]), .B(A[5]), .Y(n454) );
  NAND2X4 U510 ( .A(B[5]), .B(A[5]), .Y(n269) );
  INVX1 U511 ( .A(n263), .Y(n265) );
  NAND2X4 U512 ( .A(B[18]), .B(A[18]), .Y(n163) );
  NAND2X6 U513 ( .A(B[4]), .B(A[4]), .Y(n274) );
  NOR2X8 U514 ( .A(B[14]), .B(A[14]), .Y(n192) );
  NAND2X4 U515 ( .A(n463), .B(n54), .Y(n52) );
  INVX2 U516 ( .A(n273), .Y(n317) );
  NOR2BX1 U517 ( .AN(n262), .B(n257), .Y(n255) );
  XNOR2X4 U518 ( .A(n164), .B(n20), .Y(SUM[18]) );
  NAND2X4 U519 ( .A(B[17]), .B(A[17]), .Y(n174) );
  NAND2X4 U520 ( .A(n469), .B(n177), .Y(n175) );
  NOR2X8 U521 ( .A(B[17]), .B(A[17]), .Y(n173) );
  INVX3 U522 ( .A(n173), .Y(n304) );
  NOR2X6 U523 ( .A(n176), .B(n173), .Y(n167) );
  CLKINVX6 U524 ( .A(n247), .Y(n246) );
  OAI21X4 U525 ( .A0(n73), .A1(n2), .B0(n74), .Y(n72) );
  XOR2X4 U526 ( .A(n139), .B(n453), .Y(SUM[21]) );
  AND2X8 U527 ( .A(n483), .B(n297), .Y(n468) );
  AO21X4 U528 ( .A0(n462), .A1(n255), .B0(n256), .Y(n476) );
  OR2X2 U529 ( .A(n2), .B(n42), .Y(n470) );
  XNOR2X4 U530 ( .A(n157), .B(n19), .Y(SUM[19]) );
  NAND2X2 U531 ( .A(n4), .B(n297), .Y(n102) );
  OR2X4 U532 ( .A(n2), .B(n102), .Y(n455) );
  NAND2X6 U533 ( .A(n153), .B(n167), .Y(n147) );
  AOI21X2 U534 ( .A0(n150), .A1(n122), .B0(n123), .Y(n121) );
  AOI21X4 U535 ( .A0(n150), .A1(n301), .B0(n143), .Y(n141) );
  OAI21X4 U536 ( .A0(n252), .A1(n260), .B0(n253), .Y(n251) );
  OAI21X2 U537 ( .A0(n246), .A1(n244), .B0(n245), .Y(n243) );
  XNOR2X4 U538 ( .A(n243), .B(n29), .Y(SUM[9]) );
  OR2X2 U539 ( .A(n2), .B(n129), .Y(n456) );
  NAND2X4 U540 ( .A(n456), .B(n130), .Y(n128) );
  XNOR2X4 U541 ( .A(n128), .B(n16), .Y(SUM[22]) );
  OAI21X4 U542 ( .A0(n140), .A1(n2), .B0(n141), .Y(n139) );
  AOI21X4 U543 ( .A0(n483), .A1(n75), .B0(n76), .Y(n74) );
  NAND2X2 U544 ( .A(B[13]), .B(A[13]), .Y(n206) );
  OAI21X4 U545 ( .A0(n155), .A1(n163), .B0(n156), .Y(n154) );
  NAND2X6 U546 ( .A(B[19]), .B(A[19]), .Y(n156) );
  AOI21X2 U547 ( .A0(n483), .A1(n93), .B0(n94), .Y(n92) );
  NOR2X8 U548 ( .A(B[29]), .B(A[29]), .Y(n61) );
  NOR2X4 U549 ( .A(n6), .B(n57), .Y(n55) );
  INVX4 U550 ( .A(n59), .Y(n57) );
  NOR2X8 U551 ( .A(B[22]), .B(A[22]), .Y(n124) );
  INVX8 U552 ( .A(n147), .Y(n149) );
  OA21X4 U553 ( .A0(n241), .A1(n245), .B0(n242), .Y(n457) );
  AOI21X4 U554 ( .A0(n483), .A1(n66), .B0(n67), .Y(n65) );
  NAND2X4 U555 ( .A(B[22]), .B(A[22]), .Y(n127) );
  NOR2X4 U556 ( .A(n6), .B(n68), .Y(n66) );
  NAND2X2 U557 ( .A(n317), .B(n274), .Y(n34) );
  NOR2X8 U558 ( .A(B[27]), .B(A[27]), .Y(n79) );
  INVX4 U559 ( .A(n6), .Y(n75) );
  NAND2X2 U560 ( .A(n4), .B(n75), .Y(n73) );
  OAI21X1 U561 ( .A0(n437), .A1(n86), .B0(n89), .Y(n85) );
  INVX1 U562 ( .A(n257), .Y(n315) );
  OAI21X2 U563 ( .A0(n265), .A1(n257), .B0(n260), .Y(n256) );
  NAND2BX4 U564 ( .AN(n288), .B(n289), .Y(n38) );
  NAND2X8 U565 ( .A(n464), .B(n269), .Y(n263) );
  XNOR2X4 U566 ( .A(n72), .B(n10), .Y(SUM[28]) );
  OR2XL U567 ( .A(B[1]), .B(A[1]), .Y(n459) );
  INVX3 U568 ( .A(n51), .Y(n49) );
  INVX12 U569 ( .A(n215), .Y(n217) );
  OAI21X2 U570 ( .A0(n2), .A1(n82), .B0(n83), .Y(n81) );
  NOR2X8 U571 ( .A(B[19]), .B(A[19]), .Y(n155) );
  XNOR2X2 U572 ( .A(n108), .B(n14), .Y(SUM[24]) );
  INVX2 U573 ( .A(n319), .Y(n460) );
  INVXL U574 ( .A(n155), .Y(n302) );
  INVX3 U575 ( .A(n436), .Y(n461) );
  XOR2X4 U576 ( .A(n175), .B(n432), .Y(SUM[17]) );
  XNOR2X4 U577 ( .A(n476), .B(n31), .Y(SUM[7]) );
  XNOR2X4 U578 ( .A(n214), .B(n26), .Y(SUM[12]) );
  OAI21X1 U579 ( .A0(n246), .A1(n215), .B0(n449), .Y(n214) );
  NAND2X4 U580 ( .A(n59), .B(n481), .Y(n46) );
  AOI21X2 U581 ( .A0(n60), .A1(n481), .B0(n49), .Y(n47) );
  OAI21X4 U582 ( .A0(n173), .A1(n177), .B0(n174), .Y(n168) );
  OAI21X2 U583 ( .A0(n2), .A1(n158), .B0(n159), .Y(n157) );
  OAI21X4 U584 ( .A0(n145), .A1(n137), .B0(n138), .Y(n132) );
  OR2X8 U585 ( .A(n2), .B(n147), .Y(n471) );
  OAI21X2 U586 ( .A0(n117), .A1(n127), .B0(n118), .Y(n116) );
  AOI21X2 U587 ( .A0(n462), .A1(n262), .B0(n450), .Y(n261) );
  NOR2X4 U588 ( .A(n6), .B(n46), .Y(n44) );
  INVX4 U589 ( .A(n230), .Y(n311) );
  OAI21X4 U590 ( .A0(n223), .A1(n231), .B0(n224), .Y(n222) );
  OA21X4 U591 ( .A0(n216), .A1(n181), .B0(n182), .Y(n478) );
  AO21X4 U592 ( .A0(n277), .A1(n285), .B0(n439), .Y(n462) );
  OAI21X4 U593 ( .A0(n279), .A1(n283), .B0(n280), .Y(n278) );
  NAND2X2 U594 ( .A(n481), .B(n51), .Y(n8) );
  AOI21X2 U595 ( .A0(n483), .A1(n44), .B0(n45), .Y(n43) );
  XNOR2X4 U596 ( .A(n187), .B(n23), .Y(SUM[15]) );
  XNOR2X4 U597 ( .A(n81), .B(n11), .Y(SUM[27]) );
  XOR2X4 U598 ( .A(n261), .B(n32), .Y(SUM[6]) );
  OAI21X2 U599 ( .A0(n246), .A1(n197), .B0(n198), .Y(n196) );
  NOR2X8 U600 ( .A(B[21]), .B(A[21]), .Y(n137) );
  XNOR2X2 U601 ( .A(n225), .B(n27), .Y(SUM[11]) );
  XOR2X4 U602 ( .A(n2), .B(n22), .Y(SUM[16]) );
  NAND2X6 U603 ( .A(B[25]), .B(A[25]), .Y(n100) );
  NOR2X6 U604 ( .A(B[24]), .B(A[24]), .Y(n106) );
  NOR2BX4 U605 ( .AN(n93), .B(n86), .Y(n84) );
  NOR2X8 U606 ( .A(n99), .B(n106), .Y(n93) );
  OAI21X4 U607 ( .A0(n99), .A1(n107), .B0(n100), .Y(n94) );
  NAND2X4 U608 ( .A(B[29]), .B(A[29]), .Y(n62) );
  NAND2X4 U609 ( .A(B[27]), .B(A[27]), .Y(n80) );
  NAND2X6 U610 ( .A(B[26]), .B(A[26]), .Y(n89) );
  INVX1 U611 ( .A(n99), .Y(n296) );
  XOR2X4 U612 ( .A(n475), .B(n25), .Y(SUM[13]) );
  NOR2X8 U613 ( .A(B[11]), .B(A[11]), .Y(n223) );
  NOR2X6 U614 ( .A(B[23]), .B(A[23]), .Y(n117) );
  NAND2X2 U615 ( .A(B[23]), .B(A[23]), .Y(n118) );
  OAI21X4 U616 ( .A0(n286), .A1(n289), .B0(n287), .Y(n285) );
  NAND2X2 U617 ( .A(n459), .B(n287), .Y(n37) );
  NOR2X8 U618 ( .A(B[18]), .B(A[18]), .Y(n162) );
  INVX6 U619 ( .A(n162), .Y(n303) );
  NOR2X8 U620 ( .A(B[9]), .B(A[9]), .Y(n241) );
  XNOR2X2 U621 ( .A(n196), .B(n24), .Y(SUM[14]) );
  AOI21X2 U622 ( .A0(n462), .A1(n317), .B0(n458), .Y(n473) );
  NAND2X6 U623 ( .A(n467), .B(n457), .Y(n232) );
  INVXL U624 ( .A(n235), .Y(n233) );
  XNOR2X4 U625 ( .A(n232), .B(n28), .Y(SUM[10]) );
  INVX3 U626 ( .A(n106), .Y(n297) );
  INVXL U627 ( .A(n107), .Y(n105) );
  XNOR2X4 U628 ( .A(n41), .B(n7), .Y(SUM[31]) );
  OAI21X2 U629 ( .A0(n61), .A1(n429), .B0(n62), .Y(n60) );
  NAND2X2 U630 ( .A(n217), .B(n309), .Y(n208) );
  NAND2XL U631 ( .A(n217), .B(n199), .Y(n197) );
  INVX1 U632 ( .A(n241), .Y(n312) );
  OAI21X4 U633 ( .A0(n241), .A1(n245), .B0(n242), .Y(n236) );
  OAI21X2 U634 ( .A0(n79), .A1(n89), .B0(n80), .Y(n78) );
  NAND2X2 U635 ( .A(n4), .B(n44), .Y(n42) );
  NOR2X8 U636 ( .A(n147), .B(n113), .Y(n4) );
  INVX3 U637 ( .A(n117), .Y(n298) );
  INVXL U638 ( .A(n244), .Y(n313) );
  INVXL U639 ( .A(n213), .Y(n211) );
  INVXL U640 ( .A(n167), .Y(n165) );
  NAND2XL U641 ( .A(n310), .B(n224), .Y(n27) );
  INVXL U642 ( .A(n223), .Y(n310) );
  NAND2XL U643 ( .A(n440), .B(n195), .Y(n24) );
  INVX3 U644 ( .A(n212), .Y(n309) );
  XOR2XL U645 ( .A(n246), .B(n30), .Y(SUM[8]) );
  INVXL U646 ( .A(n185), .Y(n306) );
  INVXL U647 ( .A(n61), .Y(n292) );
  OAI21X4 U648 ( .A0(n276), .A1(n248), .B0(n249), .Y(n247) );
  NAND2XL U649 ( .A(n309), .B(n213), .Y(n26) );
  OAI2BB1X4 U650 ( .A0N(n179), .A1N(n247), .B0(n478), .Y(n477) );
  CLKINVX1 U651 ( .A(n279), .Y(n318) );
  NOR2BX1 U652 ( .AN(n199), .B(n192), .Y(n190) );
  NAND2X1 U653 ( .A(n235), .B(n311), .Y(n226) );
  NAND2XL U654 ( .A(n167), .B(n303), .Y(n158) );
  NAND2X1 U655 ( .A(n122), .B(n149), .Y(n120) );
  NAND2X1 U656 ( .A(n319), .B(n283), .Y(n36) );
  NAND2XL U657 ( .A(n149), .B(n131), .Y(n129) );
  CLKINVX1 U658 ( .A(n176), .Y(n305) );
  XOR2X1 U659 ( .A(n37), .B(n289), .Y(SUM[1]) );
  NAND2X1 U660 ( .A(n313), .B(n245), .Y(n30) );
  CLKINVX1 U661 ( .A(n163), .Y(n161) );
  NAND2X1 U662 ( .A(n444), .B(n89), .Y(n12) );
  OA21X2 U663 ( .A0(n2), .A1(n120), .B0(n121), .Y(n479) );
  NAND2X1 U664 ( .A(n302), .B(n156), .Y(n19) );
  NAND2XL U665 ( .A(n299), .B(n127), .Y(n16) );
  NAND2XL U666 ( .A(n303), .B(n163), .Y(n20) );
  NAND2XL U667 ( .A(n311), .B(n231), .Y(n28) );
  OA21X4 U668 ( .A0(n148), .A1(n113), .B0(n114), .Y(n480) );
  INVXL U669 ( .A(n231), .Y(n229) );
  CLKINVX1 U670 ( .A(n145), .Y(n143) );
  NAND2XL U671 ( .A(n297), .B(n107), .Y(n14) );
  NAND2X2 U672 ( .A(n294), .B(n80), .Y(n11) );
  INVXL U673 ( .A(n79), .Y(n294) );
  NAND2X1 U674 ( .A(n315), .B(n260), .Y(n32) );
  CLKINVX1 U675 ( .A(n38), .Y(SUM[0]) );
  NAND2X1 U676 ( .A(n482), .B(n40), .Y(n7) );
  OR2XL U677 ( .A(B[31]), .B(A[31]), .Y(n482) );
  NAND2XL U678 ( .A(B[31]), .B(A[31]), .Y(n40) );
  NAND2XL U679 ( .A(n305), .B(n177), .Y(n22) );
  AOI21XL U680 ( .A0(n461), .A1(n303), .B0(n161), .Y(n159) );
endmodule


module ALU_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n11, n15, n17, n19, n20, n21, n23, n24, n25,
         n26, n28, n29, n30, n31, n33, n34, n36, n37, n39, n41, n42, n43, n44,
         n45, n46, n48, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n64, n65, n66, n67, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n88, n89, n91, n92, n93, n95, n98,
         n99, n100, n101, n102, n104, n105, n106, n109, n112, n113, n114, n115,
         n116, n117, n119, n120, n121, n122, n123, n126, n127, n128, n129,
         n130, n131, n133, n136, n137, n138, n139, n140, n142, n143, n144,
         n145, n147, n152, n153, n154, n155, n156, n157, n158, n160, n161,
         n162, n163, n164, n165, n166, n167, n172, n173, n174, n175, n176,
         n178, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n194, n195, n196, n197, n198, n199, n204, n205, n206,
         n207, n208, n210, n211, n212, n213, n214, n215, n216, n217, n220,
         n221, n222, n223, n225, n226, n228, n229, n230, n231, n232, n234,
         n235, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n259, n261, n262, n264,
         n267, n268, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n281, n282, n283, n284, n285, n286, n287, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n301, n303, n304, n305, n306,
         n307, n308, n309, n314, n315, n316, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523;

  OAI21X4 U288 ( .A0(n275), .A1(n247), .B0(n248), .Y(n246) );
  AOI21X4 U329 ( .A0(n276), .A1(n284), .B0(n277), .Y(n275) );
  CLKINVX12 U386 ( .A(B[4]), .Y(n522) );
  NAND2X8 U387 ( .A(n198), .B(n182), .Y(n180) );
  CLKAND2X12 U388 ( .A(B[16]), .B(n460), .Y(n175) );
  CLKINVX12 U389 ( .A(n475), .Y(n4) );
  XNOR2X1 U390 ( .A(n2), .B(n486), .Y(DIFF[16]) );
  INVX20 U391 ( .A(B[9]), .Y(n341) );
  CLKINVX12 U392 ( .A(n510), .Y(n517) );
  NOR2X6 U393 ( .A(n136), .B(n143), .Y(n130) );
  CLKAND2X12 U394 ( .A(A[16]), .B(n482), .Y(n499) );
  INVX3 U395 ( .A(n482), .Y(n172) );
  INVX4 U396 ( .A(n229), .Y(n309) );
  NOR2X8 U397 ( .A(n336), .B(A[14]), .Y(n191) );
  NAND2X8 U398 ( .A(n114), .B(n130), .Y(n112) );
  NAND2X6 U399 ( .A(n336), .B(A[14]), .Y(n194) );
  CLKINVX16 U400 ( .A(B[14]), .Y(n336) );
  CLKINVX16 U401 ( .A(n2), .Y(n456) );
  NOR2X8 U402 ( .A(n329), .B(A[21]), .Y(n136) );
  AND2X4 U403 ( .A(n4), .B(n65), .Y(n453) );
  NAND2X8 U404 ( .A(n456), .B(n453), .Y(n484) );
  NAND2X2 U405 ( .A(n309), .B(n230), .Y(n28) );
  CLKINVX4 U406 ( .A(n230), .Y(n228) );
  NAND2X4 U407 ( .A(n335), .B(A[15]), .Y(n185) );
  INVX20 U408 ( .A(B[7]), .Y(n343) );
  NOR2X8 U409 ( .A(n272), .B(n267), .Y(n261) );
  NOR2X8 U410 ( .A(n522), .B(A[4]), .Y(n272) );
  OAI21X2 U411 ( .A0(n473), .A1(n472), .B0(n194), .Y(n190) );
  NOR2X2 U412 ( .A(n336), .B(A[14]), .Y(n472) );
  INVX2 U413 ( .A(n262), .Y(n264) );
  INVX8 U414 ( .A(n458), .Y(n510) );
  NAND2BXL U415 ( .AN(n240), .B(n241), .Y(n29) );
  INVX6 U416 ( .A(n112), .Y(n476) );
  NOR2X8 U417 ( .A(n335), .B(A[15]), .Y(n184) );
  INVX4 U418 ( .A(B[3]), .Y(n521) );
  NAND2X4 U419 ( .A(n341), .B(A[9]), .Y(n241) );
  NOR2X8 U420 ( .A(n325), .B(A[25]), .Y(n98) );
  NAND2X4 U421 ( .A(n325), .B(A[25]), .Y(n99) );
  OAI21X2 U422 ( .A0(n95), .A1(n85), .B0(n88), .Y(n84) );
  INVXL U423 ( .A(n93), .Y(n95) );
  NOR2X4 U424 ( .A(n214), .B(n180), .Y(n178) );
  INVX20 U425 ( .A(B[1]), .Y(n518) );
  NAND2X8 U426 ( .A(n340), .B(A[10]), .Y(n230) );
  INVX2 U427 ( .A(n275), .Y(n274) );
  XNOR2X2 U428 ( .A(n503), .B(n33), .Y(DIFF[5]) );
  AO21X2 U429 ( .A0(n274), .A1(n315), .B0(n271), .Y(n503) );
  INVX12 U430 ( .A(B[5]), .Y(n523) );
  NOR2X8 U431 ( .A(n324), .B(A[26]), .Y(n85) );
  CLKINVX12 U432 ( .A(B[26]), .Y(n324) );
  AND2X8 U433 ( .A(n93), .B(n76), .Y(n494) );
  CLKINVX2 U434 ( .A(n222), .Y(n308) );
  AOI21X4 U435 ( .A0(n274), .A1(n254), .B0(n255), .Y(n253) );
  NAND2X4 U436 ( .A(n497), .B(n259), .Y(n255) );
  INVX16 U437 ( .A(B[22]), .Y(n328) );
  CLKINVX12 U438 ( .A(B[25]), .Y(n325) );
  CLKINVX2 U439 ( .A(n5), .Y(n75) );
  NAND2X4 U440 ( .A(n234), .B(n220), .Y(n214) );
  NOR2X6 U441 ( .A(n229), .B(n222), .Y(n220) );
  INVX20 U442 ( .A(n505), .Y(n2) );
  INVX20 U443 ( .A(B[10]), .Y(n340) );
  NAND2X4 U444 ( .A(n261), .B(n249), .Y(n247) );
  CLKINVX6 U445 ( .A(B[16]), .Y(n334) );
  INVX6 U446 ( .A(B[23]), .Y(n327) );
  INVX2 U447 ( .A(n204), .Y(n306) );
  CLKINVX8 U448 ( .A(B[28]), .Y(n322) );
  NAND2X6 U449 ( .A(n520), .B(A[2]), .Y(n282) );
  INVX12 U450 ( .A(B[6]), .Y(n344) );
  CLKINVX6 U451 ( .A(A[16]), .Y(n460) );
  AOI21X1 U452 ( .A0(n167), .A1(n301), .B0(n160), .Y(n158) );
  AOI21X1 U453 ( .A0(n463), .A1(n121), .B0(n122), .Y(n120) );
  NAND2X6 U454 ( .A(n326), .B(A[24]), .Y(n106) );
  AND2X2 U455 ( .A(n4), .B(n92), .Y(n465) );
  CLKXOR2X2 U456 ( .A(n245), .B(n30), .Y(DIFF[8]) );
  NAND2X2 U457 ( .A(n304), .B(n185), .Y(n23) );
  AND2X2 U458 ( .A(n4), .B(n54), .Y(n468) );
  NAND2X4 U459 ( .A(n490), .B(n491), .Y(DIFF[31]) );
  CLKINVX4 U460 ( .A(n504), .Y(n488) );
  OR2X6 U461 ( .A(n320), .B(A[30]), .Y(n511) );
  INVX3 U462 ( .A(n59), .Y(n57) );
  AND2X4 U463 ( .A(n291), .B(n70), .Y(n485) );
  NAND2X6 U464 ( .A(n520), .B(A[2]), .Y(n474) );
  XOR2X1 U465 ( .A(n37), .B(n287), .Y(DIFF[1]) );
  INVX1 U466 ( .A(n472), .Y(n305) );
  AND2X2 U467 ( .A(n303), .B(n176), .Y(n486) );
  CLKAND2X3 U468 ( .A(n299), .B(n144), .Y(n464) );
  XNOR2X2 U469 ( .A(n231), .B(n28), .Y(DIFF[10]) );
  INVX1 U470 ( .A(n234), .Y(n232) );
  NAND2X2 U471 ( .A(n307), .B(n212), .Y(n26) );
  NAND2X2 U472 ( .A(n481), .B(n155), .Y(n19) );
  INVX2 U473 ( .A(n116), .Y(n296) );
  CLKAND2X4 U474 ( .A(n290), .B(n61), .Y(n480) );
  CLKAND2X3 U475 ( .A(n294), .B(n99), .Y(n455) );
  CLKAND2X3 U476 ( .A(n293), .B(n88), .Y(n479) );
  AND2X8 U477 ( .A(n152), .B(n166), .Y(n454) );
  OAI2BB1X4 U478 ( .A0N(n456), .A1N(n454), .B0(n478), .Y(n145) );
  INVX3 U479 ( .A(n131), .Y(n133) );
  INVX16 U480 ( .A(B[11]), .Y(n339) );
  NOR2X8 U481 ( .A(n327), .B(A[23]), .Y(n116) );
  INVX3 U482 ( .A(n487), .Y(n283) );
  NAND2X2 U483 ( .A(n301), .B(n162), .Y(n20) );
  NAND2X6 U484 ( .A(n332), .B(A[18]), .Y(n162) );
  INVX3 U485 ( .A(n167), .Y(n165) );
  AO21X4 U486 ( .A0(n167), .A1(n152), .B0(n153), .Y(n463) );
  NOR2X6 U487 ( .A(n518), .B(A[1]), .Y(n285) );
  XOR2X4 U488 ( .A(n127), .B(n457), .Y(DIFF[22]) );
  CLKAND2X8 U489 ( .A(n297), .B(n126), .Y(n457) );
  NAND2X2 U490 ( .A(n329), .B(A[21]), .Y(n137) );
  XNOR2X1 U491 ( .A(n519), .B(A[0]), .Y(DIFF[0]) );
  OAI21X4 U492 ( .A0(n112), .A1(n147), .B0(n113), .Y(n458) );
  NOR2X8 U493 ( .A(n519), .B(A[0]), .Y(n287) );
  CLKINVX2 U494 ( .A(B[0]), .Y(n519) );
  NAND2X8 U495 ( .A(n522), .B(A[4]), .Y(n273) );
  OR2XL U496 ( .A(A[8]), .B(n342), .Y(n459) );
  INVX16 U497 ( .A(B[8]), .Y(n342) );
  NOR2X4 U498 ( .A(A[1]), .B(n518), .Y(n461) );
  CLKINVX12 U499 ( .A(B[12]), .Y(n338) );
  INVX3 U500 ( .A(n466), .Y(n462) );
  OA21X2 U501 ( .A0(n240), .A1(n244), .B0(n241), .Y(n466) );
  NAND2X4 U502 ( .A(n343), .B(A[7]), .Y(n252) );
  NOR2X6 U503 ( .A(n243), .B(n240), .Y(n234) );
  OAI2BB1X2 U504 ( .A0N(n274), .A1N(n261), .B0(n264), .Y(n514) );
  AOI21X2 U505 ( .A0(n463), .A1(n299), .B0(n142), .Y(n140) );
  NOR2X8 U506 ( .A(n154), .B(n161), .Y(n152) );
  XOR2X4 U507 ( .A(n145), .B(n464), .Y(DIFF[20]) );
  NAND2X6 U508 ( .A(n518), .B(A[1]), .Y(n286) );
  XNOR2X2 U509 ( .A(n512), .B(n513), .Y(DIFF[3]) );
  OAI2BB1X4 U510 ( .A0N(n456), .A1N(n465), .B0(n91), .Y(n89) );
  NAND2X6 U511 ( .A(n342), .B(A[8]), .Y(n244) );
  INVX8 U512 ( .A(n256), .Y(n469) );
  NOR2X8 U513 ( .A(n344), .B(A[6]), .Y(n256) );
  NOR2X8 U514 ( .A(n343), .B(A[7]), .Y(n251) );
  CLKINVX2 U515 ( .A(n133), .Y(n467) );
  OAI2BB1X4 U516 ( .A0N(n456), .A1N(n468), .B0(n53), .Y(n51) );
  CLKINVX1 U517 ( .A(n273), .Y(n271) );
  CLKINVX8 U518 ( .A(n469), .Y(n470) );
  CLKBUFX2 U519 ( .A(n130), .Y(n471) );
  NAND2X6 U520 ( .A(n344), .B(A[6]), .Y(n259) );
  OAI21X4 U521 ( .A0(n5), .A1(n67), .B0(n70), .Y(n66) );
  INVX4 U522 ( .A(n67), .Y(n291) );
  NOR2X8 U523 ( .A(n322), .B(A[28]), .Y(n67) );
  OA21X4 U524 ( .A0(n204), .A1(n212), .B0(n205), .Y(n473) );
  NAND2X6 U525 ( .A(n338), .B(A[12]), .Y(n212) );
  NAND2X8 U526 ( .A(n454), .B(n476), .Y(n475) );
  NOR2BX4 U527 ( .AN(n198), .B(n472), .Y(n189) );
  INVX3 U528 ( .A(B[30]), .Y(n320) );
  OR2XL U529 ( .A(n343), .B(A[7]), .Y(n477) );
  NAND2X6 U530 ( .A(n484), .B(n64), .Y(n62) );
  INVX3 U531 ( .A(n463), .Y(n478) );
  XOR2X4 U532 ( .A(n89), .B(n479), .Y(DIFF[26]) );
  XOR2X4 U533 ( .A(n62), .B(n480), .Y(DIFF[29]) );
  OAI21X4 U534 ( .A0(n184), .A1(n194), .B0(n185), .Y(n183) );
  NOR2X8 U535 ( .A(n321), .B(A[29]), .Y(n60) );
  CLKINVX8 U536 ( .A(B[29]), .Y(n321) );
  NAND2X2 U537 ( .A(n166), .B(n301), .Y(n157) );
  INVX3 U538 ( .A(n166), .Y(n164) );
  INVX3 U539 ( .A(n175), .Y(n303) );
  NAND2BXL U540 ( .AN(n461), .B(n286), .Y(n37) );
  NAND2X8 U541 ( .A(n334), .B(n499), .Y(n500) );
  OAI21X1 U542 ( .A0(n461), .A1(n287), .B0(n286), .Y(n487) );
  CLKINVX16 U543 ( .A(B[2]), .Y(n520) );
  CLKINVX2 U544 ( .A(n215), .Y(n217) );
  NOR2X8 U545 ( .A(n340), .B(A[10]), .Y(n229) );
  NOR2X4 U546 ( .A(A[8]), .B(n342), .Y(n243) );
  NAND2XL U547 ( .A(n459), .B(n244), .Y(n30) );
  NAND2X4 U548 ( .A(n337), .B(A[13]), .Y(n205) );
  NOR2X8 U549 ( .A(n337), .B(A[13]), .Y(n204) );
  CLKINVX12 U550 ( .A(B[13]), .Y(n337) );
  INVX3 U551 ( .A(n123), .Y(n297) );
  NOR2X8 U552 ( .A(n175), .B(n172), .Y(n166) );
  CLKINVX8 U553 ( .A(B[20]), .Y(n330) );
  NOR2X6 U554 ( .A(n330), .B(A[20]), .Y(n143) );
  NAND2X6 U555 ( .A(n488), .B(n7), .Y(n491) );
  NOR2X8 U556 ( .A(n184), .B(n191), .Y(n182) );
  AOI21X4 U557 ( .A0(n114), .A1(n131), .B0(n115), .Y(n113) );
  NOR2X8 U558 ( .A(n523), .B(A[5]), .Y(n267) );
  NAND2X8 U559 ( .A(n330), .B(A[20]), .Y(n144) );
  OR2X1 U560 ( .A(n331), .B(A[19]), .Y(n481) );
  CLKINVX12 U561 ( .A(B[19]), .Y(n331) );
  NAND2X8 U562 ( .A(B[17]), .B(n483), .Y(n482) );
  CLKINVX20 U563 ( .A(A[17]), .Y(n483) );
  INVX12 U564 ( .A(B[17]), .Y(n333) );
  INVX1 U565 ( .A(n136), .Y(n298) );
  NAND2X4 U566 ( .A(n504), .B(n489), .Y(n490) );
  NOR2X8 U567 ( .A(A[9]), .B(n341), .Y(n240) );
  AND2X8 U568 ( .A(n517), .B(n295), .Y(n498) );
  XOR2X4 U569 ( .A(n71), .B(n485), .Y(DIFF[28]) );
  NAND2X1 U570 ( .A(n477), .B(n252), .Y(n31) );
  NAND2X8 U571 ( .A(n500), .B(n173), .Y(n167) );
  CLKINVX2 U572 ( .A(n517), .Y(n109) );
  INVX4 U573 ( .A(n272), .Y(n315) );
  AND2X4 U574 ( .A(n59), .B(n511), .Y(n492) );
  NAND2X8 U575 ( .A(n322), .B(A[28]), .Y(n70) );
  NAND2X2 U576 ( .A(n4), .B(n83), .Y(n81) );
  NAND2X2 U577 ( .A(n4), .B(n43), .Y(n41) );
  OAI21X4 U578 ( .A0(n230), .A1(n222), .B0(n223), .Y(n221) );
  NAND2X4 U579 ( .A(n339), .B(A[11]), .Y(n223) );
  AOI21X2 U580 ( .A0(n217), .A1(n307), .B0(n210), .Y(n208) );
  INVX6 U581 ( .A(n211), .Y(n307) );
  NOR2X8 U582 ( .A(n494), .B(n77), .Y(n5) );
  OAI21X4 U583 ( .A0(n78), .A1(n88), .B0(n79), .Y(n77) );
  AOI21X4 U584 ( .A0(n262), .A1(n249), .B0(n250), .Y(n248) );
  NOR2X8 U585 ( .A(n251), .B(n256), .Y(n249) );
  NOR2X8 U586 ( .A(n78), .B(n85), .Y(n76) );
  NAND2X8 U587 ( .A(n92), .B(n76), .Y(n6) );
  NOR2X4 U588 ( .A(n6), .B(n56), .Y(n54) );
  NOR2X6 U589 ( .A(n498), .B(n104), .Y(n102) );
  AOI21X4 U590 ( .A0(n517), .A1(n83), .B0(n84), .Y(n82) );
  AOI21X2 U591 ( .A0(n463), .A1(n471), .B0(n467), .Y(n129) );
  INVX6 U592 ( .A(B[15]), .Y(n335) );
  OAI21X1 U593 ( .A0(n245), .A1(n214), .B0(n215), .Y(n213) );
  NOR2X8 U594 ( .A(n339), .B(A[11]), .Y(n222) );
  INVX1 U595 ( .A(n161), .Y(n301) );
  AOI21X4 U596 ( .A0(n517), .A1(n43), .B0(n44), .Y(n42) );
  NAND2X6 U597 ( .A(n324), .B(A[26]), .Y(n88) );
  AOI21X4 U598 ( .A0(n517), .A1(n65), .B0(n66), .Y(n64) );
  NOR2X8 U599 ( .A(n323), .B(A[27]), .Y(n78) );
  CLKINVX12 U600 ( .A(B[27]), .Y(n323) );
  OAI21X4 U601 ( .A0(n2), .A1(n81), .B0(n82), .Y(n80) );
  INVX1 U602 ( .A(n184), .Y(n304) );
  NAND2X4 U603 ( .A(n328), .B(A[22]), .Y(n126) );
  NAND2X4 U604 ( .A(n327), .B(A[23]), .Y(n117) );
  NAND2X4 U605 ( .A(n323), .B(A[27]), .Y(n79) );
  XOR2X4 U606 ( .A(n502), .B(n507), .Y(DIFF[11]) );
  OAI21X2 U607 ( .A0(n245), .A1(n225), .B0(n226), .Y(n502) );
  NOR2X8 U608 ( .A(n521), .B(A[3]), .Y(n278) );
  OAI21X4 U609 ( .A0(n5), .A1(n45), .B0(n46), .Y(n44) );
  OAI21X4 U610 ( .A0(n60), .A1(n70), .B0(n61), .Y(n59) );
  NAND2X4 U611 ( .A(n321), .B(A[29]), .Y(n61) );
  NAND2X4 U612 ( .A(n523), .B(A[5]), .Y(n268) );
  NOR2X8 U613 ( .A(n211), .B(n204), .Y(n198) );
  AOI21X4 U614 ( .A0(n199), .A1(n182), .B0(n183), .Y(n181) );
  AOI21X4 U615 ( .A0(n517), .A1(n74), .B0(n75), .Y(n73) );
  CLKINVX6 U616 ( .A(n6), .Y(n74) );
  OAI21X2 U617 ( .A0(n2), .A1(n175), .B0(n176), .Y(n174) );
  OAI21X4 U618 ( .A0(n2), .A1(n164), .B0(n165), .Y(n163) );
  AOI21X2 U619 ( .A0(n217), .A1(n198), .B0(n199), .Y(n197) );
  OR2X4 U620 ( .A(n319), .B(A[31]), .Y(n516) );
  CLKINVX6 U621 ( .A(B[31]), .Y(n319) );
  OAI21X4 U622 ( .A0(n2), .A1(n157), .B0(n158), .Y(n156) );
  OAI21X4 U623 ( .A0(n2), .A1(n128), .B0(n129), .Y(n127) );
  OAI21X2 U624 ( .A0(n2), .A1(n139), .B0(n140), .Y(n138) );
  INVX6 U625 ( .A(B[18]), .Y(n332) );
  OAI21X4 U626 ( .A0(n154), .A1(n162), .B0(n155), .Y(n153) );
  NOR2X8 U627 ( .A(n331), .B(A[19]), .Y(n154) );
  XNOR2X4 U628 ( .A(n508), .B(n509), .Y(DIFF[24]) );
  INVX4 U629 ( .A(n470), .Y(n496) );
  NOR2BX4 U630 ( .AN(n261), .B(n470), .Y(n254) );
  NAND2X4 U631 ( .A(n331), .B(A[19]), .Y(n155) );
  NOR2X6 U632 ( .A(n326), .B(A[24]), .Y(n105) );
  CLKINVX12 U633 ( .A(B[24]), .Y(n326) );
  INVX6 U634 ( .A(n214), .Y(n216) );
  INVX4 U635 ( .A(n246), .Y(n245) );
  XOR2X2 U636 ( .A(n514), .B(n515), .Y(DIFF[6]) );
  OAI21X2 U637 ( .A0(n245), .A1(n243), .B0(n244), .Y(n242) );
  XNOR2X4 U638 ( .A(n51), .B(n8), .Y(DIFF[30]) );
  XNOR2X2 U639 ( .A(n242), .B(n29), .Y(DIFF[9]) );
  AOI21X2 U640 ( .A0(n517), .A1(n92), .B0(n93), .Y(n91) );
  XNOR2X4 U641 ( .A(n174), .B(n21), .Y(DIFF[17]) );
  XOR2X4 U642 ( .A(n501), .B(n15), .Y(DIFF[23]) );
  OAI21X4 U643 ( .A0(n2), .A1(n72), .B0(n73), .Y(n71) );
  NOR2X6 U644 ( .A(n6), .B(n67), .Y(n65) );
  XOR2X4 U645 ( .A(n100), .B(n455), .Y(DIFF[25]) );
  NOR2X8 U646 ( .A(n98), .B(n105), .Y(n92) );
  INVX6 U647 ( .A(n105), .Y(n295) );
  NOR2BX4 U648 ( .AN(n92), .B(n85), .Y(n83) );
  OAI21X4 U649 ( .A0(n101), .A1(n2), .B0(n102), .Y(n100) );
  OAI21X4 U650 ( .A0(n116), .A1(n126), .B0(n117), .Y(n115) );
  OAI21X1 U651 ( .A0(n245), .A1(n232), .B0(n466), .Y(n231) );
  NOR2X8 U652 ( .A(n328), .B(A[22]), .Y(n123) );
  XNOR2X4 U653 ( .A(n163), .B(n20), .Y(DIFF[18]) );
  NOR2BX2 U654 ( .AN(n130), .B(n123), .Y(n121) );
  OAI21X1 U655 ( .A0(n133), .A1(n123), .B0(n126), .Y(n122) );
  NOR2X8 U656 ( .A(n116), .B(n123), .Y(n114) );
  AOI21X2 U657 ( .A0(n517), .A1(n54), .B0(n55), .Y(n53) );
  CLKINVX12 U658 ( .A(B[21]), .Y(n329) );
  OAI21X4 U659 ( .A0(n204), .A1(n212), .B0(n205), .Y(n199) );
  XNOR2X4 U660 ( .A(n156), .B(n19), .Y(DIFF[19]) );
  NAND2X4 U661 ( .A(n333), .B(A[17]), .Y(n173) );
  XOR2X4 U662 ( .A(n253), .B(n31), .Y(DIFF[7]) );
  NAND2X2 U663 ( .A(n121), .B(n454), .Y(n119) );
  XNOR2X4 U664 ( .A(n80), .B(n11), .Y(DIFF[27]) );
  OAI21X4 U665 ( .A0(n282), .A1(n278), .B0(n279), .Y(n277) );
  NAND2X4 U666 ( .A(n521), .B(A[3]), .Y(n279) );
  XNOR2X4 U667 ( .A(n206), .B(n25), .Y(DIFF[13]) );
  NOR2X8 U668 ( .A(n520), .B(A[2]), .Y(n281) );
  NAND2BX4 U669 ( .AN(n281), .B(n474), .Y(n36) );
  OA21X4 U670 ( .A0(n2), .A1(n119), .B0(n120), .Y(n501) );
  NOR2X4 U671 ( .A(n338), .B(A[12]), .Y(n211) );
  NOR2X4 U672 ( .A(n332), .B(A[18]), .Y(n161) );
  OAI21X4 U673 ( .A0(n267), .A1(n273), .B0(n268), .Y(n262) );
  OAI21X4 U674 ( .A0(n136), .A1(n144), .B0(n137), .Y(n131) );
  OAI21X4 U675 ( .A0(n240), .A1(n244), .B0(n241), .Y(n235) );
  OAI21X1 U676 ( .A0(n245), .A1(n196), .B0(n197), .Y(n195) );
  OA21X4 U677 ( .A0(n2), .A1(n41), .B0(n42), .Y(n504) );
  INVXL U678 ( .A(n7), .Y(n489) );
  NOR2X4 U679 ( .A(n492), .B(n48), .Y(n46) );
  OR2X4 U680 ( .A(n245), .B(n187), .Y(n493) );
  NAND2X4 U681 ( .A(n493), .B(n188), .Y(n186) );
  AOI21X2 U682 ( .A0(n217), .A1(n189), .B0(n190), .Y(n188) );
  XNOR2X4 U683 ( .A(n186), .B(n23), .Y(DIFF[15]) );
  OAI21X4 U684 ( .A0(n98), .A1(n106), .B0(n99), .Y(n93) );
  OAI21X2 U685 ( .A0(n5), .A1(n56), .B0(n57), .Y(n55) );
  NAND2X2 U686 ( .A(n495), .B(n496), .Y(n497) );
  INVX3 U687 ( .A(n264), .Y(n495) );
  AOI21X4 U688 ( .A0(n235), .A1(n220), .B0(n221), .Y(n215) );
  NOR2X4 U689 ( .A(n6), .B(n45), .Y(n43) );
  NAND2X4 U690 ( .A(n58), .B(n511), .Y(n45) );
  NAND2X1 U691 ( .A(n234), .B(n309), .Y(n225) );
  NAND2X2 U692 ( .A(n4), .B(n74), .Y(n72) );
  NAND2X1 U693 ( .A(n4), .B(n295), .Y(n101) );
  NOR2X6 U694 ( .A(n67), .B(n60), .Y(n58) );
  INVX4 U695 ( .A(n60), .Y(n290) );
  INVX4 U696 ( .A(n78), .Y(n292) );
  NAND2X1 U697 ( .A(n454), .B(n471), .Y(n128) );
  INVXL U698 ( .A(n106), .Y(n104) );
  AOI21X4 U699 ( .A0(n167), .A1(n152), .B0(n153), .Y(n147) );
  NAND2XL U700 ( .A(n334), .B(A[16]), .Y(n176) );
  OA21X4 U701 ( .A0(n2), .A1(n475), .B0(n109), .Y(n508) );
  AND2X1 U702 ( .A(n295), .B(n106), .Y(n509) );
  OAI21X4 U703 ( .A0(n285), .A1(n287), .B0(n286), .Y(n284) );
  NOR2X4 U704 ( .A(n281), .B(n278), .Y(n276) );
  OA21X4 U705 ( .A0(n215), .A1(n180), .B0(n181), .Y(n506) );
  NAND2X1 U706 ( .A(n189), .B(n216), .Y(n187) );
  NAND2X1 U707 ( .A(n216), .B(n198), .Y(n196) );
  INVX3 U708 ( .A(n58), .Y(n56) );
  INVXL U709 ( .A(n144), .Y(n142) );
  INVXL U710 ( .A(n162), .Y(n160) );
  NAND2XL U711 ( .A(n511), .B(n50), .Y(n8) );
  OAI21X4 U712 ( .A0(n251), .A1(n259), .B0(n252), .Y(n250) );
  INVXL U713 ( .A(n278), .Y(n316) );
  AND2XL U714 ( .A(n316), .B(n279), .Y(n513) );
  XOR2XL U715 ( .A(n283), .B(n36), .Y(DIFF[2]) );
  OAI2BB1X4 U716 ( .A0N(n246), .A1N(n178), .B0(n506), .Y(n505) );
  NAND2X1 U717 ( .A(n216), .B(n307), .Y(n207) );
  XNOR2X1 U718 ( .A(n213), .B(n26), .Y(DIFF[12]) );
  CLKINVX1 U719 ( .A(n50), .Y(n48) );
  XNOR2X1 U720 ( .A(n274), .B(n34), .Y(DIFF[4]) );
  NAND2X1 U721 ( .A(n315), .B(n273), .Y(n34) );
  AND2X2 U722 ( .A(n308), .B(n223), .Y(n507) );
  NAND2X1 U723 ( .A(n306), .B(n205), .Y(n25) );
  NAND2X1 U724 ( .A(n482), .B(n173), .Y(n21) );
  XNOR2X1 U725 ( .A(n195), .B(n24), .Y(DIFF[14]) );
  NAND2X1 U726 ( .A(n305), .B(n194), .Y(n24) );
  CLKINVX1 U727 ( .A(n143), .Y(n299) );
  NAND2X1 U728 ( .A(n296), .B(n117), .Y(n15) );
  CLKINVX1 U729 ( .A(n98), .Y(n294) );
  CLKINVX1 U730 ( .A(n85), .Y(n293) );
  NAND2X1 U731 ( .A(n292), .B(n79), .Y(n11) );
  NAND2XL U732 ( .A(n454), .B(n299), .Y(n139) );
  CLKINVX1 U733 ( .A(n212), .Y(n210) );
  NAND2X1 U734 ( .A(n314), .B(n268), .Y(n33) );
  CLKINVX1 U735 ( .A(n267), .Y(n314) );
  NAND2X1 U736 ( .A(n516), .B(n39), .Y(n7) );
  NAND2X1 U737 ( .A(n319), .B(A[31]), .Y(n39) );
  OA21XL U738 ( .A0(n283), .A1(n281), .B0(n474), .Y(n512) );
  AND2XL U739 ( .A(n469), .B(n259), .Y(n515) );
  NAND2X2 U740 ( .A(n320), .B(A[30]), .Y(n50) );
  XNOR2X2 U741 ( .A(n138), .B(n17), .Y(DIFF[21]) );
  NAND2XL U742 ( .A(n298), .B(n137), .Y(n17) );
  AOI21XL U743 ( .A0(n462), .A1(n309), .B0(n228), .Y(n226) );
  OAI21X2 U744 ( .A0(n245), .A1(n207), .B0(n208), .Y(n206) );
endmodule


module ALU_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n9, n10, n11, n12, n13, n14, n17, n18, n19, n20, n21,
         n22, n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n46, n47, n51, n52, n53, n54, n55, n56,
         n58, n59, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n118, n119, n122, n123, n124, n125, n126, n127, n128, n131, n134,
         n135, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216;

  NAND2X2 U171 ( .A(n98), .B(n64), .Y(n63) );
  CLKINVX4 U172 ( .A(n63), .Y(n209) );
  NOR2X1 U173 ( .A(n216), .B(B[1]), .Y(n131) );
  OR2XL U174 ( .A(n10), .B(B[30]), .Y(n207) );
  AND2X2 U175 ( .A(n40), .B(n32), .Y(n208) );
  NOR2X8 U176 ( .A(n55), .B(n213), .Y(n46) );
  NAND2X8 U177 ( .A(n211), .B(n209), .Y(n55) );
  NOR2X4 U178 ( .A(B[13]), .B(B[14]), .Y(n74) );
  AND2X2 U179 ( .A(n58), .B(n210), .Y(n211) );
  CLKINVX2 U180 ( .A(B[17]), .Y(n210) );
  NAND2X2 U181 ( .A(n209), .B(n210), .Y(n212) );
  NOR2X4 U182 ( .A(B[9]), .B(B[10]), .Y(n92) );
  NOR2X8 U183 ( .A(B[1]), .B(B[2]), .Y(n128) );
  NOR2X4 U184 ( .A(B[5]), .B(B[6]), .Y(n112) );
  NOR2X2 U185 ( .A(n29), .B(B[25]), .Y(n27) );
  NAND2X2 U186 ( .A(n46), .B(n208), .Y(n29) );
  BUFX8 U187 ( .A(n3), .Y(n215) );
  CLKBUFX3 U188 ( .A(n3), .Y(n216) );
  NOR2X1 U189 ( .A(n215), .B(n109), .Y(n108) );
  NAND2X1 U190 ( .A(n72), .B(n69), .Y(n68) );
  INVXL U191 ( .A(n40), .Y(n39) );
  INVXL U192 ( .A(n46), .Y(n47) );
  INVXL U193 ( .A(n21), .Y(n22) );
  NAND2XL U194 ( .A(n98), .B(n82), .Y(n79) );
  INVXL U195 ( .A(n83), .Y(n82) );
  INVXL U196 ( .A(n74), .Y(n73) );
  INVXL U197 ( .A(n92), .Y(n91) );
  INVXL U198 ( .A(n98), .Y(n99) );
  NAND2BXL U199 ( .AN(n4), .B(n215), .Y(n5) );
  NOR2XL U200 ( .A(n135), .B(n134), .Y(n4) );
  INVXL U201 ( .A(n55), .Y(n56) );
  NOR2XL U202 ( .A(n119), .B(n111), .Y(n110) );
  INVXL U203 ( .A(n119), .Y(n118) );
  INVXL U204 ( .A(n14), .Y(n13) );
  OR2XL U205 ( .A(B[19]), .B(B[20]), .Y(n213) );
  OR2XL U206 ( .A(B[28]), .B(B[27]), .Y(n214) );
  INVXL U207 ( .A(n27), .Y(n26) );
  INVX1 U208 ( .A(n110), .Y(n109) );
  CLKINVX1 U209 ( .A(n79), .Y(n80) );
  NAND2X2 U210 ( .A(n135), .B(n134), .Y(n3) );
  NOR2X1 U211 ( .A(n99), .B(n91), .Y(n90) );
  CLKINVX1 U212 ( .A(n112), .Y(n111) );
  NOR2X1 U213 ( .A(n47), .B(n39), .Y(n38) );
  NOR2X1 U214 ( .A(n79), .B(n73), .Y(n72) );
  CLKINVX1 U215 ( .A(A[1]), .Y(n135) );
  CLKINVX1 U216 ( .A(n5), .Y(DIFF[0]) );
  NOR2X2 U217 ( .A(n119), .B(n103), .Y(n98) );
  NAND2X1 U218 ( .A(n112), .B(n104), .Y(n103) );
  NOR2XL U219 ( .A(B[7]), .B(B[8]), .Y(n104) );
  XNOR2XL U220 ( .A(n36), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U221 ( .A(n215), .B(n37), .Y(n36) );
  INVX1 U222 ( .A(n38), .Y(n37) );
  XNOR2XL U223 ( .A(n54), .B(B[19]), .Y(DIFF[19]) );
  NOR2X1 U224 ( .A(n215), .B(n55), .Y(n54) );
  XNOR2XL U225 ( .A(n70), .B(B[15]), .Y(DIFF[15]) );
  NOR2X1 U226 ( .A(n216), .B(n71), .Y(n70) );
  CLKINVX1 U227 ( .A(n72), .Y(n71) );
  XNOR2XL U228 ( .A(n88), .B(B[11]), .Y(DIFF[11]) );
  NOR2X1 U229 ( .A(n216), .B(n89), .Y(n88) );
  CLKINVX1 U230 ( .A(n90), .Y(n89) );
  XNOR2XL U231 ( .A(n96), .B(B[9]), .Y(DIFF[9]) );
  NOR2X1 U232 ( .A(n216), .B(n99), .Y(n96) );
  XNOR2XL U233 ( .A(n116), .B(B[5]), .Y(DIFF[5]) );
  NOR2X1 U234 ( .A(n216), .B(n119), .Y(n116) );
  XNOR2XL U235 ( .A(n20), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U236 ( .A(n215), .B(n21), .Y(n20) );
  XNOR2XL U237 ( .A(n44), .B(B[21]), .Y(DIFF[21]) );
  NOR2X1 U238 ( .A(n215), .B(n47), .Y(n44) );
  XNOR2XL U239 ( .A(n78), .B(B[13]), .Y(DIFF[13]) );
  NOR2X1 U240 ( .A(n216), .B(n79), .Y(n78) );
  XNOR2XL U241 ( .A(n108), .B(B[7]), .Y(DIFF[7]) );
  XNOR2XL U242 ( .A(n126), .B(B[3]), .Y(DIFF[3]) );
  NOR2X1 U243 ( .A(n216), .B(n127), .Y(n126) );
  CLKINVX1 U244 ( .A(n128), .Y(n127) );
  XNOR2XL U245 ( .A(n12), .B(B[29]), .Y(DIFF[29]) );
  NOR2X1 U246 ( .A(n215), .B(n13), .Y(n12) );
  XNOR2XL U247 ( .A(n28), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U248 ( .A(n215), .B(n29), .Y(n28) );
  XNOR2XL U249 ( .A(n41), .B(B[22]), .Y(DIFF[22]) );
  NOR2X1 U250 ( .A(n215), .B(n42), .Y(n41) );
  NAND2X1 U251 ( .A(n46), .B(n43), .Y(n42) );
  INVXL U252 ( .A(B[21]), .Y(n43) );
  XNOR2XL U253 ( .A(n51), .B(B[20]), .Y(DIFF[20]) );
  NOR2X1 U254 ( .A(n215), .B(n52), .Y(n51) );
  NAND2X1 U255 ( .A(n56), .B(n53), .Y(n52) );
  INVXL U256 ( .A(B[19]), .Y(n53) );
  XNOR2XL U257 ( .A(n62), .B(B[17]), .Y(DIFF[17]) );
  NOR2X1 U258 ( .A(n215), .B(n63), .Y(n62) );
  XNOR2XL U259 ( .A(n67), .B(B[16]), .Y(DIFF[16]) );
  NOR2X1 U260 ( .A(n215), .B(n68), .Y(n67) );
  INVXL U261 ( .A(B[15]), .Y(n69) );
  XNOR2XL U262 ( .A(n75), .B(B[14]), .Y(DIFF[14]) );
  NOR2X1 U263 ( .A(n216), .B(n76), .Y(n75) );
  NAND2X1 U264 ( .A(n80), .B(n77), .Y(n76) );
  INVXL U265 ( .A(B[13]), .Y(n77) );
  XNOR2XL U266 ( .A(n85), .B(B[12]), .Y(DIFF[12]) );
  NOR2X1 U267 ( .A(n216), .B(n86), .Y(n85) );
  NAND2X1 U268 ( .A(n90), .B(n87), .Y(n86) );
  INVXL U269 ( .A(B[11]), .Y(n87) );
  XNOR2XL U270 ( .A(n93), .B(B[10]), .Y(DIFF[10]) );
  NOR2X1 U271 ( .A(n216), .B(n94), .Y(n93) );
  NAND2X1 U272 ( .A(n98), .B(n95), .Y(n94) );
  INVXL U273 ( .A(B[9]), .Y(n95) );
  XNOR2XL U274 ( .A(n105), .B(B[8]), .Y(DIFF[8]) );
  NOR2X1 U275 ( .A(n215), .B(n106), .Y(n105) );
  NAND2X1 U276 ( .A(n110), .B(n107), .Y(n106) );
  INVXL U277 ( .A(B[7]), .Y(n107) );
  XNOR2XL U278 ( .A(n113), .B(B[6]), .Y(DIFF[6]) );
  NOR2X1 U279 ( .A(n216), .B(n114), .Y(n113) );
  NAND2X1 U280 ( .A(n118), .B(n115), .Y(n114) );
  INVXL U281 ( .A(B[5]), .Y(n115) );
  XNOR2XL U282 ( .A(n123), .B(B[4]), .Y(DIFF[4]) );
  NOR2X1 U283 ( .A(n216), .B(n124), .Y(n123) );
  NAND2X1 U284 ( .A(n128), .B(n125), .Y(n124) );
  INVXL U285 ( .A(B[3]), .Y(n125) );
  XNOR2XL U286 ( .A(n33), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U287 ( .A(n215), .B(n34), .Y(n33) );
  NAND2X1 U288 ( .A(n38), .B(n35), .Y(n34) );
  INVXL U289 ( .A(B[23]), .Y(n35) );
  XNOR2XL U290 ( .A(n131), .B(B[2]), .Y(DIFF[2]) );
  XNOR2XL U291 ( .A(n59), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U292 ( .A(n215), .B(n212), .Y(n59) );
  XNOR2XL U293 ( .A(n25), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U294 ( .A(n215), .B(n26), .Y(n25) );
  XNOR2XL U295 ( .A(n6), .B(B[31]), .Y(DIFF[31]) );
  NOR2X1 U296 ( .A(n216), .B(n207), .Y(n6) );
  NAND2X2 U297 ( .A(n128), .B(n122), .Y(n119) );
  NOR2XL U298 ( .A(B[3]), .B(B[4]), .Y(n122) );
  NOR2XL U299 ( .A(B[21]), .B(B[22]), .Y(n40) );
  INVXL U300 ( .A(B[18]), .Y(n58) );
  NAND2X1 U301 ( .A(n27), .B(n24), .Y(n21) );
  INVXL U302 ( .A(B[26]), .Y(n24) );
  INVX1 U303 ( .A(B[0]), .Y(n134) );
  NOR2X1 U304 ( .A(n21), .B(n214), .Y(n14) );
  NAND2X1 U305 ( .A(n14), .B(n11), .Y(n10) );
  INVXL U306 ( .A(B[29]), .Y(n11) );
  NOR2XL U307 ( .A(B[23]), .B(B[24]), .Y(n32) );
  NOR2X1 U308 ( .A(n83), .B(n65), .Y(n64) );
  NAND2X1 U309 ( .A(n74), .B(n66), .Y(n65) );
  NOR2XL U310 ( .A(B[15]), .B(B[16]), .Y(n66) );
  NAND2X1 U311 ( .A(n92), .B(n84), .Y(n83) );
  NOR2XL U312 ( .A(B[11]), .B(B[12]), .Y(n84) );
  XNOR2XL U313 ( .A(n9), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U314 ( .A(n215), .B(n10), .Y(n9) );
  XNOR2XL U315 ( .A(n17), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U316 ( .A(n215), .B(n18), .Y(n17) );
  NAND2X1 U317 ( .A(n22), .B(n19), .Y(n18) );
  INVXL U318 ( .A(B[27]), .Y(n19) );
  XOR2XL U319 ( .A(n215), .B(B[1]), .Y(DIFF[1]) );
endmodule


module ALU_DW01_inc_2 ( A, SUM );
  input [32:0] A;
  output [32:0] SUM;
  wire   n1, n2, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15, n16, n17, n18,
         n19, n21, n23, n24, n25, n26, n27, n28, n29, n30, n32, n34, n35, n36,
         n37, n38, n39, n40, n41, n43, n44, n45, n46, n48, n49, n50, n51, n52,
         n54, n55, n56, n57, n58, n59, n63, n64, n65, n66, n69, n70, n74, n75,
         n76, n77, n78, n79, n80, n81, n83, n84, n85, n87, n88, n89, n90, n91,
         n92, n94, n95, n96, n97, n98, n99, n101, n103, n104, n105, n106, n109,
         n110, n111, n112, n114, n115, n116, n117, n118, n119, n121, n122,
         n123, n124, n125, n126, n127, n128, n130, n131, n133, n134, n135,
         n137, n139, n140, n141, n142, n143, n144, n146, n147, n149, n150,
         n151, n153, n225, n226, n227;
  assign n8 = A[31];
  assign n12 = A[30];
  assign n19 = A[29];
  assign n23 = A[28];
  assign n30 = A[27];
  assign n34 = A[26];
  assign n39 = A[25];
  assign n43 = A[24];
  assign n50 = A[23];
  assign n54 = A[22];
  assign n59 = A[21];
  assign n63 = A[20];
  assign n70 = A[19];
  assign n74 = A[18];
  assign n79 = A[17];
  assign n83 = A[16];
  assign n90 = A[15];
  assign n94 = A[14];
  assign n99 = A[13];
  assign n103 = A[12];
  assign n110 = A[11];
  assign n114 = A[10];
  assign n119 = A[9];
  assign n122 = A[8];
  assign n128 = A[7];
  assign n131 = A[6];
  assign n135 = A[5];
  assign n139 = A[4];
  assign n144 = A[3];
  assign n147 = A[2];
  assign n151 = A[1];
  assign n153 = A[0];

  INVXL U190 ( .A(n78), .Y(n77) );
  INVXL U191 ( .A(n227), .Y(n85) );
  INVX1 U192 ( .A(n125), .Y(n124) );
  NOR2XL U193 ( .A(n141), .B(n134), .Y(n133) );
  NOR2BXL U194 ( .AN(n106), .B(n98), .Y(n97) );
  INVXL U195 ( .A(n118), .Y(n117) );
  NAND2XL U196 ( .A(n124), .B(n106), .Y(n105) );
  NAND2XL U197 ( .A(n37), .B(n227), .Y(n36) );
  NOR2XL U198 ( .A(n2), .B(n38), .Y(n37) );
  NAND2XL U199 ( .A(n15), .B(n227), .Y(n14) );
  NOR2XL U200 ( .A(n2), .B(n16), .Y(n15) );
  NAND2XL U201 ( .A(n28), .B(n17), .Y(n16) );
  INVXL U202 ( .A(n18), .Y(n17) );
  NAND2XL U203 ( .A(n26), .B(n227), .Y(n25) );
  NOR2XL U204 ( .A(n2), .B(n27), .Y(n26) );
  INVXL U205 ( .A(n28), .Y(n27) );
  NAND2XL U206 ( .A(n227), .B(n46), .Y(n45) );
  INVXL U207 ( .A(n2), .Y(n46) );
  NOR2BXL U208 ( .AN(n66), .B(n58), .Y(n57) );
  NAND2XL U209 ( .A(n227), .B(n66), .Y(n65) );
  NAND2XL U210 ( .A(n227), .B(n77), .Y(n76) );
  INVXL U211 ( .A(n142), .Y(n141) );
  XOR2XL U212 ( .A(n36), .B(n35), .Y(SUM[26]) );
  XOR2XL U213 ( .A(n65), .B(n64), .Y(SUM[20]) );
  INVXL U214 ( .A(n150), .Y(n149) );
  XOR2XL U215 ( .A(n25), .B(n24), .Y(SUM[28]) );
  XOR2XL U216 ( .A(n32), .B(n30), .Y(SUM[27]) );
  XOR2XL U217 ( .A(n137), .B(n135), .Y(SUM[5]) );
  XOR2XL U218 ( .A(n149), .B(n147), .Y(SUM[2]) );
  XNOR2XL U219 ( .A(n146), .B(n144), .Y(SUM[3]) );
  XOR2XL U220 ( .A(n21), .B(n19), .Y(SUM[29]) );
  XNOR2XL U221 ( .A(n124), .B(n123), .Y(SUM[8]) );
  INVXL U222 ( .A(n122), .Y(n123) );
  XOR2XL U223 ( .A(n101), .B(n99), .Y(SUM[13]) );
  XNOR2XL U224 ( .A(n130), .B(n128), .Y(SUM[7]) );
  INVXL U225 ( .A(n79), .Y(n80) );
  INVXL U226 ( .A(n50), .Y(n51) );
  INVXL U227 ( .A(n90), .Y(n91) );
  INVXL U228 ( .A(n110), .Y(n111) );
  XNOR2XL U229 ( .A(n121), .B(n119), .Y(SUM[9]) );
  XOR2XL U230 ( .A(n133), .B(n131), .Y(SUM[6]) );
  INVXL U231 ( .A(n39), .Y(n40) );
  XOR2XL U232 ( .A(n10), .B(n8), .Y(SUM[31]) );
  XOR2XL U233 ( .A(n151), .B(n153), .Y(SUM[1]) );
  NOR2X1 U234 ( .A(n78), .B(n69), .Y(n66) );
  INVXL U235 ( .A(n12), .Y(n13) );
  INVXL U236 ( .A(n23), .Y(n24) );
  INVXL U237 ( .A(n34), .Y(n35) );
  INVXL U238 ( .A(n43), .Y(n44) );
  INVXL U239 ( .A(n54), .Y(n55) );
  INVXL U240 ( .A(n83), .Y(n84) );
  INVXL U241 ( .A(n94), .Y(n95) );
  INVXL U242 ( .A(n103), .Y(n104) );
  INVXL U243 ( .A(n114), .Y(n115) );
  INVXL U244 ( .A(n139), .Y(n140) );
  INVXL U245 ( .A(n63), .Y(n64) );
  INVXL U246 ( .A(n74), .Y(n75) );
  XOR2X1 U247 ( .A(n45), .B(n44), .Y(SUM[24]) );
  XOR2X1 U248 ( .A(n56), .B(n55), .Y(SUM[22]) );
  XOR2X1 U249 ( .A(n76), .B(n75), .Y(SUM[18]) );
  XOR2X1 U250 ( .A(n105), .B(n104), .Y(SUM[12]) );
  XOR2X1 U251 ( .A(n141), .B(n140), .Y(SUM[4]) );
  XOR2X1 U252 ( .A(n14), .B(n13), .Y(SUM[30]) );
  XOR2X1 U253 ( .A(n85), .B(n84), .Y(SUM[16]) );
  XOR2X1 U254 ( .A(n116), .B(n115), .Y(SUM[10]) );
  NAND2X1 U255 ( .A(n97), .B(n124), .Y(n96) );
  NAND2X1 U256 ( .A(n124), .B(n117), .Y(n116) );
  NAND2X1 U257 ( .A(n4), .B(n227), .Y(SUM[32]) );
  NAND2X1 U258 ( .A(n227), .B(n57), .Y(n56) );
  BUFX4 U259 ( .A(n1), .Y(n227) );
  NOR2X1 U260 ( .A(n87), .B(n125), .Y(n1) );
  NAND2X1 U261 ( .A(n106), .B(n88), .Y(n87) );
  NOR2X1 U262 ( .A(n98), .B(n89), .Y(n88) );
  XOR2X1 U263 ( .A(n96), .B(n95), .Y(SUM[14]) );
  NAND2X1 U264 ( .A(n149), .B(n147), .Y(n146) );
  NOR2X1 U265 ( .A(n36), .B(n35), .Y(n32) );
  XNOR2X1 U266 ( .A(n52), .B(n51), .Y(SUM[23]) );
  NOR2X1 U267 ( .A(n56), .B(n55), .Y(n52) );
  NOR2X1 U268 ( .A(n105), .B(n104), .Y(n101) );
  NAND2X1 U269 ( .A(n133), .B(n131), .Y(n130) );
  XNOR2X1 U270 ( .A(n41), .B(n40), .Y(SUM[25]) );
  NOR2X1 U271 ( .A(n45), .B(n44), .Y(n41) );
  NOR2X1 U272 ( .A(n25), .B(n24), .Y(n21) );
  XNOR2X1 U273 ( .A(n81), .B(n80), .Y(SUM[17]) );
  NOR2X1 U274 ( .A(n85), .B(n84), .Y(n81) );
  XNOR2X1 U275 ( .A(n92), .B(n91), .Y(SUM[15]) );
  NOR2X1 U276 ( .A(n96), .B(n95), .Y(n92) );
  XNOR2X1 U277 ( .A(n112), .B(n111), .Y(SUM[11]) );
  NOR2X1 U278 ( .A(n116), .B(n115), .Y(n112) );
  NAND2X1 U279 ( .A(n124), .B(n122), .Y(n121) );
  NOR2X1 U280 ( .A(n141), .B(n140), .Y(n137) );
  CLKINVX1 U281 ( .A(n153), .Y(SUM[0]) );
  NOR2X1 U282 ( .A(n14), .B(n13), .Y(n10) );
  NAND2X2 U283 ( .A(n66), .B(n48), .Y(n2) );
  NOR2X1 U284 ( .A(n58), .B(n49), .Y(n48) );
  NAND2X1 U285 ( .A(n54), .B(n50), .Y(n49) );
  NOR2X1 U286 ( .A(n38), .B(n29), .Y(n28) );
  NAND2X1 U287 ( .A(n34), .B(n30), .Y(n29) );
  NOR2X2 U288 ( .A(n118), .B(n109), .Y(n106) );
  NAND2X1 U289 ( .A(n114), .B(n110), .Y(n109) );
  NAND2X1 U290 ( .A(n74), .B(n70), .Y(n69) );
  XNOR2X1 U291 ( .A(n225), .B(n59), .Y(SUM[21]) );
  OR2X1 U292 ( .A(n65), .B(n64), .Y(n225) );
  XNOR2X1 U293 ( .A(n226), .B(n70), .Y(SUM[19]) );
  OR2X1 U294 ( .A(n76), .B(n75), .Y(n226) );
  NOR2X1 U295 ( .A(n143), .B(n150), .Y(n142) );
  NAND2X1 U296 ( .A(n147), .B(n144), .Y(n143) );
  NAND2X1 U297 ( .A(n103), .B(n99), .Y(n98) );
  NAND2X1 U298 ( .A(n139), .B(n135), .Y(n134) );
  NAND2X1 U299 ( .A(n43), .B(n39), .Y(n38) );
  NAND2X1 U300 ( .A(n63), .B(n59), .Y(n58) );
  NAND2X1 U301 ( .A(n122), .B(n119), .Y(n118) );
  NAND2X1 U302 ( .A(n23), .B(n19), .Y(n18) );
  NAND2X1 U303 ( .A(n83), .B(n79), .Y(n78) );
  NAND2X1 U304 ( .A(n153), .B(n151), .Y(n150) );
  NOR2X1 U305 ( .A(n2), .B(n5), .Y(n4) );
  NAND2X1 U306 ( .A(n28), .B(n6), .Y(n5) );
  NOR2X1 U307 ( .A(n18), .B(n7), .Y(n6) );
  NAND2X1 U308 ( .A(n12), .B(n8), .Y(n7) );
  NAND2X1 U309 ( .A(n126), .B(n142), .Y(n125) );
  NOR2X1 U310 ( .A(n134), .B(n127), .Y(n126) );
  NAND2X1 U311 ( .A(n131), .B(n128), .Y(n127) );
  NAND2X1 U312 ( .A(n94), .B(n90), .Y(n89) );
endmodule


module ALU_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32,
         n33, n34, n36, n37, n38, n39, n40, n41, n42, n46, n47, n48, n49, n50,
         n51, n53, n54, n55, n56, n57, n58, n62, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85,
         n86, n87, n88, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n102, n103, n104, n105, n106, n107, n108, n109, n211, n212, n213,
         n214, n215, n216, n218;

  OR2XL U144 ( .A(B[16]), .B(B[17]), .Y(n211) );
  AND2X6 U145 ( .A(n64), .B(n93), .Y(n216) );
  INVX16 U146 ( .A(n216), .Y(n218) );
  XOR2XL U147 ( .A(B[1]), .B(B[0]), .Y(DIFF[1]) );
  XNOR2XL U148 ( .A(n91), .B(B[9]), .Y(DIFF[9]) );
  OR2X8 U149 ( .A(B[20]), .B(B[21]), .Y(n212) );
  BUFX3 U150 ( .A(n99), .Y(n213) );
  NAND2X1 U151 ( .A(n95), .B(n213), .Y(n94) );
  INVX1 U152 ( .A(n213), .Y(n100) );
  XNOR2XL U153 ( .A(n78), .B(B[12]), .Y(DIFF[12]) );
  NOR2XL U154 ( .A(B[1]), .B(B[0]), .Y(n109) );
  CLKINVX4 U155 ( .A(n212), .Y(n214) );
  CLKINVX4 U156 ( .A(n211), .Y(n215) );
  NOR2XL U157 ( .A(n212), .B(B[22]), .Y(n40) );
  XNOR2XL U158 ( .A(n41), .B(B[22]), .Y(DIFF[22]) );
  NOR2XL U159 ( .A(B[22]), .B(B[23]), .Y(n37) );
  NOR2XL U160 ( .A(B[6]), .B(B[7]), .Y(n95) );
  XNOR2XL U161 ( .A(n70), .B(B[14]), .Y(DIFF[14]) );
  NOR2XL U162 ( .A(B[14]), .B(B[15]), .Y(n66) );
  NOR2XL U163 ( .A(B[26]), .B(B[27]), .Y(n21) );
  NOR2XL U164 ( .A(B[12]), .B(B[13]), .Y(n72) );
  XNOR2XL U165 ( .A(n49), .B(B[20]), .Y(DIFF[20]) );
  XNOR2XL U166 ( .A(n75), .B(B[13]), .Y(DIFF[13]) );
  INVX1 U167 ( .A(n72), .Y(n73) );
  NAND2X1 U168 ( .A(n66), .B(n72), .Y(n65) );
  NOR2XL U169 ( .A(B[5]), .B(B[4]), .Y(n99) );
  INVXL U170 ( .A(B[12]), .Y(n77) );
  INVX4 U171 ( .A(n93), .Y(n92) );
  INVXL U172 ( .A(n109), .Y(n108) );
  NOR2XL U173 ( .A(n92), .B(B[8]), .Y(n91) );
  NAND2XL U174 ( .A(n51), .B(n214), .Y(n42) );
  NOR2XL U175 ( .A(n68), .B(n92), .Y(n67) );
  NOR2XL U176 ( .A(n73), .B(B[14]), .Y(n69) );
  INVXL U177 ( .A(B[20]), .Y(n48) );
  NOR2X1 U178 ( .A(n16), .B(n218), .Y(n15) );
  NOR2XL U179 ( .A(n92), .B(n87), .Y(n86) );
  NOR2XL U180 ( .A(n76), .B(n92), .Y(n75) );
  NOR2XL U181 ( .A(n71), .B(n92), .Y(n70) );
  INVXL U182 ( .A(n27), .Y(n28) );
  NAND2X2 U183 ( .A(n215), .B(n53), .Y(n50) );
  NOR2X1 U184 ( .A(n23), .B(n218), .Y(n22) );
  NOR2XL U185 ( .A(n28), .B(B[26]), .Y(n24) );
  NOR2X1 U186 ( .A(n31), .B(n218), .Y(n30) );
  INVXL U187 ( .A(B[24]), .Y(n32) );
  INVXL U188 ( .A(n215), .Y(n58) );
  XNOR2XL U189 ( .A(n46), .B(B[21]), .Y(DIFF[21]) );
  NAND2X2 U190 ( .A(n88), .B(n82), .Y(n79) );
  XNOR2XL U191 ( .A(n25), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U192 ( .A(n11), .B(n218), .Y(n10) );
  XNOR2XL U193 ( .A(n18), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U194 ( .A(n19), .B(n218), .Y(n18) );
  XNOR2XL U195 ( .A(n33), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U196 ( .A(n218), .B(n34), .Y(n33) );
  INVXL U197 ( .A(n3), .Y(n34) );
  NOR2XL U198 ( .A(n218), .B(n42), .Y(n41) );
  NAND2XL U199 ( .A(n3), .B(n17), .Y(n16) );
  NOR2XL U200 ( .A(n4), .B(B[28]), .Y(n17) );
  XOR2XL U201 ( .A(n102), .B(B[5]), .Y(DIFF[5]) );
  NAND2X1 U202 ( .A(n104), .B(n103), .Y(n102) );
  INVXL U203 ( .A(B[4]), .Y(n103) );
  XNOR2XL U204 ( .A(n104), .B(B[4]), .Y(DIFF[4]) );
  NOR2XL U205 ( .A(B[28]), .B(B[29]), .Y(n14) );
  NAND2X2 U206 ( .A(n106), .B(n109), .Y(n105) );
  XOR2XL U207 ( .A(n96), .B(B[7]), .Y(DIFF[7]) );
  NAND2X1 U208 ( .A(n97), .B(n104), .Y(n96) );
  NOR2XL U209 ( .A(n100), .B(B[6]), .Y(n97) );
  XOR2XL U210 ( .A(n98), .B(B[6]), .Y(DIFF[6]) );
  NOR2XL U211 ( .A(n4), .B(n8), .Y(n7) );
  NAND2XL U212 ( .A(n14), .B(n9), .Y(n8) );
  NAND2XL U213 ( .A(n80), .B(n72), .Y(n71) );
  NOR2X1 U214 ( .A(n79), .B(n65), .Y(n64) );
  CLKINVX1 U215 ( .A(n105), .Y(n104) );
  CLKINVX1 U216 ( .A(n79), .Y(n80) );
  CLKINVX1 U217 ( .A(n50), .Y(n51) );
  CLKINVX1 U218 ( .A(n14), .Y(n13) );
  NOR2X2 U219 ( .A(n50), .B(n36), .Y(n3) );
  NAND2X1 U220 ( .A(n214), .B(n37), .Y(n36) );
  XNOR2X1 U221 ( .A(n57), .B(B[18]), .Y(DIFF[18]) );
  NOR2XL U222 ( .A(n218), .B(n58), .Y(n57) );
  NOR2X1 U223 ( .A(B[8]), .B(B[9]), .Y(n88) );
  NOR2X1 U224 ( .A(B[24]), .B(B[25]), .Y(n27) );
  NAND2X1 U225 ( .A(n27), .B(n21), .Y(n4) );
  NOR2X1 U226 ( .A(B[10]), .B(B[11]), .Y(n82) );
  NOR2X1 U227 ( .A(B[18]), .B(B[19]), .Y(n53) );
  NOR2X2 U228 ( .A(n94), .B(n105), .Y(n93) );
  NOR2XL U229 ( .A(n92), .B(n79), .Y(n78) );
  XNOR2X1 U230 ( .A(n83), .B(B[11]), .Y(DIFF[11]) );
  NOR2XL U231 ( .A(n92), .B(n84), .Y(n83) );
  NAND2XL U232 ( .A(n88), .B(n85), .Y(n84) );
  CLKINVX1 U233 ( .A(B[10]), .Y(n85) );
  XNOR2X1 U234 ( .A(n86), .B(B[10]), .Y(DIFF[10]) );
  INVXL U235 ( .A(n88), .Y(n87) );
  XNOR2X1 U236 ( .A(n67), .B(B[15]), .Y(DIFF[15]) );
  NAND2XL U237 ( .A(n69), .B(n80), .Y(n68) );
  NAND2XL U238 ( .A(n80), .B(n77), .Y(n76) );
  NOR2X1 U239 ( .A(B[3]), .B(B[2]), .Y(n106) );
  CLKINVX1 U240 ( .A(B[30]), .Y(n9) );
  XNOR2X1 U241 ( .A(n5), .B(B[31]), .Y(DIFF[31]) );
  NOR2X1 U242 ( .A(n6), .B(n218), .Y(n5) );
  NAND2XL U243 ( .A(n3), .B(n7), .Y(n6) );
  XNOR2X1 U244 ( .A(n15), .B(B[29]), .Y(DIFF[29]) );
  XNOR2X1 U245 ( .A(n10), .B(B[30]), .Y(DIFF[30]) );
  NAND2XL U246 ( .A(n3), .B(n12), .Y(n11) );
  NOR2XL U247 ( .A(n4), .B(n13), .Y(n12) );
  NOR2XL U248 ( .A(n26), .B(n218), .Y(n25) );
  NAND2XL U249 ( .A(n3), .B(n27), .Y(n26) );
  XNOR2X1 U250 ( .A(n30), .B(B[25]), .Y(DIFF[25]) );
  NAND2XL U251 ( .A(n3), .B(n32), .Y(n31) );
  NAND2XL U252 ( .A(n3), .B(n20), .Y(n19) );
  INVXL U253 ( .A(n4), .Y(n20) );
  XNOR2X1 U254 ( .A(n22), .B(B[27]), .Y(DIFF[27]) );
  NAND2XL U255 ( .A(n3), .B(n24), .Y(n23) );
  XOR2XL U256 ( .A(n92), .B(B[8]), .Y(DIFF[8]) );
  XNOR2X1 U257 ( .A(n62), .B(B[17]), .Y(DIFF[17]) );
  NOR2XL U258 ( .A(n218), .B(B[16]), .Y(n62) );
  NOR2XL U259 ( .A(n218), .B(n50), .Y(n49) );
  NOR2XL U260 ( .A(n218), .B(n47), .Y(n46) );
  NAND2XL U261 ( .A(n51), .B(n48), .Y(n47) );
  XNOR2X1 U262 ( .A(n54), .B(B[19]), .Y(DIFF[19]) );
  NOR2XL U263 ( .A(n218), .B(n55), .Y(n54) );
  NAND2XL U264 ( .A(n215), .B(n56), .Y(n55) );
  CLKINVX1 U265 ( .A(B[18]), .Y(n56) );
  XNOR2X1 U266 ( .A(n38), .B(B[23]), .Y(DIFF[23]) );
  NOR2XL U267 ( .A(n218), .B(n39), .Y(n38) );
  NAND2XL U268 ( .A(n40), .B(n51), .Y(n39) );
  XNOR2X1 U269 ( .A(n107), .B(B[3]), .Y(DIFF[3]) );
  NOR2X1 U270 ( .A(n108), .B(B[2]), .Y(n107) );
  XOR2XL U271 ( .A(n108), .B(B[2]), .Y(DIFF[2]) );
  NAND2XL U272 ( .A(n104), .B(n213), .Y(n98) );
  XOR2XL U273 ( .A(n218), .B(B[16]), .Y(DIFF[16]) );
  CLKBUFX2 U274 ( .A(B[0]), .Y(DIFF[0]) );
endmodule


module ALU_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30, n31, n32, n33,
         n34, n36, n37, n38, n39, n40, n41, n42, n43, n46, n47, n48, n49, n50,
         n51, n53, n54, n55, n56, n57, n58, n59, n62, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85,
         n86, n87, n88, n91, n92, n93, n94, n95, n96, n97, n98, n99, n102,
         n104, n105, n106, n107, n108, n109, n211, n212, n213, n214, n215;

  XNOR2X1 U144 ( .A(n78), .B(B[12]), .Y(DIFF[12]) );
  CLKINVX2 U145 ( .A(B[12]), .Y(n77) );
  NOR2X4 U146 ( .A(B[12]), .B(B[13]), .Y(n72) );
  AND2X8 U147 ( .A(n93), .B(n64), .Y(n211) );
  INVX16 U148 ( .A(n211), .Y(n212) );
  NAND2X1 U149 ( .A(n88), .B(n82), .Y(n79) );
  CLKINVX4 U150 ( .A(n79), .Y(n80) );
  NOR2X1 U151 ( .A(n92), .B(n79), .Y(n78) );
  NOR2X6 U152 ( .A(n214), .B(B[5]), .Y(n99) );
  INVX3 U153 ( .A(n215), .Y(n214) );
  NOR2XL U154 ( .A(B[21]), .B(B[20]), .Y(n43) );
  INVX1 U155 ( .A(B[20]), .Y(n48) );
  INVXL U156 ( .A(B[4]), .Y(n215) );
  NOR2XL U157 ( .A(B[7]), .B(B[6]), .Y(n95) );
  NOR2BXL U158 ( .AN(n99), .B(B[6]), .Y(n97) );
  XOR2X1 U159 ( .A(n98), .B(B[6]), .Y(DIFF[6]) );
  CLKBUFX2 U160 ( .A(B[2]), .Y(n213) );
  XNOR2X2 U161 ( .A(n70), .B(B[14]), .Y(DIFF[14]) );
  NOR2BX1 U162 ( .AN(n72), .B(B[14]), .Y(n69) );
  XOR2X1 U163 ( .A(n92), .B(B[8]), .Y(DIFF[8]) );
  NOR2X2 U164 ( .A(n92), .B(B[8]), .Y(n91) );
  XNOR2X1 U165 ( .A(n38), .B(B[23]), .Y(DIFF[23]) );
  NAND2XL U166 ( .A(n104), .B(n215), .Y(n102) );
  NAND2XL U167 ( .A(n3), .B(n20), .Y(n19) );
  INVXL U168 ( .A(n50), .Y(n51) );
  NOR2XL U169 ( .A(n212), .B(n50), .Y(n49) );
  INVX1 U170 ( .A(n105), .Y(n104) );
  NOR2XL U171 ( .A(n108), .B(n213), .Y(n107) );
  NAND2XL U172 ( .A(n104), .B(n99), .Y(n98) );
  NAND2XL U173 ( .A(n3), .B(n27), .Y(n26) );
  INVXL U174 ( .A(n4), .Y(n20) );
  NOR2XL U175 ( .A(n4), .B(n13), .Y(n12) );
  INVXL U176 ( .A(n14), .Y(n13) );
  NOR2XL U177 ( .A(B[1]), .B(B[0]), .Y(n109) );
  NAND2XL U178 ( .A(n51), .B(n43), .Y(n42) );
  CLKINVX2 U179 ( .A(n93), .Y(n92) );
  INVXL U180 ( .A(n88), .Y(n87) );
  NOR2XL U181 ( .A(B[19]), .B(B[18]), .Y(n53) );
  NOR2BXL U182 ( .AN(n27), .B(B[26]), .Y(n24) );
  NOR2XL U183 ( .A(n4), .B(B[28]), .Y(n17) );
  NOR2X6 U184 ( .A(n50), .B(n36), .Y(n3) );
  NOR2XL U185 ( .A(B[27]), .B(B[26]), .Y(n21) );
  NOR2BXL U186 ( .AN(n43), .B(B[22]), .Y(n40) );
  XNOR2X1 U187 ( .A(n57), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U188 ( .A(n212), .B(n58), .Y(n57) );
  INVXL U189 ( .A(n59), .Y(n58) );
  CLKINVX1 U190 ( .A(n109), .Y(n108) );
  NOR2X2 U191 ( .A(n79), .B(n65), .Y(n64) );
  NAND2X1 U192 ( .A(n72), .B(n66), .Y(n65) );
  NOR2X1 U193 ( .A(n92), .B(n71), .Y(n70) );
  NAND2XL U194 ( .A(n80), .B(n72), .Y(n71) );
  NOR2X1 U195 ( .A(n92), .B(n68), .Y(n67) );
  NAND2XL U196 ( .A(n69), .B(n80), .Y(n68) );
  NOR2X1 U197 ( .A(n92), .B(n76), .Y(n75) );
  NAND2XL U198 ( .A(n80), .B(n77), .Y(n76) );
  NOR2X1 U199 ( .A(n92), .B(n87), .Y(n86) );
  NOR2XL U200 ( .A(n212), .B(n34), .Y(n33) );
  CLKINVX1 U201 ( .A(n3), .Y(n34) );
  NOR2XL U202 ( .A(n212), .B(n11), .Y(n10) );
  NAND2X1 U203 ( .A(n3), .B(n12), .Y(n11) );
  NOR2XL U204 ( .A(n212), .B(n26), .Y(n25) );
  NOR2XL U205 ( .A(n212), .B(n19), .Y(n18) );
  NOR2X1 U206 ( .A(n212), .B(n42), .Y(n41) );
  NAND2X1 U207 ( .A(n106), .B(n109), .Y(n105) );
  NOR2X1 U208 ( .A(n213), .B(B[3]), .Y(n106) );
  NAND2X1 U209 ( .A(n37), .B(n43), .Y(n36) );
  NAND2X1 U210 ( .A(n53), .B(n59), .Y(n50) );
  NOR2XL U211 ( .A(n212), .B(n55), .Y(n54) );
  CLKINVX1 U212 ( .A(B[18]), .Y(n56) );
  NOR2X1 U213 ( .A(n92), .B(n84), .Y(n83) );
  NAND2XL U214 ( .A(n88), .B(n85), .Y(n84) );
  XNOR2X1 U215 ( .A(n5), .B(B[31]), .Y(DIFF[31]) );
  NOR2XL U216 ( .A(n212), .B(n6), .Y(n5) );
  NAND2XL U217 ( .A(n3), .B(n7), .Y(n6) );
  NOR2X1 U218 ( .A(n4), .B(n8), .Y(n7) );
  NOR2XL U219 ( .A(n212), .B(n31), .Y(n30) );
  NAND2XL U220 ( .A(n3), .B(n32), .Y(n31) );
  CLKINVX1 U221 ( .A(B[24]), .Y(n32) );
  NOR2XL U222 ( .A(n212), .B(n23), .Y(n22) );
  NAND2X1 U223 ( .A(n3), .B(n24), .Y(n23) );
  NOR2XL U224 ( .A(n212), .B(n16), .Y(n15) );
  NAND2X1 U225 ( .A(n3), .B(n17), .Y(n16) );
  NOR2XL U226 ( .A(n212), .B(n39), .Y(n38) );
  NAND2X1 U227 ( .A(n40), .B(n51), .Y(n39) );
  NOR2XL U228 ( .A(n212), .B(n47), .Y(n46) );
  NAND2X1 U229 ( .A(n51), .B(n48), .Y(n47) );
  NAND2X1 U230 ( .A(n14), .B(n9), .Y(n8) );
  INVXL U231 ( .A(B[30]), .Y(n9) );
  NOR2X1 U232 ( .A(B[25]), .B(B[24]), .Y(n27) );
  NAND2X2 U233 ( .A(n27), .B(n21), .Y(n4) );
  NOR2XL U234 ( .A(B[15]), .B(B[14]), .Y(n66) );
  NOR2X4 U235 ( .A(n94), .B(n105), .Y(n93) );
  NAND2X1 U236 ( .A(n99), .B(n95), .Y(n94) );
  NAND2X1 U237 ( .A(n97), .B(n104), .Y(n96) );
  XNOR2XL U238 ( .A(n10), .B(B[30]), .Y(DIFF[30]) );
  XNOR2XL U239 ( .A(n33), .B(B[24]), .Y(DIFF[24]) );
  XNOR2XL U240 ( .A(n67), .B(B[15]), .Y(DIFF[15]) );
  XNOR2XL U241 ( .A(n30), .B(B[25]), .Y(DIFF[25]) );
  XNOR2XL U242 ( .A(n75), .B(B[13]), .Y(DIFF[13]) );
  XNOR2XL U243 ( .A(n49), .B(B[20]), .Y(DIFF[20]) );
  XNOR2XL U244 ( .A(n25), .B(B[26]), .Y(DIFF[26]) );
  XNOR2XL U245 ( .A(n18), .B(B[28]), .Y(DIFF[28]) );
  XOR2XL U246 ( .A(B[1]), .B(B[0]), .Y(DIFF[1]) );
  XOR2XL U247 ( .A(n108), .B(n213), .Y(DIFF[2]) );
  XNOR2XL U248 ( .A(n107), .B(B[3]), .Y(DIFF[3]) );
  XNOR2XL U249 ( .A(n104), .B(n214), .Y(DIFF[4]) );
  XOR2XL U250 ( .A(n102), .B(B[5]), .Y(DIFF[5]) );
  XNOR2XL U251 ( .A(n15), .B(B[29]), .Y(DIFF[29]) );
  NOR2XL U252 ( .A(B[28]), .B(B[29]), .Y(n14) );
  XOR2XL U253 ( .A(n96), .B(B[7]), .Y(DIFF[7]) );
  XNOR2XL U254 ( .A(n86), .B(B[10]), .Y(DIFF[10]) );
  INVXL U255 ( .A(B[10]), .Y(n85) );
  NOR2XL U256 ( .A(B[10]), .B(B[11]), .Y(n82) );
  XNOR2XL U257 ( .A(n91), .B(B[9]), .Y(DIFF[9]) );
  NOR2XL U258 ( .A(B[8]), .B(B[9]), .Y(n88) );
  NOR2XL U259 ( .A(B[23]), .B(B[22]), .Y(n37) );
  XOR2XL U260 ( .A(n212), .B(B[16]), .Y(DIFF[16]) );
  NOR2XL U261 ( .A(n212), .B(B[16]), .Y(n62) );
  XNOR2XL U262 ( .A(n22), .B(B[27]), .Y(DIFF[27]) );
  XNOR2XL U263 ( .A(n83), .B(B[11]), .Y(DIFF[11]) );
  NOR2XL U264 ( .A(B[16]), .B(B[17]), .Y(n59) );
  NAND2XL U265 ( .A(n59), .B(n56), .Y(n55) );
  XNOR2XL U266 ( .A(n54), .B(B[19]), .Y(DIFF[19]) );
  XNOR2XL U267 ( .A(n41), .B(B[22]), .Y(DIFF[22]) );
  XNOR2XL U268 ( .A(n46), .B(B[21]), .Y(DIFF[21]) );
  XNOR2XL U269 ( .A(n62), .B(B[17]), .Y(DIFF[17]) );
endmodule


module ALU_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388;

  NOR2X2 U764 ( .A(B[9]), .B(n129), .Y(n90) );
  INVX2 U765 ( .A(A[19]), .Y(n139) );
  INVX4 U766 ( .A(A[12]), .Y(n132) );
  OAI21X2 U767 ( .A0(n70), .A1(n73), .B0(n71), .Y(n69) );
  CLKINVX4 U768 ( .A(A[9]), .Y(n129) );
  CLKBUFX2 U769 ( .A(B[1]), .Y(n1384) );
  OAI21X4 U770 ( .A0(n84), .A1(n87), .B0(n85), .Y(n83) );
  NAND2X2 U771 ( .A(B[10]), .B(n130), .Y(n87) );
  CLKINVX8 U772 ( .A(A[11]), .Y(n131) );
  NAND2X1 U773 ( .A(B[9]), .B(n129), .Y(n91) );
  INVX2 U774 ( .A(A[8]), .Y(n128) );
  NAND2X2 U775 ( .A(n1385), .B(n122), .Y(n115) );
  CLKINVX2 U776 ( .A(A[24]), .Y(n144) );
  NOR2X4 U777 ( .A(n23), .B(n25), .Y(n21) );
  NOR2X2 U778 ( .A(B[28]), .B(n148), .Y(n17) );
  NOR2X2 U779 ( .A(B[20]), .B(n140), .Y(n47) );
  OAI21X2 U780 ( .A0(n90), .A1(n93), .B0(n91), .Y(n89) );
  INVX4 U781 ( .A(A[3]), .Y(n123) );
  NOR2X4 U782 ( .A(n78), .B(n1383), .Y(n74) );
  NOR2X2 U783 ( .A(B[12]), .B(n132), .Y(n78) );
  NOR2X6 U784 ( .A(n5), .B(n19), .Y(n3) );
  CLKINVX3 U785 ( .A(A[28]), .Y(n148) );
  NOR2X8 U786 ( .A(B[31]), .B(n151), .Y(n1379) );
  NAND2X1 U787 ( .A(B[7]), .B(n127), .Y(n100) );
  NAND2X1 U788 ( .A(B[0]), .B(n120), .Y(n119) );
  INVX1 U789 ( .A(A[0]), .Y(n120) );
  OAI31X4 U790 ( .A0(n1380), .A1(n29), .A2(A[24]), .B0(n30), .Y(n28) );
  CLKINVX1 U791 ( .A(B[24]), .Y(n1380) );
  OAI21X4 U792 ( .A0(n112), .A1(n115), .B0(n113), .Y(n111) );
  NAND2X1 U793 ( .A(B[14]), .B(n134), .Y(n73) );
  NOR2X2 U794 ( .A(B[6]), .B(n126), .Y(n101) );
  CLKINVX2 U795 ( .A(A[14]), .Y(n134) );
  CLKBUFX6 U796 ( .A(B[5]), .Y(n1388) );
  NOR2X2 U797 ( .A(B[10]), .B(n130), .Y(n86) );
  NOR2X4 U798 ( .A(n1382), .B(n147), .Y(n1381) );
  INVX8 U799 ( .A(A[27]), .Y(n147) );
  NOR2X6 U800 ( .A(n1382), .B(n147), .Y(n23) );
  NAND2X1 U801 ( .A(B[25]), .B(n145), .Y(n30) );
  CLKINVX6 U802 ( .A(A[25]), .Y(n145) );
  OAI21X4 U803 ( .A0(n26), .A1(n1381), .B0(n24), .Y(n22) );
  NAND2X1 U804 ( .A(B[26]), .B(n146), .Y(n26) );
  NOR2X4 U805 ( .A(n1385), .B(n122), .Y(n114) );
  AOI21X4 U806 ( .A0(n104), .A1(n97), .B0(n98), .Y(n96) );
  OAI21X2 U807 ( .A0(n99), .A1(n102), .B0(n100), .Y(n98) );
  CLKBUFX3 U808 ( .A(B[2]), .Y(n1385) );
  INVX3 U809 ( .A(A[16]), .Y(n136) );
  OAI21X4 U810 ( .A0(n59), .A1(n62), .B0(n60), .Y(n58) );
  NOR2X4 U811 ( .A(B[17]), .B(n137), .Y(n59) );
  NAND2X1 U812 ( .A(B[16]), .B(n136), .Y(n62) );
  NOR2X2 U813 ( .A(B[26]), .B(n146), .Y(n25) );
  NOR2X4 U814 ( .A(n17), .B(n15), .Y(n13) );
  NOR2X6 U815 ( .A(B[29]), .B(n149), .Y(n15) );
  NOR2X2 U816 ( .A(B[30]), .B(n150), .Y(n11) );
  NOR2X4 U817 ( .A(n99), .B(n101), .Y(n97) );
  NOR2X4 U818 ( .A(B[7]), .B(n127), .Y(n99) );
  INVX4 U819 ( .A(A[6]), .Y(n126) );
  AOI21X4 U820 ( .A0(n89), .A1(n82), .B0(n83), .Y(n81) );
  NOR2X4 U821 ( .A(n86), .B(n84), .Y(n82) );
  NOR2X4 U822 ( .A(B[23]), .B(n143), .Y(n39) );
  INVX2 U823 ( .A(A[23]), .Y(n143) );
  NAND2X1 U824 ( .A(B[31]), .B(n151), .Y(n10) );
  NOR2X2 U825 ( .A(B[18]), .B(n138), .Y(n55) );
  NOR2X8 U826 ( .A(B[19]), .B(n139), .Y(n53) );
  INVX6 U827 ( .A(A[18]), .Y(n138) );
  NAND2X2 U828 ( .A(B[20]), .B(n140), .Y(n48) );
  NOR2X1 U829 ( .A(B[24]), .B(n144), .Y(n31) );
  OAI21X4 U830 ( .A0(n15), .A1(n18), .B0(n16), .Y(n14) );
  NAND2X2 U831 ( .A(B[28]), .B(n148), .Y(n18) );
  NAND2X2 U832 ( .A(B[29]), .B(n149), .Y(n16) );
  NOR2X6 U833 ( .A(n1388), .B(n125), .Y(n105) );
  INVX6 U834 ( .A(A[5]), .Y(n125) );
  NOR2X4 U835 ( .A(n107), .B(n105), .Y(n103) );
  NOR2X2 U836 ( .A(n1387), .B(n124), .Y(n107) );
  NOR2X4 U837 ( .A(B[11]), .B(n131), .Y(n84) );
  NAND2X1 U838 ( .A(B[11]), .B(n131), .Y(n85) );
  CLKINVX2 U839 ( .A(A[4]), .Y(n124) );
  OAI21X2 U840 ( .A0(n105), .A1(n108), .B0(n106), .Y(n104) );
  NAND2X2 U841 ( .A(n1387), .B(n124), .Y(n108) );
  BUFX20 U842 ( .A(B[27]), .Y(n1382) );
  INVX3 U843 ( .A(A[29]), .Y(n149) );
  CLKINVX3 U844 ( .A(A[13]), .Y(n133) );
  INVX6 U845 ( .A(A[26]), .Y(n146) );
  CLKINVX4 U846 ( .A(A[20]), .Y(n140) );
  OAI21X4 U847 ( .A0(n50), .A1(n35), .B0(n36), .Y(n34) );
  AOI21X4 U848 ( .A0(n44), .A1(n37), .B0(n38), .Y(n36) );
  NOR2X4 U849 ( .A(n39), .B(n41), .Y(n37) );
  NOR2X6 U850 ( .A(n80), .B(n66), .Y(n64) );
  NAND2X1 U851 ( .A(B[8]), .B(n128), .Y(n93) );
  NOR2X1 U852 ( .A(B[13]), .B(n133), .Y(n76) );
  NAND2X1 U853 ( .A(B[19]), .B(n139), .Y(n54) );
  NAND2X2 U854 ( .A(B[30]), .B(n150), .Y(n12) );
  NOR2X2 U855 ( .A(n1386), .B(n123), .Y(n112) );
  AOI21X4 U856 ( .A0(n28), .A1(n21), .B0(n22), .Y(n20) );
  OAI21X4 U857 ( .A0(n20), .A1(n5), .B0(n6), .Y(n4) );
  NOR2X4 U858 ( .A(B[25]), .B(n145), .Y(n29) );
  NOR2X2 U859 ( .A(B[14]), .B(n134), .Y(n72) );
  NAND2X6 U860 ( .A(n7), .B(n13), .Y(n5) );
  OAI21X2 U861 ( .A0(n39), .A1(n42), .B0(n40), .Y(n38) );
  OAI21X1 U862 ( .A0(n45), .A1(n48), .B0(n46), .Y(n44) );
  CLKINVX8 U863 ( .A(A[21]), .Y(n141) );
  INVX6 U864 ( .A(A[30]), .Y(n150) );
  NAND2X2 U865 ( .A(n103), .B(n97), .Y(n95) );
  AOI21X4 U866 ( .A0(n110), .A1(n116), .B0(n111), .Y(n109) );
  OAI21X4 U867 ( .A0(n81), .A1(n66), .B0(n67), .Y(n65) );
  AOI21X4 U868 ( .A0(n75), .A1(n68), .B0(n69), .Y(n67) );
  OAI21X4 U869 ( .A0(n63), .A1(n1), .B0(n2), .Y(GE_LT_GT_LE) );
  AOI21X4 U870 ( .A0(n34), .A1(n3), .B0(n4), .Y(n2) );
  OAI21X4 U871 ( .A0(n109), .A1(n95), .B0(n96), .Y(n94) );
  AOI21X4 U872 ( .A0(n14), .A1(n7), .B0(n8), .Y(n6) );
  OAI21X2 U873 ( .A0(n1379), .A1(n12), .B0(n10), .Y(n8) );
  NAND2X1 U874 ( .A(B[21]), .B(n141), .Y(n46) );
  NAND2X4 U875 ( .A(n51), .B(n57), .Y(n49) );
  NOR2X4 U876 ( .A(n1379), .B(n11), .Y(n7) );
  AOI21X4 U877 ( .A0(n94), .A1(n64), .B0(n65), .Y(n63) );
  NAND2X4 U878 ( .A(n27), .B(n21), .Y(n19) );
  NOR2X1 U879 ( .A(n29), .B(n31), .Y(n27) );
  NAND2X2 U880 ( .A(B[12]), .B(n132), .Y(n79) );
  AOI21X4 U881 ( .A0(n58), .A1(n51), .B0(n52), .Y(n50) );
  NAND2X2 U882 ( .A(n1382), .B(n147), .Y(n24) );
  OAI21X4 U883 ( .A0(n117), .A1(n119), .B0(n118), .Y(n116) );
  NOR2X4 U884 ( .A(n1384), .B(n121), .Y(n117) );
  NAND2X2 U885 ( .A(n1384), .B(n121), .Y(n118) );
  NOR2X4 U886 ( .A(n61), .B(n59), .Y(n57) );
  NOR2X2 U887 ( .A(B[16]), .B(n136), .Y(n61) );
  NAND2X1 U888 ( .A(B[22]), .B(n142), .Y(n42) );
  NOR2X2 U889 ( .A(n114), .B(n112), .Y(n110) );
  NOR2X2 U890 ( .A(B[22]), .B(n142), .Y(n41) );
  NOR2X1 U891 ( .A(B[8]), .B(n128), .Y(n92) );
  NOR2X4 U892 ( .A(B[21]), .B(n141), .Y(n45) );
  OAI21X4 U893 ( .A0(n1383), .A1(n79), .B0(n77), .Y(n75) );
  NAND2X2 U894 ( .A(n3), .B(n33), .Y(n1) );
  NOR2X4 U895 ( .A(n49), .B(n35), .Y(n33) );
  NAND2X6 U896 ( .A(n74), .B(n68), .Y(n66) );
  NOR2X2 U897 ( .A(B[15]), .B(n135), .Y(n70) );
  INVX4 U898 ( .A(A[15]), .Y(n135) );
  NAND2X2 U899 ( .A(n88), .B(n82), .Y(n80) );
  NOR2X1 U900 ( .A(n92), .B(n90), .Y(n88) );
  NAND2X4 U901 ( .A(n37), .B(n43), .Y(n35) );
  NOR2X4 U902 ( .A(n45), .B(n47), .Y(n43) );
  CLKINVX8 U903 ( .A(A[7]), .Y(n127) );
  BUFX4 U904 ( .A(n76), .Y(n1383) );
  NAND2X1 U905 ( .A(n1388), .B(n125), .Y(n106) );
  CLKINVX6 U906 ( .A(A[31]), .Y(n151) );
  NOR2X4 U907 ( .A(n53), .B(n55), .Y(n51) );
  OAI21X2 U908 ( .A0(n53), .A1(n56), .B0(n54), .Y(n52) );
  NOR2X4 U909 ( .A(n70), .B(n72), .Y(n68) );
  CLKINVX8 U910 ( .A(A[1]), .Y(n121) );
  NAND2XL U911 ( .A(B[23]), .B(n143), .Y(n40) );
  NAND2XL U912 ( .A(n1386), .B(n123), .Y(n113) );
  NAND2XL U913 ( .A(B[15]), .B(n135), .Y(n71) );
  CLKINVX1 U914 ( .A(A[17]), .Y(n137) );
  CLKINVX1 U915 ( .A(A[2]), .Y(n122) );
  CLKINVX1 U916 ( .A(A[22]), .Y(n142) );
  CLKINVX1 U917 ( .A(A[10]), .Y(n130) );
  CLKBUFX3 U918 ( .A(B[4]), .Y(n1387) );
  CLKBUFX3 U919 ( .A(B[3]), .Y(n1386) );
  NAND2XL U920 ( .A(B[13]), .B(n133), .Y(n77) );
  NAND2XL U921 ( .A(B[6]), .B(n126), .Y(n102) );
  NAND2X1 U922 ( .A(B[18]), .B(n138), .Y(n56) );
  NAND2X1 U923 ( .A(B[17]), .B(n137), .Y(n60) );
endmodule


module ALU_DW01_add_8 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n100, n101, n102, n103, n104, n105, n107, n110,
         n111, n112, n113, n114, n116, n117, n118, n119, n120, n121, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n138, n139, n140, n141, n142, n143, n145, n148, n149, n150, n151,
         n152, n154, n155, n156, n157, n158, n159, n160, n161, n164, n165,
         n166, n167, n168, n169, n170, n172, n173, n174, n175, n176, n177,
         n178, n179, n184, n185, n186, n187, n188, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n206,
         n207, n208, n209, n210, n211, n213, n216, n217, n218, n219, n220,
         n222, n223, n224, n225, n226, n227, n228, n229, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n271, n272, n273, n274,
         n276, n279, n280, n281, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n438, n439, n440, n441,
         n442, n443, n444;

  AOI21X1 U369 ( .A0(n274), .A1(n261), .B0(n262), .Y(n260) );
  NOR2X4 U370 ( .A(n226), .B(n192), .Y(n190) );
  INVX1 U371 ( .A(n247), .Y(n245) );
  NAND2XL U372 ( .A(n4), .B(n64), .Y(n62) );
  OAI21X2 U373 ( .A0(n184), .A1(n188), .B0(n185), .Y(n179) );
  INVX3 U374 ( .A(n159), .Y(n161) );
  INVX1 U375 ( .A(n285), .Y(n283) );
  INVX1 U376 ( .A(n187), .Y(n316) );
  AND2XL U377 ( .A(n4), .B(n42), .Y(n438) );
  XNOR2X4 U378 ( .A(n236), .B(n27), .Y(SUM[11]) );
  BUFX20 U379 ( .A(n2), .Y(n444) );
  XNOR2X4 U380 ( .A(n61), .B(n8), .Y(SUM[30]) );
  NOR2X2 U381 ( .A(B[8]), .B(A[8]), .Y(n255) );
  NAND2X4 U382 ( .A(n246), .B(n232), .Y(n226) );
  NOR2X2 U383 ( .A(n241), .B(n234), .Y(n232) );
  NOR2X4 U384 ( .A(n255), .B(n252), .Y(n246) );
  NOR2X4 U385 ( .A(n187), .B(n184), .Y(n178) );
  NOR2X2 U386 ( .A(B[16]), .B(A[16]), .Y(n187) );
  NAND2X2 U387 ( .A(n178), .B(n314), .Y(n169) );
  NAND2X2 U388 ( .A(n178), .B(n164), .Y(n158) );
  INVX3 U389 ( .A(n178), .Y(n176) );
  XNOR2X4 U390 ( .A(n92), .B(n11), .Y(SUM[27]) );
  XNOR2X4 U391 ( .A(n81), .B(n10), .Y(SUM[28]) );
  OAI21X4 U392 ( .A0(n444), .A1(n82), .B0(n83), .Y(n81) );
  NOR2X2 U393 ( .A(B[30]), .B(A[30]), .Y(n59) );
  AOI21X2 U394 ( .A0(n3), .A1(n53), .B0(n54), .Y(n52) );
  CLKINVX12 U395 ( .A(n441), .Y(n3) );
  OAI21X1 U396 ( .A0(n5), .A1(n55), .B0(n56), .Y(n54) );
  CLKINVX6 U397 ( .A(n173), .Y(n314) );
  NOR2X2 U398 ( .A(B[18]), .B(A[18]), .Y(n173) );
  OAI21X1 U399 ( .A0(n444), .A1(n158), .B0(n159), .Y(n157) );
  AOI21X2 U400 ( .A0(n179), .A1(n164), .B0(n165), .Y(n159) );
  CLKINVX3 U401 ( .A(n158), .Y(n160) );
  XNOR2X4 U402 ( .A(n101), .B(n12), .Y(SUM[26]) );
  AOI21X4 U403 ( .A0(n258), .A1(n190), .B0(n191), .Y(n2) );
  NAND2X1 U404 ( .A(B[6]), .B(A[6]), .Y(n271) );
  OAI21X1 U405 ( .A0(n263), .A1(n271), .B0(n264), .Y(n262) );
  AOI21XL U406 ( .A0(n3), .A1(n64), .B0(n65), .Y(n63) );
  NOR2X1 U407 ( .A(n6), .B(n66), .Y(n64) );
  OAI21X2 U408 ( .A0(n252), .A1(n256), .B0(n253), .Y(n247) );
  NAND2X2 U409 ( .A(n324), .B(n256), .Y(n30) );
  OAI21X1 U410 ( .A0(n257), .A1(n255), .B0(n256), .Y(n254) );
  NAND2X1 U411 ( .A(B[8]), .B(A[8]), .Y(n256) );
  AOI21X1 U412 ( .A0(n247), .A1(n322), .B0(n240), .Y(n238) );
  OAI21X2 U413 ( .A0(n279), .A1(n285), .B0(n280), .Y(n274) );
  NAND2X2 U414 ( .A(n328), .B(n285), .Y(n34) );
  NAND2X2 U415 ( .A(B[4]), .B(A[4]), .Y(n285) );
  INVX3 U416 ( .A(n274), .Y(n276) );
  AOI21X1 U417 ( .A0(n286), .A1(n273), .B0(n274), .Y(n272) );
  XNOR2X4 U418 ( .A(n130), .B(n15), .Y(SUM[23]) );
  XNOR2X4 U419 ( .A(n198), .B(n23), .Y(SUM[15]) );
  NAND2X2 U420 ( .A(B[2]), .B(A[2]), .Y(n294) );
  XNOR2X4 U421 ( .A(n207), .B(n24), .Y(SUM[14]) );
  NAND2X4 U422 ( .A(B[26]), .B(A[26]), .Y(n100) );
  XNOR2X4 U423 ( .A(n218), .B(n25), .Y(SUM[13]) );
  OAI21X4 U424 ( .A0(n257), .A1(n219), .B0(n220), .Y(n218) );
  XNOR2X4 U425 ( .A(n139), .B(n16), .Y(SUM[22]) );
  XNOR2X4 U426 ( .A(n150), .B(n17), .Y(SUM[21]) );
  OAI21X2 U427 ( .A0(n444), .A1(n151), .B0(n152), .Y(n150) );
  OAI21X1 U428 ( .A0(n290), .A1(n294), .B0(n291), .Y(n289) );
  NOR2X6 U429 ( .A(n117), .B(n110), .Y(n104) );
  NOR2X2 U430 ( .A(B[25]), .B(A[25]), .Y(n110) );
  NOR2X2 U431 ( .A(B[24]), .B(A[24]), .Y(n117) );
  XNOR2X4 U432 ( .A(n72), .B(n9), .Y(SUM[29]) );
  OAI21X2 U433 ( .A0(n444), .A1(n73), .B0(n74), .Y(n72) );
  OAI2BB1X4 U434 ( .A0N(n438), .A1N(n439), .B0(n41), .Y(SUM[32]) );
  INVXL U435 ( .A(n2), .Y(n439) );
  NAND2X2 U436 ( .A(B[9]), .B(A[9]), .Y(n253) );
  NOR2X2 U437 ( .A(B[9]), .B(A[9]), .Y(n252) );
  NAND2X2 U438 ( .A(B[1]), .B(A[1]), .Y(n298) );
  NOR2X2 U439 ( .A(B[1]), .B(A[1]), .Y(n297) );
  NAND2X2 U440 ( .A(B[16]), .B(A[16]), .Y(n188) );
  NOR2X2 U441 ( .A(B[17]), .B(A[17]), .Y(n184) );
  NAND2X2 U442 ( .A(B[24]), .B(A[24]), .Y(n118) );
  OAI21X4 U443 ( .A0(n227), .A1(n192), .B0(n193), .Y(n191) );
  NAND2X2 U444 ( .A(n142), .B(n126), .Y(n124) );
  CLKXOR2X2 U445 ( .A(n443), .B(n35), .Y(SUM[3]) );
  CLKINVX8 U446 ( .A(n440), .Y(n4) );
  AOI21XL U447 ( .A0(n3), .A1(n42), .B0(n43), .Y(n41) );
  NAND2X1 U448 ( .A(n201), .B(n228), .Y(n199) );
  INVX1 U449 ( .A(n287), .Y(n286) );
  OAI21X1 U450 ( .A0(n297), .A1(n300), .B0(n298), .Y(n296) );
  NOR2X2 U451 ( .A(n155), .B(n148), .Y(n142) );
  NOR2X2 U452 ( .A(n223), .B(n216), .Y(n210) );
  NOR2X2 U453 ( .A(n77), .B(n70), .Y(n68) );
  OA21XL U454 ( .A0(n295), .A1(n293), .B0(n294), .Y(n443) );
  INVXL U455 ( .A(n297), .Y(n331) );
  OR2X4 U456 ( .A(n158), .B(n124), .Y(n440) );
  NOR2X2 U457 ( .A(n6), .B(n55), .Y(n53) );
  CLKINVX3 U458 ( .A(n226), .Y(n228) );
  INVXL U459 ( .A(n6), .Y(n84) );
  NAND2X2 U460 ( .A(n210), .B(n194), .Y(n192) );
  NOR2XL U461 ( .A(n6), .B(n44), .Y(n42) );
  AOI21X1 U462 ( .A0(n3), .A1(n84), .B0(n85), .Y(n83) );
  INVXL U463 ( .A(n5), .Y(n85) );
  NAND2X2 U464 ( .A(n68), .B(n57), .Y(n55) );
  INVXL U465 ( .A(n227), .Y(n229) );
  AOI21XL U466 ( .A0(n3), .A1(n104), .B0(n105), .Y(n103) );
  AOI21XL U467 ( .A0(n161), .A1(n142), .B0(n143), .Y(n141) );
  AOI21XL U468 ( .A0(n229), .A1(n210), .B0(n211), .Y(n209) );
  INVXL U469 ( .A(n69), .Y(n67) );
  INVXL U470 ( .A(n179), .Y(n177) );
  NAND2XL U471 ( .A(n246), .B(n322), .Y(n237) );
  NAND2XL U472 ( .A(n133), .B(n160), .Y(n131) );
  OAI21X4 U473 ( .A0(n287), .A1(n259), .B0(n260), .Y(n258) );
  NAND2X2 U474 ( .A(n273), .B(n261), .Y(n259) );
  OA21X4 U475 ( .A0(n159), .A1(n124), .B0(n125), .Y(n441) );
  XOR2X4 U476 ( .A(n442), .B(n7), .Y(SUM[31]) );
  OA21X4 U477 ( .A0(n444), .A1(n51), .B0(n52), .Y(n442) );
  NOR2BXL U478 ( .AN(n210), .B(n203), .Y(n201) );
  INVXL U479 ( .A(n242), .Y(n240) );
  NOR2BXL U480 ( .AN(n142), .B(n135), .Y(n133) );
  NOR2BXL U481 ( .AN(n104), .B(n97), .Y(n95) );
  NOR2XL U482 ( .A(n6), .B(n77), .Y(n75) );
  CLKXOR2X1 U483 ( .A(n295), .B(n36), .Y(SUM[2]) );
  XOR2X1 U484 ( .A(n37), .B(n300), .Y(SUM[1]) );
  NOR2XL U485 ( .A(B[12]), .B(A[12]), .Y(n223) );
  NOR2XL U486 ( .A(B[20]), .B(A[20]), .Y(n155) );
  NAND2XL U487 ( .A(B[12]), .B(A[12]), .Y(n224) );
  NAND2XL U488 ( .A(B[20]), .B(A[20]), .Y(n156) );
  NAND2X2 U489 ( .A(B[0]), .B(A[0]), .Y(n300) );
  NAND2XL U490 ( .A(B[18]), .B(A[18]), .Y(n174) );
  NAND2XL U491 ( .A(B[14]), .B(A[14]), .Y(n206) );
  NOR2XL U492 ( .A(B[10]), .B(A[10]), .Y(n241) );
  NOR2XL U493 ( .A(B[4]), .B(A[4]), .Y(n284) );
  NOR2X1 U494 ( .A(B[14]), .B(A[14]), .Y(n203) );
  NOR2X1 U495 ( .A(B[6]), .B(A[6]), .Y(n268) );
  NOR2X1 U496 ( .A(B[13]), .B(A[13]), .Y(n216) );
  NOR2X1 U497 ( .A(B[21]), .B(A[21]), .Y(n148) );
  NOR2X1 U498 ( .A(B[5]), .B(A[5]), .Y(n279) );
  NAND2XL U499 ( .A(B[13]), .B(A[13]), .Y(n217) );
  NAND2XL U500 ( .A(B[21]), .B(A[21]), .Y(n149) );
  NAND2XL U501 ( .A(B[5]), .B(A[5]), .Y(n280) );
  NOR2X1 U502 ( .A(B[23]), .B(A[23]), .Y(n128) );
  NOR2X1 U503 ( .A(B[11]), .B(A[11]), .Y(n234) );
  NOR2X1 U504 ( .A(B[19]), .B(A[19]), .Y(n166) );
  NOR2X1 U505 ( .A(B[15]), .B(A[15]), .Y(n196) );
  NOR2X1 U506 ( .A(B[27]), .B(A[27]), .Y(n90) );
  NOR2X1 U507 ( .A(B[7]), .B(A[7]), .Y(n263) );
  NOR2X1 U508 ( .A(B[3]), .B(A[3]), .Y(n290) );
  NAND2XL U509 ( .A(B[25]), .B(A[25]), .Y(n111) );
  NAND2XL U510 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U511 ( .A(B[2]), .B(A[2]), .Y(n293) );
  NAND2XL U512 ( .A(B[11]), .B(A[11]), .Y(n235) );
  NAND2XL U513 ( .A(B[15]), .B(A[15]), .Y(n197) );
  NAND2XL U514 ( .A(B[19]), .B(A[19]), .Y(n167) );
  NAND2XL U515 ( .A(B[3]), .B(A[3]), .Y(n291) );
  NAND2XL U516 ( .A(B[7]), .B(A[7]), .Y(n264) );
  NAND2XL U517 ( .A(B[28]), .B(A[28]), .Y(n80) );
  NOR2X1 U518 ( .A(B[28]), .B(A[28]), .Y(n77) );
  NAND2XL U519 ( .A(B[30]), .B(A[30]), .Y(n60) );
  NAND2XL U520 ( .A(B[22]), .B(A[22]), .Y(n138) );
  NOR2X1 U521 ( .A(B[22]), .B(A[22]), .Y(n135) );
  NOR2X1 U522 ( .A(B[26]), .B(A[26]), .Y(n97) );
  NOR2X1 U523 ( .A(B[29]), .B(A[29]), .Y(n70) );
  NAND2XL U524 ( .A(B[29]), .B(A[29]), .Y(n71) );
  NOR2X1 U525 ( .A(B[31]), .B(A[31]), .Y(n48) );
  NAND2XL U526 ( .A(B[23]), .B(A[23]), .Y(n129) );
  NAND2XL U527 ( .A(B[27]), .B(A[27]), .Y(n91) );
  NAND2XL U528 ( .A(B[31]), .B(A[31]), .Y(n49) );
  NAND2BXL U529 ( .AN(n299), .B(n300), .Y(n38) );
  NAND2X1 U530 ( .A(n4), .B(n84), .Y(n82) );
  NAND2X1 U531 ( .A(n4), .B(n53), .Y(n51) );
  INVX3 U532 ( .A(n258), .Y(n257) );
  NAND2X2 U533 ( .A(n104), .B(n88), .Y(n6) );
  OAI21XL U534 ( .A0(n5), .A1(n66), .B0(n67), .Y(n65) );
  CLKINVX1 U535 ( .A(n68), .Y(n66) );
  CLKINVX1 U536 ( .A(n296), .Y(n295) );
  NAND2X1 U537 ( .A(n68), .B(n46), .Y(n44) );
  NAND2XL U538 ( .A(n228), .B(n320), .Y(n219) );
  NAND2XL U539 ( .A(n160), .B(n312), .Y(n151) );
  NAND2XL U540 ( .A(n4), .B(n308), .Y(n113) );
  NAND2XL U541 ( .A(n228), .B(n210), .Y(n208) );
  NAND2XL U542 ( .A(n160), .B(n142), .Y(n140) );
  NAND2XL U543 ( .A(n4), .B(n104), .Y(n102) );
  NAND2XL U544 ( .A(n4), .B(n75), .Y(n73) );
  NAND2XL U545 ( .A(n4), .B(n95), .Y(n93) );
  CLKINVX1 U546 ( .A(n3), .Y(n121) );
  AOI21X2 U547 ( .A0(n105), .A1(n88), .B0(n89), .Y(n5) );
  OAI21XL U548 ( .A0(n90), .A1(n100), .B0(n91), .Y(n89) );
  AOI21X2 U549 ( .A0(n247), .A1(n232), .B0(n233), .Y(n227) );
  OAI21XL U550 ( .A0(n234), .A1(n242), .B0(n235), .Y(n233) );
  OAI21XL U551 ( .A0(n166), .A1(n174), .B0(n167), .Y(n165) );
  OAI21X1 U552 ( .A0(n216), .A1(n224), .B0(n217), .Y(n211) );
  OAI21X1 U553 ( .A0(n110), .A1(n118), .B0(n111), .Y(n105) );
  NOR2X1 U554 ( .A(n268), .B(n263), .Y(n261) );
  AOI21X1 U555 ( .A0(n296), .A1(n288), .B0(n289), .Y(n287) );
  NOR2X1 U556 ( .A(n293), .B(n290), .Y(n288) );
  AOI21X1 U557 ( .A0(n211), .A1(n194), .B0(n195), .Y(n193) );
  OAI21XL U558 ( .A0(n196), .A1(n206), .B0(n197), .Y(n195) );
  AOI21X1 U559 ( .A0(n69), .A1(n57), .B0(n58), .Y(n56) );
  CLKINVX1 U560 ( .A(n60), .Y(n58) );
  NAND2X1 U561 ( .A(n301), .B(n49), .Y(n7) );
  CLKINVX1 U562 ( .A(n48), .Y(n301) );
  NOR2X1 U563 ( .A(n97), .B(n90), .Y(n88) );
  NOR2X1 U564 ( .A(n173), .B(n166), .Y(n164) );
  AOI21X1 U565 ( .A0(n143), .A1(n126), .B0(n127), .Y(n125) );
  OAI21XL U566 ( .A0(n128), .A1(n138), .B0(n129), .Y(n127) );
  NAND2X1 U567 ( .A(n329), .B(n291), .Y(n35) );
  CLKINVX1 U568 ( .A(n290), .Y(n329) );
  OAI21X1 U569 ( .A0(n70), .A1(n80), .B0(n71), .Y(n69) );
  OAI21X1 U570 ( .A0(n148), .A1(n156), .B0(n149), .Y(n143) );
  XNOR2X1 U571 ( .A(n286), .B(n34), .Y(SUM[4]) );
  NOR2X1 U572 ( .A(n284), .B(n279), .Y(n273) );
  NAND2X1 U573 ( .A(n317), .B(n197), .Y(n23) );
  OAI21XL U574 ( .A0(n257), .A1(n199), .B0(n200), .Y(n198) );
  CLKINVX1 U575 ( .A(n196), .Y(n317) );
  NAND2X1 U576 ( .A(n318), .B(n206), .Y(n24) );
  OAI21XL U577 ( .A0(n257), .A1(n208), .B0(n209), .Y(n207) );
  CLKINVX1 U578 ( .A(n203), .Y(n318) );
  NAND2X1 U579 ( .A(n319), .B(n217), .Y(n25) );
  CLKINVX1 U580 ( .A(n216), .Y(n319) );
  NAND2X1 U581 ( .A(n321), .B(n235), .Y(n27) );
  OAI21XL U582 ( .A0(n257), .A1(n237), .B0(n238), .Y(n236) );
  CLKINVX1 U583 ( .A(n234), .Y(n321) );
  XNOR2X1 U584 ( .A(n254), .B(n29), .Y(SUM[9]) );
  NAND2X1 U585 ( .A(n323), .B(n253), .Y(n29) );
  CLKINVX1 U586 ( .A(n252), .Y(n323) );
  XNOR2X1 U587 ( .A(n225), .B(n26), .Y(SUM[12]) );
  NAND2X1 U588 ( .A(n320), .B(n224), .Y(n26) );
  OAI21XL U589 ( .A0(n257), .A1(n226), .B0(n227), .Y(n225) );
  XNOR2X1 U590 ( .A(n243), .B(n28), .Y(SUM[10]) );
  NAND2X1 U591 ( .A(n322), .B(n242), .Y(n28) );
  OAI21XL U592 ( .A0(n257), .A1(n244), .B0(n245), .Y(n243) );
  INVXL U593 ( .A(n246), .Y(n244) );
  OAI21XL U594 ( .A0(n5), .A1(n44), .B0(n45), .Y(n43) );
  AOI21XL U595 ( .A0(n69), .A1(n46), .B0(n47), .Y(n45) );
  OAI21XL U596 ( .A0(n48), .A1(n60), .B0(n49), .Y(n47) );
  CLKINVX1 U597 ( .A(n59), .Y(n57) );
  CLKINVX1 U598 ( .A(n241), .Y(n322) );
  CLKINVX1 U599 ( .A(n223), .Y(n320) );
  CLKINVX1 U600 ( .A(n155), .Y(n312) );
  CLKINVX1 U601 ( .A(n117), .Y(n308) );
  NAND2X1 U602 ( .A(n330), .B(n294), .Y(n36) );
  CLKINVX1 U603 ( .A(n293), .Y(n330) );
  OAI21XL U604 ( .A0(n276), .A1(n268), .B0(n271), .Y(n267) );
  AOI21X1 U605 ( .A0(n229), .A1(n320), .B0(n222), .Y(n220) );
  CLKINVX1 U606 ( .A(n224), .Y(n222) );
  AOI21XL U607 ( .A0(n3), .A1(n308), .B0(n116), .Y(n114) );
  CLKINVX1 U608 ( .A(n118), .Y(n116) );
  AOI21XL U609 ( .A0(n161), .A1(n312), .B0(n154), .Y(n152) );
  CLKINVX1 U610 ( .A(n156), .Y(n154) );
  AOI21XL U611 ( .A0(n179), .A1(n314), .B0(n172), .Y(n170) );
  CLKINVX1 U612 ( .A(n174), .Y(n172) );
  AOI21XL U613 ( .A0(n3), .A1(n75), .B0(n76), .Y(n74) );
  OAI21XL U614 ( .A0(n5), .A1(n77), .B0(n80), .Y(n76) );
  AOI21X1 U615 ( .A0(n229), .A1(n201), .B0(n202), .Y(n200) );
  OAI21XL U616 ( .A0(n213), .A1(n203), .B0(n206), .Y(n202) );
  INVXL U617 ( .A(n211), .Y(n213) );
  AOI21XL U618 ( .A0(n3), .A1(n95), .B0(n96), .Y(n94) );
  OAI21XL U619 ( .A0(n107), .A1(n97), .B0(n100), .Y(n96) );
  INVXL U620 ( .A(n105), .Y(n107) );
  AOI21XL U621 ( .A0(n161), .A1(n133), .B0(n134), .Y(n132) );
  OAI21XL U622 ( .A0(n145), .A1(n135), .B0(n138), .Y(n134) );
  INVXL U623 ( .A(n143), .Y(n145) );
  XNOR2X1 U624 ( .A(n186), .B(n21), .Y(SUM[17]) );
  NAND2X1 U625 ( .A(n315), .B(n185), .Y(n21) );
  OAI21XL U626 ( .A0(n444), .A1(n187), .B0(n188), .Y(n186) );
  CLKINVX1 U627 ( .A(n184), .Y(n315) );
  NAND2X1 U628 ( .A(n305), .B(n91), .Y(n11) );
  OAI21XL U629 ( .A0(n444), .A1(n93), .B0(n94), .Y(n92) );
  CLKINVX1 U630 ( .A(n90), .Y(n305) );
  NAND2X1 U631 ( .A(n306), .B(n100), .Y(n12) );
  OAI21XL U632 ( .A0(n444), .A1(n102), .B0(n103), .Y(n101) );
  CLKINVX1 U633 ( .A(n97), .Y(n306) );
  XNOR2X1 U634 ( .A(n112), .B(n13), .Y(SUM[25]) );
  NAND2X1 U635 ( .A(n307), .B(n111), .Y(n13) );
  OAI21XL U636 ( .A0(n444), .A1(n113), .B0(n114), .Y(n112) );
  CLKINVX1 U637 ( .A(n110), .Y(n307) );
  NAND2X1 U638 ( .A(n309), .B(n129), .Y(n15) );
  OAI21XL U639 ( .A0(n444), .A1(n131), .B0(n132), .Y(n130) );
  CLKINVX1 U640 ( .A(n128), .Y(n309) );
  NAND2X1 U641 ( .A(n310), .B(n138), .Y(n16) );
  OAI21XL U642 ( .A0(n444), .A1(n140), .B0(n141), .Y(n139) );
  CLKINVX1 U643 ( .A(n135), .Y(n310) );
  NAND2X1 U644 ( .A(n311), .B(n149), .Y(n17) );
  CLKINVX1 U645 ( .A(n148), .Y(n311) );
  XNOR2X1 U646 ( .A(n168), .B(n19), .Y(SUM[19]) );
  NAND2X1 U647 ( .A(n313), .B(n167), .Y(n19) );
  OAI21XL U648 ( .A0(n444), .A1(n169), .B0(n170), .Y(n168) );
  CLKINVX1 U649 ( .A(n166), .Y(n313) );
  XNOR2X1 U650 ( .A(n119), .B(n14), .Y(SUM[24]) );
  NAND2X1 U651 ( .A(n308), .B(n118), .Y(n14) );
  OAI21XL U652 ( .A0(n444), .A1(n120), .B0(n121), .Y(n119) );
  INVX1 U653 ( .A(n4), .Y(n120) );
  XNOR2X1 U654 ( .A(n157), .B(n18), .Y(SUM[20]) );
  NAND2X1 U655 ( .A(n312), .B(n156), .Y(n18) );
  XNOR2X1 U656 ( .A(n175), .B(n20), .Y(SUM[18]) );
  NAND2X1 U657 ( .A(n314), .B(n174), .Y(n20) );
  OAI21XL U658 ( .A0(n444), .A1(n176), .B0(n177), .Y(n175) );
  NAND2X1 U659 ( .A(n304), .B(n80), .Y(n10) );
  CLKINVX1 U660 ( .A(n77), .Y(n304) );
  NAND2XL U661 ( .A(n57), .B(n60), .Y(n8) );
  OAI21XL U662 ( .A0(n444), .A1(n62), .B0(n63), .Y(n61) );
  NAND2X1 U663 ( .A(n303), .B(n71), .Y(n9) );
  CLKINVX1 U664 ( .A(n70), .Y(n303) );
  NOR2X1 U665 ( .A(n135), .B(n128), .Y(n126) );
  NOR2X1 U666 ( .A(n203), .B(n196), .Y(n194) );
  NOR2X1 U667 ( .A(n59), .B(n48), .Y(n46) );
  NAND2X1 U668 ( .A(n331), .B(n298), .Y(n37) );
  XOR2X1 U669 ( .A(n265), .B(n31), .Y(SUM[7]) );
  NAND2X1 U670 ( .A(n325), .B(n264), .Y(n31) );
  AOI21X1 U671 ( .A0(n286), .A1(n266), .B0(n267), .Y(n265) );
  CLKINVX1 U672 ( .A(n263), .Y(n325) );
  XOR2X1 U673 ( .A(n272), .B(n32), .Y(SUM[6]) );
  NAND2X1 U674 ( .A(n326), .B(n271), .Y(n32) );
  CLKINVX1 U675 ( .A(n268), .Y(n326) );
  XOR2X1 U676 ( .A(n444), .B(n22), .Y(SUM[16]) );
  NAND2X1 U677 ( .A(n316), .B(n188), .Y(n22) );
  XOR2X1 U678 ( .A(n257), .B(n30), .Y(SUM[8]) );
  CLKINVX1 U679 ( .A(n255), .Y(n324) );
  CLKINVX1 U680 ( .A(n284), .Y(n328) );
  XOR2X1 U681 ( .A(n281), .B(n33), .Y(SUM[5]) );
  NAND2X1 U682 ( .A(n327), .B(n280), .Y(n33) );
  AOI21X1 U683 ( .A0(n286), .A1(n328), .B0(n283), .Y(n281) );
  CLKINVX1 U684 ( .A(n279), .Y(n327) );
  NOR2BXL U685 ( .AN(n273), .B(n268), .Y(n266) );
  NAND2X1 U686 ( .A(B[10]), .B(A[10]), .Y(n242) );
  CLKINVX1 U687 ( .A(n38), .Y(SUM[0]) );
  NOR2XL U688 ( .A(B[0]), .B(A[0]), .Y(n299) );
endmodule


module ALU_DW_rightsh_5 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n3, n4, n5, n6, n7, n10, n11, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n109, n113, n114,
         n115, n116, n117, n118, n119, n120, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n199, n200, n201, n202, n205, n206, n211, n212, n213,
         n214, n219, n220, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414;

  NOR2BX4 U5 ( .AN(n34), .B(n394), .Y(B[30]) );
  NOR2BX4 U126 ( .AN(n105), .B(n414), .Y(n73) );
  MXI2X4 U256 ( .A(n57), .B(n55), .S0(n323), .Y(n382) );
  CLKINVX20 U257 ( .A(n397), .Y(n323) );
  OR2X4 U258 ( .A(SH[19]), .B(SH[9]), .Y(n214) );
  MX2X6 U259 ( .A(n83), .B(n87), .S0(n404), .Y(n51) );
  NOR2X6 U260 ( .A(n362), .B(n394), .Y(B[22]) );
  BUFX16 U261 ( .A(SH[4]), .Y(n407) );
  NOR2X2 U262 ( .A(n370), .B(n395), .Y(B[11]) );
  NAND2X6 U263 ( .A(n392), .B(n393), .Y(n199) );
  NOR2X6 U264 ( .A(n213), .B(n214), .Y(n393) );
  OR2X2 U265 ( .A(SH[13]), .B(SH[25]), .Y(n219) );
  BUFX20 U266 ( .A(n396), .Y(n397) );
  MX2X4 U267 ( .A(A[9]), .B(A[8]), .S0(n341), .Y(n340) );
  CLKMX2X6 U268 ( .A(n81), .B(n77), .S0(n337), .Y(n45) );
  CLKINVX20 U269 ( .A(n404), .Y(n337) );
  MX2X1 U270 ( .A(A[0]), .B(A[1]), .S0(n400), .Y(n164) );
  BUFX20 U271 ( .A(SH[2]), .Y(n401) );
  CLKMX2X6 U272 ( .A(n187), .B(n195), .S0(n405), .Y(n155) );
  MX2X6 U273 ( .A(n176), .B(n184), .S0(n406), .Y(n144) );
  CLKMX2X6 U274 ( .A(A[20]), .B(A[21]), .S0(n399), .Y(n184) );
  CLKMX2X6 U275 ( .A(n146), .B(n162), .S0(n410), .Y(n114) );
  NOR2BX4 U276 ( .AN(n122), .B(n412), .Y(n90) );
  CLKMX2X6 U277 ( .A(n68), .B(n325), .S0(n402), .Y(n36) );
  CLKMX2X6 U278 ( .A(n71), .B(n75), .S0(n404), .Y(n39) );
  AND2X8 U279 ( .A(n107), .B(n329), .Y(n75) );
  MX2X2 U280 ( .A(n171), .B(n179), .S0(n406), .Y(n139) );
  MX2X2 U281 ( .A(A[8]), .B(A[7]), .S0(n341), .Y(n171) );
  MX2X4 U282 ( .A(n36), .B(n38), .S0(n397), .Y(n4) );
  BUFX20 U283 ( .A(n411), .Y(n412) );
  BUFX20 U284 ( .A(SH[3]), .Y(n405) );
  NOR2X4 U285 ( .A(n201), .B(n202), .Y(n361) );
  NAND2X2 U286 ( .A(n385), .B(n386), .Y(n202) );
  AND3X4 U287 ( .A(n153), .B(n328), .C(n329), .Y(n89) );
  MX2X4 U288 ( .A(n85), .B(n89), .S0(n404), .Y(n53) );
  CLKMX2X2 U289 ( .A(n166), .B(n174), .S0(n406), .Y(n134) );
  NAND2X4 U290 ( .A(n344), .B(n345), .Y(n186) );
  CLKINVX3 U291 ( .A(n399), .Y(n349) );
  NOR2X4 U292 ( .A(n219), .B(n220), .Y(n390) );
  MXI2X2 U293 ( .A(n53), .B(n55), .S0(n397), .Y(n378) );
  NOR2X2 U294 ( .A(n324), .B(n395), .Y(B[12]) );
  NOR2X4 U295 ( .A(n363), .B(n394), .Y(B[23]) );
  MXI2X2 U296 ( .A(n61), .B(n63), .S0(n397), .Y(n365) );
  INVX12 U297 ( .A(n409), .Y(n328) );
  CLKINVX8 U298 ( .A(n399), .Y(n346) );
  BUFX16 U299 ( .A(n411), .Y(n413) );
  INVX12 U300 ( .A(n405), .Y(n342) );
  AND2X4 U301 ( .A(n353), .B(n354), .Y(n324) );
  MX2X6 U302 ( .A(n145), .B(n161), .S0(n410), .Y(n113) );
  NOR2X6 U303 ( .A(n364), .B(n395), .Y(B[18]) );
  CLKMX2X6 U304 ( .A(A[15]), .B(A[16]), .S0(n400), .Y(n179) );
  CLKMX2X6 U305 ( .A(n190), .B(n182), .S0(n342), .Y(n150) );
  NOR2X2 U306 ( .A(n367), .B(n394), .Y(B[28]) );
  BUFX20 U307 ( .A(n3), .Y(n395) );
  CLKAND2X12 U308 ( .A(n189), .B(n342), .Y(n157) );
  CLKMX2X6 U309 ( .A(A[25]), .B(A[26]), .S0(n399), .Y(n189) );
  MX2X6 U310 ( .A(n84), .B(n88), .S0(n404), .Y(n52) );
  CLKMX2X6 U311 ( .A(n137), .B(n153), .S0(n410), .Y(n105) );
  NOR2X6 U312 ( .A(n333), .B(n413), .Y(n79) );
  NAND2X6 U313 ( .A(A[24]), .B(n399), .Y(n356) );
  INVX3 U314 ( .A(n78), .Y(n327) );
  CLKINVX8 U315 ( .A(n82), .Y(n326) );
  NOR2X4 U316 ( .A(n377), .B(n395), .Y(B[8]) );
  MX2X6 U317 ( .A(A[11]), .B(A[12]), .S0(n400), .Y(n175) );
  CLKAND2X12 U318 ( .A(n130), .B(n329), .Y(n98) );
  CLKMX2X6 U319 ( .A(n181), .B(n173), .S0(n342), .Y(n141) );
  NOR2BX4 U320 ( .AN(n67), .B(n397), .Y(n35) );
  CLKMX2X6 U321 ( .A(n75), .B(n79), .S0(n404), .Y(n43) );
  NOR2X6 U322 ( .A(n384), .B(n394), .Y(B[24]) );
  INVX12 U323 ( .A(n400), .Y(n341) );
  NOR2BX4 U324 ( .AN(n104), .B(n414), .Y(n325) );
  MX2X6 U325 ( .A(n136), .B(n152), .S0(n408), .Y(n104) );
  NAND2X4 U326 ( .A(A[27]), .B(n357), .Y(n358) );
  CLKAND2X12 U327 ( .A(n154), .B(n328), .Y(n122) );
  CLKBUFX6 U328 ( .A(SH[5]), .Y(n411) );
  CLKAND2X8 U329 ( .A(n118), .B(n329), .Y(n86) );
  INVX16 U330 ( .A(n412), .Y(n329) );
  CLKAND2X8 U331 ( .A(n190), .B(n342), .Y(n158) );
  CLKMX2X6 U332 ( .A(n93), .B(n97), .S0(n403), .Y(n61) );
  NOR2X2 U333 ( .A(SH[28]), .B(SH[24]), .Y(n388) );
  CLKMX2X6 U334 ( .A(n91), .B(n95), .S0(n403), .Y(n59) );
  NOR2BX2 U335 ( .AN(n6), .B(n395), .Y(B[2]) );
  CLKAND2X12 U336 ( .A(n124), .B(n329), .Y(n92) );
  NAND2X2 U337 ( .A(n48), .B(n352), .Y(n353) );
  MXI2X6 U338 ( .A(n326), .B(n327), .S0(n337), .Y(n46) );
  CLKMX2X6 U339 ( .A(A[13]), .B(A[14]), .S0(n400), .Y(n177) );
  MX2X4 U340 ( .A(A[14]), .B(A[15]), .S0(n400), .Y(n178) );
  CLKAND2X8 U341 ( .A(n106), .B(n329), .Y(n74) );
  CLKMX2X3 U342 ( .A(n174), .B(n182), .S0(n406), .Y(n142) );
  NOR2X2 U343 ( .A(n369), .B(n394), .Y(B[27]) );
  CLKAND2X8 U344 ( .A(n109), .B(n329), .Y(n77) );
  CLKMX2X2 U345 ( .A(n167), .B(n175), .S0(n406), .Y(n135) );
  MXI2X4 U346 ( .A(n63), .B(n65), .S0(n397), .Y(n369) );
  CLKAND2X8 U347 ( .A(n126), .B(n329), .Y(n94) );
  MXI2X4 U348 ( .A(n52), .B(n50), .S0(n330), .Y(n376) );
  MXI2X4 U349 ( .A(n159), .B(n143), .S0(n328), .Y(n333) );
  CLKMX2X6 U350 ( .A(n94), .B(n98), .S0(n403), .Y(n62) );
  MXI2X4 U351 ( .A(n142), .B(n158), .S0(n410), .Y(n331) );
  CLKAND2X12 U352 ( .A(n113), .B(n329), .Y(n81) );
  NOR2X2 U353 ( .A(n366), .B(n394), .Y(B[26]) );
  MX2X2 U354 ( .A(A[6]), .B(A[7]), .S0(n400), .Y(n170) );
  CLKAND2X12 U355 ( .A(n128), .B(n329), .Y(n96) );
  MXI2X4 U356 ( .A(n54), .B(n52), .S0(n330), .Y(n371) );
  BUFX12 U357 ( .A(n396), .Y(n398) );
  CLKINVX12 U358 ( .A(n397), .Y(n330) );
  MXI2X4 U359 ( .A(n56), .B(n54), .S0(n330), .Y(n364) );
  NOR2X2 U360 ( .A(n332), .B(n413), .Y(n80) );
  MXI2X4 U361 ( .A(n144), .B(n160), .S0(n410), .Y(n332) );
  NAND2X6 U362 ( .A(n334), .B(n335), .Y(n60) );
  MX2X2 U363 ( .A(n42), .B(n44), .S0(n398), .Y(n10) );
  NOR2X4 U364 ( .A(n331), .B(n413), .Y(n78) );
  MXI2X2 U365 ( .A(n46), .B(n48), .S0(n398), .Y(n380) );
  CLKMX2X6 U366 ( .A(A[18]), .B(A[19]), .S0(n400), .Y(n182) );
  CLKMX2X3 U367 ( .A(A[2]), .B(A[3]), .S0(n400), .Y(n166) );
  CLKMX2X6 U368 ( .A(A[26]), .B(A[27]), .S0(n399), .Y(n190) );
  CLKMX2X3 U369 ( .A(n134), .B(n150), .S0(n408), .Y(n102) );
  MXI2X2 U370 ( .A(n56), .B(n58), .S0(n397), .Y(n383) );
  NAND2X4 U371 ( .A(A[28]), .B(n399), .Y(n359) );
  CLKAND2X8 U372 ( .A(n192), .B(n342), .Y(n160) );
  CLKMX2X6 U373 ( .A(n184), .B(n192), .S0(n405), .Y(n152) );
  MX2X2 U374 ( .A(n82), .B(n86), .S0(n404), .Y(n50) );
  NAND2X4 U375 ( .A(n92), .B(n337), .Y(n334) );
  NAND2X4 U376 ( .A(n96), .B(n403), .Y(n335) );
  BUFX20 U377 ( .A(n401), .Y(n403) );
  OR2X8 U378 ( .A(SH[30]), .B(n343), .Y(n205) );
  MX2X2 U379 ( .A(n80), .B(n84), .S0(n404), .Y(n48) );
  CLKMX2X6 U380 ( .A(A[24]), .B(A[25]), .S0(n399), .Y(n188) );
  MX2X4 U381 ( .A(A[12]), .B(A[13]), .S0(n400), .Y(n176) );
  MX2X2 U382 ( .A(A[1]), .B(A[2]), .S0(n400), .Y(n165) );
  NAND2X6 U383 ( .A(n358), .B(n359), .Y(n191) );
  MXI2X2 U384 ( .A(n51), .B(n53), .S0(n398), .Y(n379) );
  CLKMX2X6 U385 ( .A(A[28]), .B(A[29]), .S0(n399), .Y(n192) );
  NOR2X6 U386 ( .A(SH[29]), .B(SH[17]), .Y(n387) );
  NOR2BX4 U387 ( .AN(n10), .B(n395), .Y(B[6]) );
  MX2X6 U388 ( .A(A[9]), .B(A[10]), .S0(n400), .Y(n173) );
  MX2X4 U389 ( .A(n74), .B(n78), .S0(n404), .Y(n42) );
  MX2X4 U390 ( .A(A[30]), .B(A[31]), .S0(n399), .Y(n194) );
  BUFX4 U391 ( .A(SH[4]), .Y(n408) );
  CLKMX2X3 U392 ( .A(n169), .B(n177), .S0(n406), .Y(n137) );
  NOR2X2 U393 ( .A(n373), .B(n395), .Y(B[5]) );
  CLKMX2X2 U394 ( .A(A[5]), .B(A[6]), .S0(n400), .Y(n169) );
  CLKMX2X6 U395 ( .A(n141), .B(n157), .S0(n410), .Y(n109) );
  MXI2X4 U396 ( .A(n64), .B(n66), .S0(n397), .Y(n367) );
  OR2X2 U397 ( .A(SH[7]), .B(SH[21]), .Y(n220) );
  CLKMX2X6 U398 ( .A(n147), .B(n163), .S0(n410), .Y(n115) );
  NOR2BX4 U399 ( .AN(n122), .B(n412), .Y(n336) );
  NOR2BX4 U400 ( .AN(n97), .B(n403), .Y(n65) );
  MXI2X2 U401 ( .A(n65), .B(n67), .S0(n397), .Y(n368) );
  NOR2X1 U402 ( .A(SH[20]), .B(SH[18]), .Y(n389) );
  CLKMX2X6 U403 ( .A(n336), .B(n94), .S0(n403), .Y(n58) );
  NOR2X2 U404 ( .A(n381), .B(n395), .Y(B[13]) );
  NOR2X2 U405 ( .A(n365), .B(n394), .Y(B[25]) );
  NAND2X2 U406 ( .A(A[23]), .B(n399), .Y(n345) );
  INVX2 U407 ( .A(n399), .Y(n357) );
  MXI2X2 U408 ( .A(n40), .B(n42), .S0(n398), .Y(n374) );
  CLKMX2X6 U409 ( .A(n79), .B(n83), .S0(n404), .Y(n47) );
  OR2X2 U410 ( .A(SH[23]), .B(SH[27]), .Y(n213) );
  CLKMX2X6 U411 ( .A(n186), .B(n178), .S0(n342), .Y(n146) );
  NOR2X6 U412 ( .A(n375), .B(n395), .Y(B[9]) );
  MX2X4 U413 ( .A(A[19]), .B(A[20]), .S0(n399), .Y(n183) );
  MXI2X4 U414 ( .A(n140), .B(n156), .S0(n410), .Y(n339) );
  NOR2X8 U415 ( .A(n199), .B(n200), .Y(n360) );
  MX2X4 U416 ( .A(n325), .B(n76), .S0(n404), .Y(n40) );
  CLKMX2X6 U417 ( .A(n80), .B(n76), .S0(n337), .Y(n44) );
  CLKMX2X2 U418 ( .A(A[4]), .B(A[5]), .S0(n400), .Y(n168) );
  CLKMX2X6 U419 ( .A(A[30]), .B(A[31]), .S0(n399), .Y(n338) );
  CLKMX2X3 U420 ( .A(n38), .B(n40), .S0(n398), .Y(n6) );
  MXI2X4 U421 ( .A(n60), .B(n62), .S0(n397), .Y(n384) );
  CLKBUFX12 U422 ( .A(SH[3]), .Y(n406) );
  MX2X6 U423 ( .A(A[10]), .B(A[11]), .S0(n400), .Y(n174) );
  NAND2X4 U424 ( .A(A[23]), .B(n346), .Y(n355) );
  NOR2X2 U425 ( .A(n382), .B(n3), .Y(B[19]) );
  NOR2BX4 U426 ( .AN(n127), .B(n412), .Y(n95) );
  NOR2X4 U427 ( .A(n339), .B(n413), .Y(n76) );
  CLKBUFX20 U428 ( .A(n407), .Y(n409) );
  BUFX12 U429 ( .A(n413), .Y(n414) );
  NOR2X1 U430 ( .A(SH[6]), .B(SH[22]), .Y(n386) );
  MXI2X2 U431 ( .A(n41), .B(n43), .S0(n398), .Y(n373) );
  CLKMX2X4 U432 ( .A(n43), .B(n45), .S0(n398), .Y(n11) );
  MX2X4 U433 ( .A(A[16]), .B(A[17]), .S0(n400), .Y(n180) );
  MX2X6 U434 ( .A(n180), .B(n188), .S0(n406), .Y(n148) );
  NOR2BX4 U435 ( .AN(n162), .B(n409), .Y(n130) );
  CLKMX2X3 U436 ( .A(n135), .B(n151), .S0(n408), .Y(n103) );
  MX2X6 U437 ( .A(n183), .B(n191), .S0(n405), .Y(n151) );
  NOR2X2 U438 ( .A(SH[26]), .B(SH[8]), .Y(n391) );
  CLKMX2X6 U439 ( .A(n186), .B(n338), .S0(n405), .Y(n154) );
  NOR2BX2 U440 ( .AN(n35), .B(n394), .Y(B[31]) );
  NOR2BX4 U441 ( .AN(A[31]), .B(n399), .Y(n195) );
  OR2X4 U442 ( .A(SH[31]), .B(SH[15]), .Y(n212) );
  NAND2X6 U443 ( .A(n355), .B(n356), .Y(n187) );
  CLKMX2X3 U444 ( .A(n165), .B(n173), .S0(n406), .Y(n133) );
  CLKMX2X6 U445 ( .A(n70), .B(n74), .S0(n402), .Y(n38) );
  CLKMX2X2 U446 ( .A(n164), .B(n340), .S0(n406), .Y(n132) );
  CLKMX2X6 U447 ( .A(n86), .B(n90), .S0(n403), .Y(n54) );
  CLKMX2X6 U448 ( .A(n180), .B(n340), .S0(n342), .Y(n140) );
  NOR2BX4 U449 ( .AN(n96), .B(n403), .Y(n64) );
  OR2X2 U450 ( .A(SH[10]), .B(SH[12]), .Y(n211) );
  NAND2X4 U451 ( .A(A[21]), .B(n346), .Y(n347) );
  NOR2X2 U452 ( .A(n368), .B(n394), .Y(B[29]) );
  NOR2X2 U453 ( .A(n380), .B(n395), .Y(B[10]) );
  NAND2X2 U454 ( .A(A[22]), .B(n399), .Y(n348) );
  OR2X8 U455 ( .A(n205), .B(n206), .Y(n200) );
  NAND2X2 U456 ( .A(n389), .B(n388), .Y(n206) );
  NAND2X4 U457 ( .A(A[22]), .B(n346), .Y(n344) );
  NOR2BX2 U458 ( .AN(n66), .B(n397), .Y(n34) );
  MX2X2 U459 ( .A(n69), .B(n73), .S0(n402), .Y(n37) );
  NOR2BX4 U460 ( .AN(n158), .B(n409), .Y(n126) );
  CLKMX2X6 U461 ( .A(n181), .B(n189), .S0(n406), .Y(n149) );
  CLKMX2X6 U462 ( .A(n81), .B(n85), .S0(n404), .Y(n49) );
  NOR2BX4 U463 ( .AN(n7), .B(n395), .Y(B[3]) );
  CLKMX2X6 U464 ( .A(A[29]), .B(A[30]), .S0(n399), .Y(n193) );
  NOR2X2 U465 ( .A(n378), .B(n395), .Y(B[17]) );
  CLKMX2X6 U466 ( .A(n88), .B(n92), .S0(n403), .Y(n56) );
  NOR2BX4 U467 ( .AN(n156), .B(n409), .Y(n124) );
  CLKBUFX20 U468 ( .A(SH[0]), .Y(n399) );
  MXI2X4 U469 ( .A(n49), .B(n51), .S0(n398), .Y(n381) );
  NOR2BX4 U470 ( .AN(n195), .B(n405), .Y(n163) );
  NOR2BX4 U471 ( .AN(n99), .B(n403), .Y(n67) );
  BUFX20 U472 ( .A(n407), .Y(n410) );
  MX2X2 U473 ( .A(n179), .B(n187), .S0(n406), .Y(n147) );
  NOR2BX4 U474 ( .AN(n100), .B(n414), .Y(n68) );
  NOR2BX4 U475 ( .AN(n101), .B(n414), .Y(n69) );
  NOR2BX4 U476 ( .AN(n102), .B(n414), .Y(n70) );
  NAND2BX2 U477 ( .AN(SH[11]), .B(n387), .Y(n343) );
  NOR2BX4 U478 ( .AN(n157), .B(n409), .Y(n125) );
  MXI2X2 U479 ( .A(n57), .B(n59), .S0(n397), .Y(n372) );
  CLKMX2X6 U480 ( .A(n89), .B(n93), .S0(n403), .Y(n57) );
  MXI2X4 U481 ( .A(n59), .B(n61), .S0(n397), .Y(n363) );
  NAND2X2 U482 ( .A(A[18]), .B(n399), .Y(n351) );
  NAND2X4 U483 ( .A(n390), .B(n391), .Y(n201) );
  MXI2X1 U484 ( .A(n62), .B(n64), .S0(n397), .Y(n366) );
  NAND2X4 U485 ( .A(n347), .B(n348), .Y(n185) );
  CLKMX2X3 U486 ( .A(n170), .B(n178), .S0(n406), .Y(n138) );
  CLKMX2X6 U487 ( .A(n87), .B(n91), .S0(n403), .Y(n55) );
  NOR2BX4 U488 ( .AN(n98), .B(n403), .Y(n66) );
  MXI2X4 U489 ( .A(n58), .B(n60), .S0(n397), .Y(n362) );
  NOR2BX4 U490 ( .AN(n103), .B(n414), .Y(n71) );
  MX2X2 U491 ( .A(n95), .B(n99), .S0(n403), .Y(n63) );
  MX2X1 U492 ( .A(A[3]), .B(A[4]), .S0(n400), .Y(n167) );
  MXI2X4 U493 ( .A(n45), .B(n47), .S0(n398), .Y(n375) );
  NOR2BX4 U494 ( .AN(n125), .B(n412), .Y(n93) );
  NOR2BX4 U495 ( .AN(n151), .B(n409), .Y(n119) );
  NOR2BX4 U496 ( .AN(n116), .B(n413), .Y(n84) );
  NOR2BX4 U497 ( .AN(n148), .B(n410), .Y(n116) );
  CLKMX2X3 U498 ( .A(n132), .B(n148), .S0(n408), .Y(n100) );
  CLKMX2X3 U499 ( .A(n168), .B(n176), .S0(n406), .Y(n136) );
  MXI2X4 U500 ( .A(n44), .B(n46), .S0(n398), .Y(n377) );
  MX2X4 U501 ( .A(n73), .B(n77), .S0(n404), .Y(n41) );
  NOR2X2 U502 ( .A(n374), .B(n395), .Y(B[4]) );
  NOR2BX4 U503 ( .AN(n117), .B(n413), .Y(n85) );
  NOR2BX4 U504 ( .AN(n149), .B(n410), .Y(n117) );
  CLKBUFX2 U505 ( .A(SH[2]), .Y(n402) );
  NOR2BX4 U506 ( .AN(n131), .B(n412), .Y(n99) );
  NOR2BX4 U507 ( .AN(n163), .B(n409), .Y(n131) );
  NOR2BX4 U508 ( .AN(n129), .B(n412), .Y(n97) );
  NOR2BX4 U509 ( .AN(n161), .B(n409), .Y(n129) );
  CLKMX2X3 U510 ( .A(n139), .B(n155), .S0(n410), .Y(n107) );
  CLKMX2X3 U511 ( .A(n37), .B(n39), .S0(n397), .Y(n5) );
  NOR2BX4 U512 ( .AN(n160), .B(n409), .Y(n128) );
  MXI2X2 U513 ( .A(n47), .B(n49), .S0(n398), .Y(n370) );
  NOR2BX4 U514 ( .AN(n5), .B(n395), .Y(B[1]) );
  NOR2BX4 U515 ( .AN(n194), .B(n405), .Y(n162) );
  NOR2BX4 U516 ( .AN(n114), .B(n413), .Y(n82) );
  NOR2BX4 U517 ( .AN(n115), .B(n413), .Y(n83) );
  CLKMX2X2 U518 ( .A(n133), .B(n149), .S0(n408), .Y(n101) );
  BUFX20 U519 ( .A(SH[0]), .Y(n400) );
  NOR2BX4 U520 ( .AN(n123), .B(n412), .Y(n91) );
  NOR2BX4 U521 ( .AN(n155), .B(n409), .Y(n123) );
  NOR2BX4 U522 ( .AN(n119), .B(n412), .Y(n87) );
  NOR2BX4 U523 ( .AN(n4), .B(n395), .Y(B[0]) );
  NAND2X8 U524 ( .A(n360), .B(n361), .Y(n3) );
  CLKMX2X4 U525 ( .A(n138), .B(n154), .S0(n410), .Y(n106) );
  NOR2BX4 U526 ( .AN(n120), .B(n412), .Y(n88) );
  NOR2BX4 U527 ( .AN(n152), .B(n409), .Y(n120) );
  CLKMX2X4 U528 ( .A(n177), .B(n185), .S0(n406), .Y(n145) );
  NAND2X2 U529 ( .A(A[17]), .B(n349), .Y(n350) );
  NAND2X4 U530 ( .A(n350), .B(n351), .Y(n181) );
  NAND2X2 U531 ( .A(n50), .B(n398), .Y(n354) );
  INVXL U532 ( .A(n398), .Y(n352) );
  NOR2BX4 U533 ( .AN(n191), .B(n405), .Y(n159) );
  CLKMX2X2 U534 ( .A(n175), .B(n183), .S0(n406), .Y(n143) );
  CLKMX2X4 U535 ( .A(n185), .B(n193), .S0(n405), .Y(n153) );
  BUFX20 U536 ( .A(n401), .Y(n404) );
  NOR2BX4 U537 ( .AN(n193), .B(n405), .Y(n161) );
  NOR2X2 U538 ( .A(SH[16]), .B(SH[14]), .Y(n385) );
  NOR2BX4 U539 ( .AN(n188), .B(n405), .Y(n156) );
  NOR2BX4 U540 ( .AN(n11), .B(n394), .Y(B[7]) );
  NOR2X2 U541 ( .A(n383), .B(n394), .Y(B[20]) );
  BUFX20 U542 ( .A(n3), .Y(n394) );
  NOR2BX4 U543 ( .AN(n159), .B(n409), .Y(n127) );
  NOR2X4 U544 ( .A(n211), .B(n212), .Y(n392) );
  NOR2X1 U545 ( .A(n379), .B(n395), .Y(B[15]) );
  NOR2BX4 U546 ( .AN(n150), .B(n410), .Y(n118) );
  NOR2X2 U547 ( .A(n376), .B(n395), .Y(B[14]) );
  CLKMX2X3 U548 ( .A(n39), .B(n41), .S0(n398), .Y(n7) );
  CLKBUFX2 U549 ( .A(SH[1]), .Y(n396) );
  NOR2X2 U550 ( .A(n371), .B(n395), .Y(B[16]) );
  NOR2X2 U551 ( .A(n372), .B(n394), .Y(B[21]) );
endmodule


module ALU_DW_leftsh_5 ( A, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  wire   n3, n4, n5, n6, n10, n13, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n199, n200, n201, n202, n207, n208,
         n211, n212, n213, n214, n215, n216, n217, n218, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407;

  NOR2BX4 U35 ( .AN(n4), .B(n388), .Y(B[0]) );
  NOR2BX4 U67 ( .AN(n36), .B(n390), .Y(n4) );
  MX2X4 U69 ( .A(n98), .B(n94), .S0(n396), .Y(n66) );
  NOR2BX4 U98 ( .AN(n69), .B(n397), .Y(n37) );
  NOR2BX4 U99 ( .AN(n68), .B(n397), .Y(n36) );
  NOR2BX4 U105 ( .AN(n126), .B(n405), .Y(n94) );
  NOR2BX4 U131 ( .AN(n100), .B(n407), .Y(n68) );
  NOR2BX4 U160 ( .AN(n135), .B(n402), .Y(n103) );
  NOR2BX4 U162 ( .AN(n133), .B(n402), .Y(n101) );
  NOR2BX4 U163 ( .AN(n132), .B(n402), .Y(n100) );
  MX2X2 U255 ( .A(A[26]), .B(A[25]), .S0(n393), .Y(n190) );
  CLKAND2X12 U256 ( .A(n140), .B(n338), .Y(n108) );
  NOR2X4 U257 ( .A(n362), .B(n388), .Y(B[16]) );
  CLKAND2X12 U258 ( .A(n107), .B(n337), .Y(n75) );
  BUFX12 U259 ( .A(SH[4]), .Y(n401) );
  CLKAND2X12 U260 ( .A(n116), .B(n337), .Y(n84) );
  MX2X4 U261 ( .A(n184), .B(n176), .S0(n400), .Y(n152) );
  CLKINVX12 U262 ( .A(SH[13]), .Y(n331) );
  MX2X6 U263 ( .A(n178), .B(n170), .S0(n329), .Y(n146) );
  NAND2X4 U264 ( .A(n141), .B(n338), .Y(n322) );
  CLKMX2X6 U265 ( .A(n173), .B(n165), .S0(n328), .Y(n141) );
  INVX12 U266 ( .A(n402), .Y(n338) );
  AND2X8 U267 ( .A(n341), .B(n342), .Y(n321) );
  NAND2X8 U268 ( .A(n354), .B(n355), .Y(n3) );
  CLKMX2X6 U269 ( .A(n86), .B(n82), .S0(n398), .Y(n54) );
  MX2X4 U270 ( .A(A[13]), .B(A[12]), .S0(n392), .Y(n177) );
  CLKAND2X12 U271 ( .A(n114), .B(n335), .Y(n82) );
  NAND2X4 U272 ( .A(n73), .B(n397), .Y(n352) );
  MX2X4 U273 ( .A(n47), .B(n45), .S0(n390), .Y(n353) );
  MX2X4 U274 ( .A(n79), .B(n75), .S0(n397), .Y(n47) );
  NAND2X6 U275 ( .A(n324), .B(n325), .Y(n52) );
  MX2X6 U276 ( .A(A[9]), .B(A[8]), .S0(n392), .Y(n173) );
  CLKMX2X6 U277 ( .A(n176), .B(n168), .S0(n328), .Y(n144) );
  MXI2X4 U278 ( .A(n140), .B(n156), .S0(n338), .Y(n333) );
  BUFX12 U279 ( .A(SH[1]), .Y(n389) );
  CLKMX2X6 U280 ( .A(n76), .B(n72), .S0(n397), .Y(n44) );
  NOR2X4 U281 ( .A(n211), .B(n212), .Y(n385) );
  OR2X4 U282 ( .A(SH[31]), .B(SH[15]), .Y(n212) );
  NOR2X4 U283 ( .A(n373), .B(n387), .Y(B[19]) );
  CLKMX2X6 U284 ( .A(n85), .B(n81), .S0(n398), .Y(n53) );
  MX2X6 U285 ( .A(n80), .B(n76), .S0(n397), .Y(n48) );
  NOR2X6 U286 ( .A(n376), .B(n388), .Y(B[8]) );
  CLKMX2X6 U287 ( .A(n172), .B(n180), .S0(n326), .Y(n148) );
  BUFX6 U288 ( .A(n404), .Y(n407) );
  BUFX20 U289 ( .A(n334), .Y(n406) );
  BUFX20 U290 ( .A(SH[0]), .Y(n392) );
  NOR2X4 U291 ( .A(n201), .B(n202), .Y(n355) );
  INVX3 U292 ( .A(n329), .Y(n326) );
  NAND2X4 U293 ( .A(n346), .B(n347), .Y(n49) );
  INVX8 U294 ( .A(n399), .Y(n332) );
  INVX2 U295 ( .A(n392), .Y(n343) );
  NOR2X4 U296 ( .A(n372), .B(n388), .Y(B[23]) );
  CLKMX2X3 U297 ( .A(A[25]), .B(A[24]), .S0(n393), .Y(n189) );
  CLKMX2X3 U298 ( .A(A[27]), .B(A[26]), .S0(n393), .Y(n191) );
  MXI2X4 U299 ( .A(n63), .B(n61), .S0(n391), .Y(n358) );
  MX2X4 U300 ( .A(n95), .B(n91), .S0(n398), .Y(n63) );
  NAND2X4 U301 ( .A(n84), .B(n323), .Y(n324) );
  NAND2X2 U302 ( .A(n80), .B(n398), .Y(n325) );
  INVXL U303 ( .A(n398), .Y(n323) );
  CLKAND2X12 U304 ( .A(n112), .B(n335), .Y(n80) );
  BUFX20 U305 ( .A(n395), .Y(n398) );
  NOR2X2 U306 ( .A(SH[6]), .B(SH[22]), .Y(n380) );
  CLKMX2X6 U307 ( .A(n42), .B(n40), .S0(n390), .Y(n10) );
  CLKMX2X3 U308 ( .A(A[24]), .B(A[23]), .S0(n393), .Y(n188) );
  NAND2X6 U309 ( .A(n60), .B(n340), .Y(n341) );
  BUFX20 U310 ( .A(SH[0]), .Y(n393) );
  CLKAND2X12 U311 ( .A(n171), .B(n332), .Y(n139) );
  NAND2X6 U312 ( .A(n348), .B(n349), .Y(n42) );
  BUFX20 U313 ( .A(n389), .Y(n391) );
  BUFX20 U314 ( .A(n389), .Y(n390) );
  CLKINVX8 U315 ( .A(n391), .Y(n340) );
  CLKAND2X8 U316 ( .A(n164), .B(n327), .Y(n132) );
  CLKINVX20 U317 ( .A(n400), .Y(n327) );
  MX2X4 U318 ( .A(n148), .B(n132), .S0(n403), .Y(n116) );
  CLKMX2X6 U319 ( .A(n172), .B(n164), .S0(n400), .Y(n140) );
  BUFX20 U320 ( .A(SH[3]), .Y(n328) );
  BUFX20 U321 ( .A(SH[3]), .Y(n329) );
  BUFX8 U322 ( .A(SH[3]), .Y(n399) );
  NOR2X8 U323 ( .A(n215), .B(n216), .Y(n381) );
  OR2X4 U324 ( .A(SH[29]), .B(SH[17]), .Y(n215) );
  OR2X4 U325 ( .A(SH[28]), .B(SH[24]), .Y(n217) );
  NOR2X4 U326 ( .A(n330), .B(n405), .Y(n89) );
  MXI2X2 U327 ( .A(n153), .B(n137), .S0(n403), .Y(n330) );
  MX2X6 U328 ( .A(A[15]), .B(A[14]), .S0(n393), .Y(n179) );
  MX2X4 U329 ( .A(A[19]), .B(A[18]), .S0(n393), .Y(n183) );
  CLKAND2X8 U330 ( .A(n104), .B(n337), .Y(n72) );
  CLKAND2X12 U331 ( .A(n120), .B(n337), .Y(n88) );
  CLKMX2X3 U332 ( .A(n187), .B(n179), .S0(n328), .Y(n155) );
  NOR2X6 U333 ( .A(n217), .B(n218), .Y(n382) );
  MX2X4 U334 ( .A(A[14]), .B(A[13]), .S0(n392), .Y(n178) );
  NOR2X6 U335 ( .A(n339), .B(n387), .Y(B[7]) );
  MXI2X4 U336 ( .A(n49), .B(n47), .S0(n390), .Y(n371) );
  CLKAND2X8 U337 ( .A(n165), .B(n332), .Y(n133) );
  NOR2X4 U338 ( .A(SH[7]), .B(SH[21]), .Y(n384) );
  NOR2X2 U339 ( .A(n370), .B(n387), .Y(B[12]) );
  NOR2BX4 U340 ( .AN(n331), .B(SH[25]), .Y(n383) );
  MX2X4 U341 ( .A(A[5]), .B(A[4]), .S0(n392), .Y(n169) );
  CLKMX2X6 U342 ( .A(n89), .B(n85), .S0(n398), .Y(n57) );
  NOR2X1 U343 ( .A(n375), .B(n387), .Y(B[29]) );
  MXI2X4 U344 ( .A(n65), .B(n63), .S0(n391), .Y(n375) );
  CLKAND2X8 U345 ( .A(n166), .B(n332), .Y(n134) );
  CLKMX2X6 U346 ( .A(n166), .B(n174), .S0(n332), .Y(n142) );
  INVX20 U347 ( .A(n406), .Y(n335) );
  CLKAND2X12 U348 ( .A(n119), .B(n335), .Y(n87) );
  CLKBUFX12 U349 ( .A(n334), .Y(n405) );
  NOR2X4 U350 ( .A(n333), .B(n405), .Y(n92) );
  NOR2X2 U351 ( .A(n371), .B(n387), .Y(B[13]) );
  CLKAND2X12 U352 ( .A(n102), .B(n337), .Y(n70) );
  CLKMX2X6 U353 ( .A(n87), .B(n83), .S0(n398), .Y(n55) );
  CLKAND2X12 U354 ( .A(n101), .B(n337), .Y(n69) );
  CLKAND2X12 U355 ( .A(n103), .B(n337), .Y(n71) );
  CLKAND2X12 U356 ( .A(n106), .B(n337), .Y(n74) );
  INVX20 U357 ( .A(n407), .Y(n337) );
  BUFX8 U358 ( .A(SH[5]), .Y(n334) );
  CLKMX2X6 U359 ( .A(n152), .B(n136), .S0(n403), .Y(n120) );
  NOR2X6 U360 ( .A(n321), .B(n388), .Y(B[24]) );
  NAND2X6 U361 ( .A(n385), .B(n386), .Y(n199) );
  MXI2X4 U362 ( .A(n56), .B(n58), .S0(n340), .Y(n359) );
  CLKAND2X12 U363 ( .A(n122), .B(n337), .Y(n90) );
  CLKMX2X6 U364 ( .A(A[3]), .B(A[2]), .S0(n392), .Y(n167) );
  NOR2BX2 U365 ( .AN(n37), .B(n390), .Y(n5) );
  CLKBUFX6 U366 ( .A(SH[2]), .Y(n395) );
  MXI2X2 U367 ( .A(n46), .B(n44), .S0(n390), .Y(n367) );
  MX2X2 U368 ( .A(n188), .B(n180), .S0(n328), .Y(n156) );
  NOR2X6 U369 ( .A(n360), .B(n387), .Y(B[18]) );
  MX2X4 U370 ( .A(n96), .B(n92), .S0(n398), .Y(n64) );
  NAND2X4 U371 ( .A(A[2]), .B(n343), .Y(n344) );
  CLKMX2X6 U372 ( .A(A[12]), .B(A[11]), .S0(n392), .Y(n176) );
  MX2X4 U373 ( .A(n93), .B(n89), .S0(n398), .Y(n61) );
  CLKMX2X3 U374 ( .A(n186), .B(n178), .S0(n328), .Y(n154) );
  NOR2BX4 U375 ( .AN(n71), .B(n397), .Y(n39) );
  BUFX20 U376 ( .A(n393), .Y(n394) );
  OR2X1 U377 ( .A(SH[20]), .B(SH[18]), .Y(n218) );
  NOR2X6 U378 ( .A(n359), .B(n388), .Y(B[22]) );
  CLKMX2X3 U379 ( .A(n67), .B(n65), .S0(n391), .Y(n35) );
  CLKMX2X3 U380 ( .A(n195), .B(n187), .S0(n328), .Y(n163) );
  CLKMX2X6 U381 ( .A(A[31]), .B(A[30]), .S0(n394), .Y(n195) );
  NOR2X2 U382 ( .A(n363), .B(n388), .Y(B[21]) );
  CLKMX2X6 U383 ( .A(A[6]), .B(A[5]), .S0(n392), .Y(n170) );
  MX2X4 U384 ( .A(A[18]), .B(A[17]), .S0(n393), .Y(n182) );
  CLKMX2X6 U385 ( .A(A[1]), .B(A[0]), .S0(n392), .Y(n165) );
  MX2X2 U386 ( .A(n83), .B(n79), .S0(n398), .Y(n51) );
  NOR2BX4 U387 ( .AN(n70), .B(n397), .Y(n38) );
  NAND2X4 U388 ( .A(n70), .B(n397), .Y(n349) );
  MX2X4 U389 ( .A(n150), .B(n134), .S0(n403), .Y(n118) );
  CLKMX2X3 U390 ( .A(n192), .B(n184), .S0(n328), .Y(n160) );
  CLKMX2X3 U391 ( .A(n194), .B(n186), .S0(n328), .Y(n162) );
  CLKMX2X3 U392 ( .A(n193), .B(n185), .S0(n328), .Y(n161) );
  BUFX20 U393 ( .A(n3), .Y(n388) );
  OR2X1 U394 ( .A(SH[10]), .B(SH[12]), .Y(n211) );
  NOR2BX4 U395 ( .AN(n5), .B(n388), .Y(B[1]) );
  NOR2X2 U396 ( .A(n365), .B(n387), .Y(B[4]) );
  CLKBUFX2 U397 ( .A(SH[5]), .Y(n404) );
  NOR2BX4 U398 ( .AN(A[0]), .B(n392), .Y(n164) );
  CLKMX2X4 U399 ( .A(n38), .B(n36), .S0(n390), .Y(n6) );
  NOR2X2 U400 ( .A(SH[16]), .B(SH[14]), .Y(n379) );
  MX2X4 U401 ( .A(A[16]), .B(A[15]), .S0(n394), .Y(n180) );
  CLKMX2X6 U402 ( .A(A[10]), .B(A[9]), .S0(n392), .Y(n174) );
  NAND2X6 U403 ( .A(n381), .B(n382), .Y(n200) );
  CLKMX2X3 U404 ( .A(n161), .B(n145), .S0(n403), .Y(n129) );
  NOR2BX2 U405 ( .AN(n35), .B(n387), .Y(B[31]) );
  MX2X1 U406 ( .A(A[29]), .B(A[28]), .S0(n393), .Y(n193) );
  NOR2BX2 U407 ( .AN(n130), .B(n405), .Y(n98) );
  MX2X1 U408 ( .A(n162), .B(n146), .S0(n403), .Y(n130) );
  NOR2X8 U409 ( .A(n199), .B(n200), .Y(n354) );
  MX2X4 U410 ( .A(n154), .B(n138), .S0(n403), .Y(n122) );
  CLKMX2X2 U411 ( .A(n160), .B(n144), .S0(n403), .Y(n128) );
  CLKMX2X4 U412 ( .A(A[21]), .B(A[20]), .S0(n393), .Y(n185) );
  CLKAND2X12 U413 ( .A(n118), .B(n335), .Y(n86) );
  CLKMX2X6 U414 ( .A(n88), .B(n84), .S0(n398), .Y(n56) );
  MXI2X4 U415 ( .A(n43), .B(n41), .S0(n390), .Y(n339) );
  CLKMX2X6 U416 ( .A(n175), .B(n167), .S0(n329), .Y(n143) );
  MX2X6 U417 ( .A(A[11]), .B(A[10]), .S0(n392), .Y(n175) );
  MX2X1 U418 ( .A(A[28]), .B(A[27]), .S0(n393), .Y(n192) );
  NOR2BX4 U419 ( .AN(n144), .B(n402), .Y(n112) );
  MXI2X2 U420 ( .A(n50), .B(n48), .S0(n390), .Y(n366) );
  OR2X4 U421 ( .A(SH[11]), .B(SH[30]), .Y(n216) );
  NOR2X2 U422 ( .A(n358), .B(n388), .Y(B[27]) );
  CLKMX2X3 U423 ( .A(n149), .B(n133), .S0(n403), .Y(n117) );
  CLKMX2X6 U424 ( .A(n90), .B(n86), .S0(n398), .Y(n336) );
  NOR2BX4 U425 ( .AN(n167), .B(n400), .Y(n135) );
  CLKMX2X6 U426 ( .A(n72), .B(n68), .S0(n397), .Y(n40) );
  MXI2X4 U427 ( .A(n64), .B(n62), .S0(n391), .Y(n357) );
  CLKAND2X12 U428 ( .A(n110), .B(n337), .Y(n78) );
  NAND2X2 U429 ( .A(n383), .B(n384), .Y(n207) );
  CLKAND2X12 U430 ( .A(n105), .B(n337), .Y(n73) );
  MXI2X4 U431 ( .A(n50), .B(n52), .S0(n340), .Y(n362) );
  CLKMX2X6 U432 ( .A(n91), .B(n87), .S0(n398), .Y(n59) );
  OR2X4 U433 ( .A(SH[19]), .B(SH[9]), .Y(n214) );
  NAND2X4 U434 ( .A(n336), .B(n391), .Y(n342) );
  MX2X6 U435 ( .A(n177), .B(n169), .S0(n329), .Y(n145) );
  NOR2BX4 U436 ( .AN(n145), .B(n403), .Y(n113) );
  CLKMX2X3 U437 ( .A(n181), .B(n173), .S0(n329), .Y(n149) );
  CLKMX2X6 U438 ( .A(n182), .B(n174), .S0(n399), .Y(n150) );
  CLKMX2X6 U439 ( .A(A[22]), .B(A[21]), .S0(n393), .Y(n186) );
  CLKBUFX20 U440 ( .A(n401), .Y(n402) );
  CLKAND2X12 U441 ( .A(n137), .B(n338), .Y(n105) );
  CLKMX2X6 U442 ( .A(n90), .B(n86), .S0(n398), .Y(n58) );
  NAND2X4 U443 ( .A(n344), .B(n345), .Y(n166) );
  NOR2X2 U444 ( .A(n377), .B(n388), .Y(B[30]) );
  NOR2X1 U445 ( .A(n367), .B(n388), .Y(B[10]) );
  NOR2BX4 U446 ( .AN(n136), .B(n402), .Y(n104) );
  MXI2X4 U447 ( .A(n44), .B(n42), .S0(n390), .Y(n376) );
  CLKMX2X6 U448 ( .A(n45), .B(n43), .S0(n390), .Y(n13) );
  NOR2X8 U449 ( .A(n322), .B(n406), .Y(n77) );
  CLKMX2X2 U450 ( .A(n183), .B(n175), .S0(n400), .Y(n151) );
  CLKMX2X4 U451 ( .A(n157), .B(n141), .S0(n403), .Y(n125) );
  CLKMX2X6 U452 ( .A(A[7]), .B(A[6]), .S0(n392), .Y(n171) );
  CLKMX2X6 U453 ( .A(n75), .B(n71), .S0(n397), .Y(n43) );
  CLKMX2X6 U454 ( .A(n92), .B(n88), .S0(n398), .Y(n60) );
  CLKMX2X6 U455 ( .A(n73), .B(n69), .S0(n397), .Y(n41) );
  CLKMX2X4 U456 ( .A(A[30]), .B(A[29]), .S0(n394), .Y(n194) );
  NOR2BX4 U457 ( .AN(n147), .B(n403), .Y(n115) );
  NOR2X1 U458 ( .A(n364), .B(n387), .Y(B[20]) );
  MX2X4 U459 ( .A(n97), .B(n93), .S0(n396), .Y(n65) );
  NOR2BX4 U460 ( .AN(n129), .B(n405), .Y(n97) );
  NOR2BX4 U461 ( .AN(n139), .B(n402), .Y(n107) );
  NAND2X2 U462 ( .A(A[1]), .B(n392), .Y(n345) );
  MXI2X4 U463 ( .A(n54), .B(n52), .S0(n391), .Y(n360) );
  MXI2X2 U464 ( .A(n62), .B(n60), .S0(n391), .Y(n374) );
  CLKMX2X6 U465 ( .A(n179), .B(n171), .S0(n400), .Y(n147) );
  MXI2X4 U466 ( .A(n59), .B(n57), .S0(n391), .Y(n372) );
  CLKMX2X6 U467 ( .A(n78), .B(n74), .S0(n397), .Y(n46) );
  CLKMX2X2 U468 ( .A(n189), .B(n181), .S0(n328), .Y(n157) );
  MXI2X1 U469 ( .A(n48), .B(n46), .S0(n390), .Y(n370) );
  MXI2X2 U470 ( .A(n56), .B(n54), .S0(n391), .Y(n364) );
  NOR2BX2 U471 ( .AN(n128), .B(n405), .Y(n96) );
  MXI2X4 U472 ( .A(n55), .B(n53), .S0(n391), .Y(n373) );
  NAND2X6 U473 ( .A(n351), .B(n352), .Y(n45) );
  BUFX20 U474 ( .A(n401), .Y(n403) );
  MXI2X1 U475 ( .A(n41), .B(n39), .S0(n390), .Y(n356) );
  NOR2BX4 U476 ( .AN(n134), .B(n402), .Y(n102) );
  NOR2BX4 U477 ( .AN(n115), .B(n406), .Y(n83) );
  NAND2X2 U478 ( .A(n77), .B(n397), .Y(n347) );
  MXI2X4 U479 ( .A(n61), .B(n59), .S0(n391), .Y(n361) );
  INVX4 U480 ( .A(n397), .Y(n350) );
  BUFX20 U481 ( .A(n395), .Y(n397) );
  NOR2BX4 U482 ( .AN(n138), .B(n402), .Y(n106) );
  NOR2BX4 U483 ( .AN(n170), .B(n400), .Y(n138) );
  NOR2BX4 U484 ( .AN(n123), .B(n405), .Y(n91) );
  MX2X2 U485 ( .A(n155), .B(n139), .S0(n403), .Y(n123) );
  NOR2BX4 U486 ( .AN(n131), .B(n405), .Y(n99) );
  CLKMX2X2 U487 ( .A(n163), .B(n147), .S0(n403), .Y(n131) );
  MX2X2 U488 ( .A(A[17]), .B(A[16]), .S0(n393), .Y(n181) );
  NOR2BX4 U489 ( .AN(n117), .B(n406), .Y(n85) );
  NOR2BX4 U490 ( .AN(n143), .B(n402), .Y(n111) );
  CLKBUFX2 U491 ( .A(SH[2]), .Y(n396) );
  BUFX20 U492 ( .A(SH[3]), .Y(n400) );
  MXI2X2 U493 ( .A(n53), .B(n51), .S0(n391), .Y(n368) );
  NOR2BX4 U494 ( .AN(n169), .B(n328), .Y(n137) );
  NOR2BX4 U495 ( .AN(n168), .B(n329), .Y(n136) );
  CLKMX2X6 U496 ( .A(A[4]), .B(A[3]), .S0(n392), .Y(n168) );
  CLKMX2X6 U497 ( .A(n82), .B(n78), .S0(n398), .Y(n50) );
  MX2X4 U498 ( .A(A[20]), .B(A[19]), .S0(n393), .Y(n184) );
  CLKMX2X6 U499 ( .A(A[8]), .B(A[7]), .S0(n392), .Y(n172) );
  NAND2X4 U500 ( .A(n74), .B(n350), .Y(n348) );
  NOR2BX4 U501 ( .AN(n127), .B(n405), .Y(n95) );
  MX2X2 U502 ( .A(n159), .B(n143), .S0(n403), .Y(n127) );
  NAND2X6 U503 ( .A(n77), .B(n350), .Y(n351) );
  NOR2BX4 U504 ( .AN(n13), .B(n387), .Y(B[9]) );
  OR2X4 U505 ( .A(SH[27]), .B(SH[23]), .Y(n213) );
  CLKMX2X3 U506 ( .A(n151), .B(n135), .S0(n403), .Y(n119) );
  MXI2X1 U507 ( .A(n40), .B(n38), .S0(n390), .Y(n365) );
  NOR2BX4 U508 ( .AN(n125), .B(n405), .Y(n93) );
  OR2X2 U509 ( .A(n207), .B(n208), .Y(n201) );
  BUFX20 U510 ( .A(n3), .Y(n387) );
  CLKMX2X4 U511 ( .A(n158), .B(n142), .S0(n403), .Y(n126) );
  CLKMX2X4 U512 ( .A(n190), .B(n182), .S0(n329), .Y(n158) );
  NOR2X2 U513 ( .A(n374), .B(n387), .Y(B[26]) );
  CLKMX2X4 U514 ( .A(n94), .B(n90), .S0(n398), .Y(n62) );
  NOR2X4 U515 ( .A(n361), .B(n387), .Y(B[25]) );
  NAND2X4 U516 ( .A(n81), .B(n350), .Y(n346) );
  NOR2BX4 U517 ( .AN(n108), .B(n406), .Y(n76) );
  NOR2BX4 U518 ( .AN(n111), .B(n406), .Y(n79) );
  CLKMX2X4 U519 ( .A(A[23]), .B(A[22]), .S0(n393), .Y(n187) );
  CLKMX2X2 U520 ( .A(n185), .B(n177), .S0(n328), .Y(n153) );
  NOR2BX4 U521 ( .AN(n113), .B(n406), .Y(n81) );
  MXI2X2 U522 ( .A(n57), .B(n55), .S0(n391), .Y(n363) );
  MXI2X1 U523 ( .A(n51), .B(n49), .S0(n391), .Y(n369) );
  OR2X4 U524 ( .A(SH[26]), .B(SH[8]), .Y(n208) );
  NOR2X2 U525 ( .A(n368), .B(n388), .Y(B[17]) );
  NOR2BX2 U526 ( .AN(n6), .B(n388), .Y(B[2]) );
  MXI2X2 U527 ( .A(n66), .B(n64), .S0(n391), .Y(n377) );
  NOR2X2 U528 ( .A(n369), .B(n388), .Y(B[15]) );
  NOR2BX4 U529 ( .AN(n142), .B(n402), .Y(n110) );
  CLKMX2X4 U530 ( .A(n99), .B(n95), .S0(n396), .Y(n67) );
  NOR2X4 U531 ( .A(n213), .B(n214), .Y(n386) );
  NOR2BX4 U532 ( .AN(n146), .B(n403), .Y(n114) );
  NOR2X2 U533 ( .A(n357), .B(n388), .Y(B[28]) );
  NOR2BX4 U534 ( .AN(n353), .B(n388), .Y(B[11]) );
  NOR2BX4 U535 ( .AN(n10), .B(n388), .Y(B[6]) );
  NOR2X1 U536 ( .A(n356), .B(n388), .Y(B[5]) );
  NOR2X1 U537 ( .A(n366), .B(n388), .Y(B[14]) );
  NOR2X4 U538 ( .A(n378), .B(n388), .Y(B[3]) );
  MXI2X2 U539 ( .A(n39), .B(n37), .S0(n390), .Y(n378) );
  CLKMX2X2 U540 ( .A(n191), .B(n183), .S0(n329), .Y(n159) );
  NAND2X1 U541 ( .A(n379), .B(n380), .Y(n202) );
endmodule


module ALU ( clk, rst_n, ALUOp_regD, funct_regD, ALUinA, ALUinB, ALUout, 
        stall_muldiv );
  input [5:0] ALUOp_regD;
  input [5:0] funct_regD;
  input [31:0] ALUinA;
  input [31:0] ALUinB;
  output [31:0] ALUout;
  input clk, rst_n;
  output stall_muldiv;
  wire   \halfresult[32] , \stateplus2[0] , \stateplus4[1] , N953, N954, N955,
         N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966,
         N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977,
         N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988,
         N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999,
         N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009,
         N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1049, N1050, N1051,
         N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061,
         N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071,
         N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081,
         N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091,
         N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101,
         N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111,
         N1112, N1145, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1133,
         n1134, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1148, n1149, n1150, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1, n2, n3,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1132, n1135, n1136, n1137,
         n1147, n1151, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
  wire   [31:0] reg_lo;
  wire   [31:0] subaluinA;
  wire   [6:0] state;
  wire   [31:0] subaluinB;
  wire   [32:0] tempresult;
  wire   [31:0] hi_com;
  wire   [31:0] lo_com;
  wire   [31:0] ALUinA_com;
  wire   [31:0] ALUinB_com;
  wire   [6:0] stateplus1;
  wire   [6:0] state_next;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFFRX4 \reg_lo_reg[3]  ( .D(n1222), .CK(clk), .RN(n223), .Q(reg_lo[3]), .QN(
        n1127) );
  DFFRX4 \reg_lo_reg[2]  ( .D(n1193), .CK(clk), .RN(n223), .Q(reg_lo[2]), .QN(
        n1128) );
  DFFRX4 \reg_lo_reg[1]  ( .D(n1192), .CK(clk), .RN(n223), .Q(reg_lo[1]), .QN(
        n1129) );
  DFFRX4 \state_reg[0]  ( .D(state_next[0]), .CK(clk), .RN(n223), .Q(
        \stateplus2[0] ), .QN(n26) );
  DFFRX4 \state_reg[6]  ( .D(state_next[6]), .CK(clk), .RN(n227), .Q(state[6]), 
        .QN(n206) );
  DFFRX4 \state_reg[1]  ( .D(state_next[1]), .CK(clk), .RN(n227), .Q(
        \stateplus4[1] ), .QN(n19) );
  DFFRX4 \state_reg[5]  ( .D(state_next[5]), .CK(clk), .RN(n227), .Q(state[5]), 
        .QN(n25) );
  DFFRX4 \state_reg[4]  ( .D(state_next[4]), .CK(clk), .RN(n228), .Q(state[4]), 
        .QN(n204) );
  DFFRX4 \state_reg[3]  ( .D(state_next[3]), .CK(clk), .RN(n228), .Q(state[3]), 
        .QN(n203) );
  ALU_DW01_inc_0 add_1216 ( .A({state[6:2], \stateplus4[1] , \stateplus2[0] }), 
        .SUM(stateplus1) );
  ALU_DW01_add_6 r436 ( .A({n279, n278, n277, n92, n146, n275, n274, n273, 
        n272, n271, n83, n81, n268, n93, n266, n85, n264, n263, n262, n261, 
        n94, n78, n86, n257, n256, n255, n82, n88, n89, n251, n250, n249}), 
        .B({n248, ALUinB[30], n147, n247, n150, n246, n245, n244, ALUinB[23], 
        n131, ALUinB[21], n119, n133, ALUinB[18], n237, n222, n116, n213, n243, 
        n209, n215, n126, ALUinB[9], n218, n104, n136, n74, n406, n404, n96, 
        n398, n400}), .CI(1'b0), .SUM({N984, N983, N982, N981, N980, N979, 
        N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, 
        N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, 
        N954, N953}) );
  ALU_DW01_sub_4 r437 ( .A({n279, n278, n277, n276, n145, n275, n274, n273, 
        n272, n271, n83, n81, n268, n93, n266, n85, n264, n263, n262, n261, 
        n94, n78, n86, n257, n256, n80, n254, n88, n89, n251, n250, n249}), 
        .B({n248, ALUinB[30], n147, n247, n149, n246, n245, n244, ALUinB[23], 
        n131, ALUinB[21], n120, n134, ALUinB[18], n237, n221, n115, n211, n243, 
        n209, n216, n126, ALUinB[9], n218, n104, n137, n74, n406, n404, n402, 
        n398, n400}), .CI(1'b0), .DIFF({N1016, N1015, N1014, N1013, N1012, 
        N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, 
        N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, 
        N990, N989, N988, N987, N986, N985}) );
  ALU_DW01_sub_5 sub_0_root_add_0_root_add_1209_ni ( .A({n1573, n1573, n1573, 
        n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, 
        n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, 
        n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573, n1573}), .B({
        subaluinA[31:28], n64, subaluinA[26], n63, subaluinA[24:16], n69, 
        subaluinA[14:12], n66, subaluinA[10:0]}), .CI(1'b0), .DIFF(hi_com) );
  ALU_DW01_inc_2 add_1211 ( .A({1'b1, n1099, n1100, n1101, n1102, n1103, n1104, 
        n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
        n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
        n1125, n1126, n1127, n1128, n1129, n1130}), .SUM({\halfresult[32] , 
        lo_com}) );
  ALU_DW01_sub_7 sub_add_1212_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({n279, n278, n277, n92, n145, n275, n274, n273, n272, 
        n271, n83, n81, n268, n93, n266, n85, n264, n263, n262, n261, n94, n78, 
        n86, n257, n256, n80, n254, n88, n89, n251, n250, n249}), .CI(1'b0), 
        .DIFF(ALUinA_com) );
  ALU_DW01_sub_6 sub_add_1213_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({n248, ALUinB[30], n147, n247, n149, n246, n245, n244, 
        ALUinB[23], n131, ALUinB[21], n120, n134, ALUinB[18], n236, n222, n116, 
        n212, n243, n208, n216, n125, ALUinB[9], n218, n105, n137, n75, n406, 
        n404, n96, n398, n400}), .CI(1'b0), .DIFF({ALUinB_com[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  ALU_DW_cmp_1 r440 ( .A({n279, n278, n277, n92, n146, n275, n274, n273, n272, 
        n271, n83, n81, n268, n93, n266, n85, n264, n263, n262, n261, n94, 
        n259, n86, n257, n256, n80, n82, n253, n89, n251, n250, n249}), .B({
        n248, ALUinB[30], n148, n247, n149, n246, n245, n244, ALUinB[23], n131, 
        ALUinB[21], n120, n134, ALUinB[18], n236, n222, n115, n213, n243, n208, 
        n216, n125, ALUinB[9], n219, n105, n136, n74, n406, n404, n96, n398, 
        n400}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N1145)
         );
  ALU_DW01_add_8 add_1205 ( .A({1'b0, subaluinA[31:28], n20, subaluinA[26], 
        n63, subaluinA[24:16], n70, subaluinA[14:12], n67, subaluinA[10:0]}), 
        .B({1'b0, subaluinB}), .CI(1'b0), .SUM(tempresult) );
  ALU_DW_rightsh_5 r439 ( .A({n279, n278, n277, n276, n145, n275, n274, n273, 
        n272, n271, n270, n269, n268, n267, n266, n265, n264, n263, n262, n261, 
        n260, n259, n258, n257, n87, n80, n254, n253, n89, n251, n250, n249}), 
        .DATA_TC(1'b0), .SH({n248, ALUinB[30], n148, n247, n150, n246, n245, 
        n244, ALUinB[23], n131, ALUinB[21], n120, n134, ALUinB[18], n237, n222, 
        n115, n212, n243, n209, n215, n126, ALUinB[9], n219, n105, n136, n74, 
        n406, n404, n96, n398, n400}), .B({N1112, N1111, N1110, N1109, N1108, 
        N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, 
        N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, 
        N1087, N1086, N1085, N1084, N1083, N1082, N1081}) );
  ALU_DW_leftsh_5 sll_1444 ( .A({n279, n278, n277, n276, n145, n275, n274, 
        n273, n272, n271, n270, n269, n268, n267, n266, n265, n264, n263, n262, 
        n261, n260, n259, n258, n257, n87, n255, n254, n253, n252, n251, n250, 
        n249}), .SH({n248, ALUinB[30], n148, n247, n150, n246, n245, n244, 
        ALUinB[23], n131, ALUinB[21], n119, n134, ALUinB[18], n236, n221, n116, 
        n212, n243, n209, n216, n126, ALUinB[9], n219, n105, n136, n74, n406, 
        n404, n96, n398, n400}), .B({N1080, N1079, N1078, N1077, N1076, N1075, 
        N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, 
        N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, 
        N1054, N1053, N1052, N1051, N1050, N1049}) );
  DFFRX1 \operand_reg[31]  ( .D(n1098), .CK(clk), .RN(n223), .Q(n1066) );
  DFFRX1 \operand_reg[0]  ( .D(n1067), .CK(clk), .RN(n227), .Q(n1035) );
  DFFRX1 \operand_reg[29]  ( .D(n1096), .CK(clk), .RN(n223), .Q(n1064), .QN(
        n39) );
  DFFRX1 \operand_reg[28]  ( .D(n1095), .CK(clk), .RN(n223), .Q(n1063), .QN(
        n56) );
  DFFRX1 \operand_reg[30]  ( .D(n1097), .CK(clk), .RN(n223), .Q(n1065), .QN(
        n41) );
  DFFRX1 \operand_reg[3]  ( .D(n1070), .CK(clk), .RN(n229), .Q(n1038), .QN(n24) );
  DFFRX1 \operand_reg[1]  ( .D(n1068), .CK(clk), .RN(n227), .Q(n1036), .QN(n22) );
  DFFRX1 \operand_reg[2]  ( .D(n1069), .CK(clk), .RN(n229), .Q(n1037), .QN(n23) );
  DFFRX1 \operand_reg[18]  ( .D(n1085), .CK(clk), .RN(n230), .Q(n1053), .QN(
        n33) );
  DFFRX1 \operand_reg[23]  ( .D(n1090), .CK(clk), .RN(n229), .Q(n1058), .QN(
        n34) );
  DFFRX1 \operand_reg[15]  ( .D(n1082), .CK(clk), .RN(n230), .Q(n1050), .QN(
        n43) );
  DFFRX1 \operand_reg[7]  ( .D(n1074), .CK(clk), .RN(n229), .Q(n1042), .QN(n50) );
  DFFRX1 \operand_reg[20]  ( .D(n1087), .CK(clk), .RN(n230), .Q(n1055), .QN(
        n47) );
  DFFRX1 \operand_reg[12]  ( .D(n1079), .CK(clk), .RN(n228), .Q(n1047), .QN(
        n42) );
  DFFRX1 \operand_reg[27]  ( .D(n1094), .CK(clk), .RN(n223), .Q(n1062), .QN(
        n55) );
  DFFRX1 \operand_reg[24]  ( .D(n1091), .CK(clk), .RN(n229), .Q(n1059), .QN(
        n32) );
  DFFRX1 \operand_reg[19]  ( .D(n1086), .CK(clk), .RN(n230), .Q(n1054), .QN(
        n37) );
  DFFRX1 \operand_reg[22]  ( .D(n1089), .CK(clk), .RN(n229), .Q(n1057), .QN(
        n38) );
  DFFRX1 \operand_reg[21]  ( .D(n1088), .CK(clk), .RN(n229), .Q(n1056), .QN(
        n40) );
  DFFRX1 \operand_reg[13]  ( .D(n1080), .CK(clk), .RN(n228), .Q(n1048), .QN(
        n46) );
  DFFRX1 \operand_reg[5]  ( .D(n1072), .CK(clk), .RN(n229), .Q(n1040), .QN(n51) );
  DFFRX1 \operand_reg[6]  ( .D(n1073), .CK(clk), .RN(n229), .Q(n1041), .QN(n52) );
  DFFRX1 \operand_reg[14]  ( .D(n1081), .CK(clk), .RN(n230), .Q(n1049), .QN(
        n57) );
  DFFRX1 \operand_reg[25]  ( .D(n1092), .CK(clk), .RN(n229), .Q(n1060), .QN(
        n45) );
  DFFRX1 \operand_reg[10]  ( .D(n1077), .CK(clk), .RN(n228), .Q(n1045), .QN(
        n44) );
  DFFRX1 \operand_reg[17]  ( .D(n1084), .CK(clk), .RN(n230), .Q(n1052), .QN(
        n35) );
  DFFRX1 \operand_reg[26]  ( .D(n1093), .CK(clk), .RN(n223), .Q(n1061), .QN(
        n53) );
  DFFRX1 \operand_reg[16]  ( .D(n1083), .CK(clk), .RN(n230), .Q(n1051), .QN(
        n36) );
  DFFRX1 \operand_reg[11]  ( .D(n1078), .CK(clk), .RN(n228), .Q(n1046), .QN(
        n54) );
  DFFRX1 \operand_reg[9]  ( .D(n1076), .CK(clk), .RN(n228), .Q(n1044), .QN(n48) );
  DFFRX1 \operand_reg[8]  ( .D(n1075), .CK(clk), .RN(n229), .Q(n1043), .QN(n49) );
  DFFRX1 \reg_lo_reg[20]  ( .D(n1174), .CK(clk), .RN(n230), .Q(reg_lo[20]), 
        .QN(n1110) );
  DFFRX1 \reg_lo_reg[15]  ( .D(n1179), .CK(clk), .RN(n227), .Q(reg_lo[15]), 
        .QN(n1115) );
  DFFRX1 \reg_lo_reg[14]  ( .D(n1180), .CK(clk), .RN(n227), .Q(reg_lo[14]), 
        .QN(n1116) );
  DFFRX1 \reg_lo_reg[6]  ( .D(n1188), .CK(clk), .RN(n228), .Q(reg_lo[6]), .QN(
        n1124) );
  DFFRX1 \reg_lo_reg[19]  ( .D(n1175), .CK(clk), .RN(n227), .Q(reg_lo[19]), 
        .QN(n1111) );
  DFFRX1 \reg_lo_reg[18]  ( .D(n1176), .CK(clk), .RN(n227), .Q(reg_lo[18]), 
        .QN(n1112) );
  DFFRX1 \reg_lo_reg[11]  ( .D(n1183), .CK(clk), .RN(n226), .Q(reg_lo[11]), 
        .QN(n1119) );
  DFFRX1 \reg_lo_reg[17]  ( .D(n1177), .CK(clk), .RN(n227), .Q(reg_lo[17]), 
        .QN(n1113) );
  DFFRX1 \reg_lo_reg[26]  ( .D(n1168), .CK(clk), .RN(n231), .Q(reg_lo[26]), 
        .QN(n1104) );
  DFFRX1 \reg_lo_reg[28]  ( .D(n1166), .CK(clk), .RN(n231), .Q(reg_lo[28]), 
        .QN(n1102) );
  DFFRX1 \reg_lo_reg[13]  ( .D(n1181), .CK(clk), .RN(n227), .Q(reg_lo[13]), 
        .QN(n1117) );
  DFFRX1 \reg_lo_reg[29]  ( .D(n1165), .CK(clk), .RN(n231), .Q(reg_lo[29]), 
        .QN(n1101) );
  DFFRX1 \reg_lo_reg[24]  ( .D(n1170), .CK(clk), .RN(n230), .Q(reg_lo[24]), 
        .QN(n1106) );
  DFFRX1 \reg_lo_reg[16]  ( .D(n1178), .CK(clk), .RN(n227), .Q(reg_lo[16]), 
        .QN(n1114) );
  DFFRX1 \reg_lo_reg[23]  ( .D(n1171), .CK(clk), .RN(n230), .Q(reg_lo[23]), 
        .QN(n1107) );
  DFFRX1 \reg_lo_reg[10]  ( .D(n1184), .CK(clk), .RN(n226), .Q(reg_lo[10]), 
        .QN(n1120) );
  DFFRX1 \reg_lo_reg[30]  ( .D(n1164), .CK(clk), .RN(n231), .Q(reg_lo[30]), 
        .QN(n1100) );
  DFFRX1 \reg_lo_reg[25]  ( .D(n1169), .CK(clk), .RN(n231), .Q(reg_lo[25]), 
        .QN(n1105) );
  DFFRX1 \reg_lo_reg[8]  ( .D(n1186), .CK(clk), .RN(n226), .Q(reg_lo[8]), .QN(
        n1122) );
  DFFRX1 \reg_lo_reg[9]  ( .D(n1185), .CK(clk), .RN(n226), .Q(reg_lo[9]), .QN(
        n1121) );
  DFFRX1 \reg_lo_reg[5]  ( .D(n1189), .CK(clk), .RN(n228), .Q(reg_lo[5]), .QN(
        n1125) );
  DFFRX1 \reg_lo_reg[21]  ( .D(n1173), .CK(clk), .RN(n230), .Q(reg_lo[21]), 
        .QN(n1109) );
  DFFRX1 \reg_lo_reg[0]  ( .D(n1191), .CK(clk), .RN(n223), .Q(reg_lo[0]), .QN(
        n1130) );
  DFFRX2 \reg_lo_reg[4]  ( .D(n1190), .CK(clk), .RN(n228), .Q(reg_lo[4]), .QN(
        n1126) );
  DFFRX2 \reg_lo_reg[31]  ( .D(n1163), .CK(clk), .RN(n231), .Q(reg_lo[31]), 
        .QN(n1099) );
  DFFRX1 \reg_hi_reg[0]  ( .D(n1226), .CK(clk), .RN(n226), .Q(subaluinA[0]), 
        .QN(n1162) );
  DFFRX1 \reg_hi_reg[20]  ( .D(n1213), .CK(clk), .RN(n224), .Q(subaluinA[20]), 
        .QN(n1142) );
  DFFRX1 \reg_hi_reg[8]  ( .D(n1201), .CK(clk), .RN(n225), .Q(subaluinA[8]), 
        .QN(n1154) );
  DFFRX1 \reg_hi_reg[12]  ( .D(n1205), .CK(clk), .RN(n225), .Q(subaluinA[12]), 
        .QN(n1150) );
  DFFRX1 \reg_hi_reg[18]  ( .D(n1211), .CK(clk), .RN(n225), .Q(subaluinA[18]), 
        .QN(n1144) );
  DFFRX1 \reg_hi_reg[16]  ( .D(n1209), .CK(clk), .RN(n225), .Q(subaluinA[16]), 
        .QN(n1146) );
  DFFRX1 \reg_hi_reg[24]  ( .D(n1217), .CK(clk), .RN(n224), .Q(subaluinA[24]), 
        .QN(n1138) );
  DFFRX1 \reg_hi_reg[21]  ( .D(n1214), .CK(clk), .RN(n224), .Q(subaluinA[21]), 
        .QN(n1141) );
  DFFRX1 \reg_hi_reg[23]  ( .D(n1216), .CK(clk), .RN(n224), .Q(subaluinA[23]), 
        .QN(n1139) );
  DFFRX1 \reg_hi_reg[31]  ( .D(n1225), .CK(clk), .RN(n223), .Q(subaluinA[31]), 
        .QN(n1131) );
  DFFRX1 \reg_hi_reg[6]  ( .D(n1199), .CK(clk), .RN(n226), .Q(subaluinA[6]), 
        .QN(n1156) );
  DFFRX1 \reg_hi_reg[14]  ( .D(n1207), .CK(clk), .RN(n225), .Q(subaluinA[14]), 
        .QN(n1148) );
  DFFRX1 \reg_hi_reg[22]  ( .D(n1215), .CK(clk), .RN(n224), .Q(subaluinA[22]), 
        .QN(n1140) );
  DFFRX1 \reg_hi_reg[2]  ( .D(n1195), .CK(clk), .RN(n226), .Q(subaluinA[2]), 
        .QN(n1160) );
  DFFRX1 \reg_hi_reg[4]  ( .D(n1197), .CK(clk), .RN(n226), .Q(subaluinA[4]), 
        .QN(n1158) );
  DFFRX1 \reg_hi_reg[10]  ( .D(n1203), .CK(clk), .RN(n225), .Q(subaluinA[10]), 
        .QN(n1152) );
  DFFRX1 \reg_hi_reg[3]  ( .D(n1196), .CK(clk), .RN(n226), .Q(subaluinA[3]), 
        .QN(n1159) );
  DFFRX1 \reg_hi_reg[7]  ( .D(n1200), .CK(clk), .RN(n225), .Q(subaluinA[7]), 
        .QN(n1155) );
  DFFRX2 \reg_hi_reg[5]  ( .D(n1198), .CK(clk), .RN(n226), .Q(subaluinA[5]), 
        .QN(n1157) );
  DFFRX4 \reg_hi_reg[1]  ( .D(n1194), .CK(clk), .RN(n226), .Q(subaluinA[1]), 
        .QN(n1161) );
  DFFRX2 \reg_hi_reg[9]  ( .D(n1202), .CK(clk), .RN(n225), .Q(subaluinA[9]), 
        .QN(n1153) );
  DFFRX2 \reg_hi_reg[17]  ( .D(n1210), .CK(clk), .RN(n225), .Q(subaluinA[17]), 
        .QN(n1145) );
  DFFRX1 \operand_reg[4]  ( .D(n1071), .CK(clk), .RN(rst_n), .Q(n1039), .QN(
        n788) );
  DFFRX1 \reg_hi_reg[29]  ( .D(n1223), .CK(clk), .RN(n224), .Q(subaluinA[29]), 
        .QN(n1133) );
  DFFRX1 \reg_hi_reg[15]  ( .D(n1208), .CK(clk), .RN(n225), .Q(n652) );
  DFFRX1 \reg_hi_reg[25]  ( .D(n1218), .CK(clk), .RN(n224), .QN(n21) );
  DFFRX1 \reg_hi_reg[11]  ( .D(n1204), .CK(clk), .RN(n225), .Q(n628) );
  DFFRX1 \reg_hi_reg[30]  ( .D(n1224), .CK(clk), .RN(n224), .Q(subaluinA[30]), 
        .QN(n738) );
  DFFRX1 \reg_lo_reg[22]  ( .D(n1172), .CK(clk), .RN(n230), .Q(reg_lo[22]), 
        .QN(n1108) );
  DFFRX1 \reg_lo_reg[12]  ( .D(n1182), .CK(clk), .RN(n226), .Q(reg_lo[12]), 
        .QN(n1118) );
  DFFRX1 \reg_lo_reg[7]  ( .D(n1187), .CK(clk), .RN(n228), .Q(reg_lo[7]), .QN(
        n1123) );
  DFFRX1 \reg_lo_reg[27]  ( .D(n1167), .CK(clk), .RN(n231), .Q(reg_lo[27]), 
        .QN(n1103) );
  DFFRX1 \reg_hi_reg[26]  ( .D(n1219), .CK(clk), .RN(n224), .Q(subaluinA[26]), 
        .QN(n1481) );
  DFFRX1 \state_reg[2]  ( .D(state_next[2]), .CK(clk), .RN(rst_n), .Q(state[2]), .QN(n846) );
  DFFRX4 \reg_hi_reg[19]  ( .D(n1212), .CK(clk), .RN(n224), .Q(subaluinA[19]), 
        .QN(n1143) );
  DFFRX4 \reg_hi_reg[28]  ( .D(n1221), .CK(clk), .RN(n224), .Q(subaluinA[28]), 
        .QN(n1134) );
  DFFRX4 \reg_hi_reg[27]  ( .D(n1220), .CK(clk), .RN(n224), .Q(n20), .QN(n31)
         );
  DFFRX4 \reg_hi_reg[13]  ( .D(n1206), .CK(clk), .RN(n225), .Q(subaluinA[13]), 
        .QN(n1149) );
  CLKINVX20 U3 ( .A(n124), .Y(n126) );
  INVX20 U4 ( .A(n220), .Y(n221) );
  NAND2BX1 U5 ( .AN(n250), .B(n123), .Y(n987) );
  BUFX16 U6 ( .A(ALUinA[6]), .Y(n255) );
  BUFX16 U7 ( .A(ALUinA[20]), .Y(n269) );
  CLKAND2X3 U8 ( .A(N1001), .B(n1541), .Y(n1) );
  CLKAND2X3 U9 ( .A(N969), .B(n1542), .Y(n2) );
  AND2X4 U10 ( .A(N1065), .B(n152), .Y(n3) );
  NOR3X4 U11 ( .A(n1), .B(n2), .C(n3), .Y(n1355) );
  OA21X4 U12 ( .A0(n280), .A1(n1357), .B0(n1356), .Y(n12) );
  NAND2X8 U13 ( .A(n12), .B(n1355), .Y(ALUout[16]) );
  INVX16 U14 ( .A(n154), .Y(n1542) );
  AND4X1 U15 ( .A(n1353), .B(n1352), .C(n1351), .D(n1350), .Y(n1357) );
  AND3X8 U16 ( .A(n1564), .B(n397), .C(N1105), .Y(n1458) );
  INVX2 U17 ( .A(n207), .Y(n208) );
  NAND2X6 U18 ( .A(n100), .B(n1367), .Y(ALUout[17]) );
  NAND2X6 U19 ( .A(N980), .B(n1542), .Y(n13) );
  NAND2X6 U20 ( .A(N1012), .B(n1541), .Y(n14) );
  AND2X8 U21 ( .A(n13), .B(n14), .Y(n1500) );
  CLKINVX12 U22 ( .A(n1463), .Y(n1541) );
  INVX20 U23 ( .A(n405), .Y(n404) );
  INVX8 U24 ( .A(ALUinB[3]), .Y(n405) );
  AOI22X4 U25 ( .A0(N1059), .A1(n152), .B0(N1091), .B1(n1443), .Y(n189) );
  CLKINVX6 U26 ( .A(n243), .Y(n1315) );
  INVX20 U27 ( .A(ALUinB[0]), .Y(n401) );
  AOI222X4 U28 ( .A0(subaluinA[4]), .A1(n241), .B0(n1030), .B1(n242), .C0(
        reg_lo[4]), .C1(n389), .Y(n1132) );
  NAND2BX4 U29 ( .AN(n85), .B(n1347), .Y(n1349) );
  INVX8 U30 ( .A(n221), .Y(n1347) );
  INVX4 U31 ( .A(N1002), .Y(n1368) );
  BUFX20 U32 ( .A(ALUinA[21]), .Y(n83) );
  BUFX20 U33 ( .A(ALUinA[11]), .Y(n94) );
  INVX6 U34 ( .A(n408), .Y(n869) );
  INVX6 U35 ( .A(n549), .Y(n822) );
  BUFX12 U36 ( .A(ALUinA[28]), .Y(n276) );
  BUFX12 U37 ( .A(ALUinA[28]), .Y(n92) );
  BUFX20 U38 ( .A(ALUinA[5]), .Y(n254) );
  INVX20 U39 ( .A(n207), .Y(n209) );
  CLKAND2X2 U40 ( .A(n245), .B(n274), .Y(n1465) );
  INVX12 U41 ( .A(ALUinB[6]), .Y(n135) );
  INVX12 U42 ( .A(n135), .Y(n136) );
  CLKINVX16 U51 ( .A(n214), .Y(n216) );
  INVX16 U52 ( .A(ALUinB[11]), .Y(n214) );
  INVX3 U53 ( .A(n1480), .Y(n1478) );
  NAND2BX1 U54 ( .AN(n275), .B(n1477), .Y(n1480) );
  CLKINVX20 U55 ( .A(n235), .Y(n237) );
  INVX20 U56 ( .A(ALUinB[17]), .Y(n235) );
  INVX12 U57 ( .A(ALUinB[22]), .Y(n130) );
  NOR2X2 U58 ( .A(n130), .B(n77), .Y(n15) );
  INVX20 U59 ( .A(n130), .Y(n131) );
  BUFX8 U60 ( .A(n793), .Y(n321) );
  BUFX8 U61 ( .A(n793), .Y(n322) );
  INVX6 U62 ( .A(n794), .Y(n791) );
  BUFX16 U63 ( .A(n791), .Y(n320) );
  OR2X8 U64 ( .A(n1555), .B(n1553), .Y(n16) );
  INVX4 U65 ( .A(n504), .Y(n883) );
  BUFX3 U66 ( .A(n883), .Y(n375) );
  BUFX4 U67 ( .A(n883), .Y(n374) );
  CLKXOR2X2 U68 ( .A(n90), .B(n248), .Y(n1558) );
  NAND2BX1 U69 ( .AN(n251), .B(n127), .Y(n1000) );
  INVX20 U70 ( .A(n103), .Y(n104) );
  INVX3 U71 ( .A(n217), .Y(n219) );
  INVX20 U72 ( .A(n220), .Y(n222) );
  INVX3 U73 ( .A(n124), .Y(n125) );
  CLKINVX4 U74 ( .A(n249), .Y(n918) );
  NAND2BXL U75 ( .AN(n88), .B(n407), .Y(n1029) );
  INVX16 U76 ( .A(n210), .Y(n213) );
  AND2X1 U77 ( .A(n209), .B(n261), .Y(n159) );
  AOI2BB1X1 U78 ( .A0N(n392), .A1N(n159), .B0(n387), .Y(n1307) );
  OAI211X4 U79 ( .A0(n280), .A1(n1227), .B0(n1151), .C0(n1147), .Y(ALUout[4])
         );
  NOR3X6 U80 ( .A(n1261), .B(n30), .C(n1258), .Y(n1262) );
  CLKINVX8 U81 ( .A(N981), .Y(n71) );
  INVX12 U82 ( .A(n403), .Y(n402) );
  BUFX20 U83 ( .A(ALUinA[3]), .Y(n89) );
  INVX6 U84 ( .A(N1145), .Y(n929) );
  INVX4 U85 ( .A(n103), .Y(n105) );
  NAND2BXL U86 ( .AN(n86), .B(n1275), .Y(n1277) );
  BUFX8 U87 ( .A(ALUinA[11]), .Y(n260) );
  NAND2XL U88 ( .A(n967), .B(n91), .Y(n17) );
  NAND2X6 U89 ( .A(N1081), .B(n18), .Y(n927) );
  INVX3 U90 ( .A(n17), .Y(n18) );
  INVXL U91 ( .A(n976), .Y(n91) );
  INVX8 U92 ( .A(funct_regD[5]), .Y(n967) );
  NAND4X8 U93 ( .A(n1572), .B(n1571), .C(n1570), .D(n1569), .Y(ALUout[31]) );
  AOI22X1 U94 ( .A0(N1054), .A1(n170), .B0(N990), .B1(n239), .Y(n1237) );
  INVX12 U95 ( .A(ALUinB[2]), .Y(n403) );
  NAND3X8 U96 ( .A(n1490), .B(n1489), .C(n1488), .Y(ALUout[26]) );
  INVX8 U97 ( .A(ALUinB[1]), .Y(n399) );
  OAI211X1 U98 ( .A0(n1503), .A1(n1149), .B0(n1323), .C0(n1322), .Y(n1324) );
  AND2X8 U99 ( .A(n992), .B(n991), .Y(n170) );
  INVX8 U100 ( .A(n1137), .Y(n1443) );
  INVX1 U101 ( .A(n271), .Y(n77) );
  INVX3 U102 ( .A(n986), .Y(n988) );
  INVX8 U103 ( .A(funct_regD[1]), .Y(n976) );
  NAND2X6 U104 ( .A(n144), .B(n924), .Y(n951) );
  CLKMX2X4 U105 ( .A(n1512), .B(n381), .S0(n29), .Y(n1513) );
  CLKMX2X2 U106 ( .A(n1298), .B(n382), .S0(n1297), .Y(n1301) );
  INVX1 U107 ( .A(n1412), .Y(n1409) );
  AND2X8 U108 ( .A(n170), .B(n396), .Y(n152) );
  BUFX20 U109 ( .A(ALUinB[13]), .Y(n243) );
  BUFX4 U110 ( .A(n796), .Y(n323) );
  AOI222X1 U111 ( .A0(n932), .A1(n973), .B0(funct_regD[0]), .B1(n931), .C0(n79), .C1(n991), .Y(n950) );
  INVX3 U112 ( .A(n1383), .Y(n1381) );
  INVXL U113 ( .A(n379), .Y(n102) );
  NAND2X2 U114 ( .A(n380), .B(n1000), .Y(n1005) );
  NAND2BX1 U115 ( .AN(n983), .B(n991), .Y(n936) );
  NAND2X6 U116 ( .A(N1090), .B(n1443), .Y(n121) );
  AND2X6 U117 ( .A(n1417), .B(n1419), .Y(n154) );
  INVX3 U118 ( .A(n79), .Y(n957) );
  CLKINVX3 U119 ( .A(n152), .Y(n110) );
  CLKMX2X2 U120 ( .A(n382), .B(n1348), .S0(n1349), .Y(n1353) );
  NAND2X1 U121 ( .A(n158), .B(n240), .Y(n1362) );
  NAND4X4 U122 ( .A(n1498), .B(n1497), .C(n1496), .D(n1495), .Y(n1499) );
  NAND2X1 U123 ( .A(n380), .B(n1228), .Y(n1233) );
  CLKMX2X2 U124 ( .A(n381), .B(n1410), .S0(n1408), .Y(n1411) );
  INVX1 U125 ( .A(n1417), .Y(n1418) );
  OAI31X1 U126 ( .A0(n906), .A1(n905), .A2(n904), .B0(n903), .Y(n915) );
  INVX3 U127 ( .A(n1558), .Y(n903) );
  AOI222XL U128 ( .A0(n351), .A1(subaluinA[28]), .B0(tempresult[29]), .B1(n824), .C0(tempresult[30]), .C1(n354), .Y(n725) );
  CLKBUFX3 U129 ( .A(n328), .Y(n327) );
  INVX6 U130 ( .A(n316), .Y(n315) );
  INVX4 U131 ( .A(n358), .Y(n355) );
  AOI221X1 U132 ( .A0(n735), .A1(n943), .B0(hi_com[0]), .B1(n319), .C0(n557), 
        .Y(n562) );
  BUFX4 U133 ( .A(n824), .Y(n328) );
  BUFX20 U134 ( .A(ALUinA[8]), .Y(n257) );
  BUFX20 U135 ( .A(ALUinA[19]), .Y(n268) );
  INVX4 U136 ( .A(n212), .Y(n1328) );
  INVX4 U137 ( .A(ALUinB[18]), .Y(n1369) );
  NAND3X4 U138 ( .A(n176), .B(n1327), .C(n1326), .Y(ALUout[13]) );
  NAND3X4 U139 ( .A(n167), .B(n168), .C(n169), .Y(ALUout[15]) );
  AOI222XL U140 ( .A0(tempresult[28]), .A1(n353), .B0(tempresult[31]), .B1(
        n343), .C0(tempresult[27]), .C1(n824), .Y(n714) );
  AOI222XL U141 ( .A0(tempresult[23]), .A1(n353), .B0(tempresult[26]), .B1(
        n343), .C0(tempresult[22]), .C1(n824), .Y(n685) );
  OA22X2 U142 ( .A0(n312), .A1(n707), .B0(n314), .B1(n701), .Y(n704) );
  CLKBUFX2 U143 ( .A(rst_n), .Y(n232) );
  CLKBUFX2 U144 ( .A(rst_n), .Y(n233) );
  CLKBUFX2 U145 ( .A(rst_n), .Y(n234) );
  BUFX2 U146 ( .A(n369), .Y(n365) );
  INVX1 U147 ( .A(n873), .Y(n823) );
  INVX1 U148 ( .A(n746), .Y(n825) );
  BUFX2 U149 ( .A(n350), .Y(n349) );
  INVX1 U150 ( .A(n876), .Y(n368) );
  BUFX2 U151 ( .A(n368), .Y(n366) );
  BUFX2 U152 ( .A(n368), .Y(n367) );
  INVX1 U153 ( .A(n1560), .Y(n1510) );
  INVX3 U154 ( .A(n1505), .Y(n1551) );
  OR4X2 U155 ( .A(n929), .B(n947), .C(n939), .D(n981), .Y(n27) );
  AND4X6 U156 ( .A(n1302), .B(n1301), .C(n1300), .D(n1299), .Y(n28) );
  AND2X6 U157 ( .A(n1509), .B(n1508), .Y(n29) );
  INVX3 U158 ( .A(n938), .Y(n973) );
  OR2X8 U159 ( .A(n1260), .B(n1259), .Y(n30) );
  BUFX2 U160 ( .A(n172), .Y(n316) );
  INVX3 U161 ( .A(n870), .Y(n350) );
  INVX1 U162 ( .A(n734), .Y(n95) );
  OAI211X4 U163 ( .A0(n910), .A1(n421), .B0(n420), .C0(reg_lo[3]), .Y(n886) );
  CLKINVX1 U164 ( .A(n886), .Y(n892) );
  INVX4 U165 ( .A(n21), .Y(n63) );
  AOI222X4 U166 ( .A0(n824), .A1(n284), .B0(n286), .B1(n348), .C0(
        ALUinA_com[26]), .C1(n325), .Y(n434) );
  AND3X1 U167 ( .A(n204), .B(n846), .C(n203), .Y(n200) );
  NAND2X2 U168 ( .A(n196), .B(n410), .Y(n419) );
  AND4X4 U169 ( .A(n413), .B(n206), .C(n409), .D(n417), .Y(n196) );
  AOI222X1 U170 ( .A0(lo_com[22]), .A1(n371), .B0(n285), .B1(n361), .C0(n286), 
        .C1(n331), .Y(n802) );
  INVX12 U171 ( .A(n335), .Y(n331) );
  AOI222X1 U172 ( .A0(lo_com[16]), .A1(n372), .B0(n291), .B1(n362), .C0(n292), 
        .C1(n332), .Y(n462) );
  INVX8 U173 ( .A(n334), .Y(n332) );
  AOI222X4 U174 ( .A0(tempresult[12]), .A1(n354), .B0(tempresult[15]), .B1(
        n344), .C0(tempresult[11]), .C1(n824), .Y(n619) );
  INVX2 U175 ( .A(n358), .Y(n354) );
  OA22X1 U176 ( .A0(n313), .A1(n623), .B0(n315), .B1(n617), .Y(n620) );
  AO21X4 U177 ( .A0(n412), .A1(n907), .B0(n1129), .Y(n871) );
  OA22X1 U178 ( .A0(n1013), .A1(n908), .B0(n1129), .B1(n907), .Y(n914) );
  AOI222X4 U179 ( .A0(lo_com[30]), .A1(n372), .B0(tempresult[2]), .B1(n362), 
        .C0(tempresult[1]), .C1(n332), .Y(n507) );
  AOI222X1 U180 ( .A0(lo_com[27]), .A1(n371), .B0(reg_lo[31]), .B1(n361), .C0(
        n281), .C1(n331), .Y(n797) );
  INVX12 U181 ( .A(n364), .Y(n361) );
  AOI222X1 U182 ( .A0(lo_com[14]), .A1(n372), .B0(n293), .B1(n362), .C0(n294), 
        .C1(n333), .Y(n452) );
  INVX8 U183 ( .A(n334), .Y(n333) );
  NAND2X2 U184 ( .A(n206), .B(n1130), .Y(n796) );
  INVX8 U185 ( .A(tempresult[30]), .Y(n747) );
  NAND4X2 U186 ( .A(n721), .B(n720), .C(n719), .D(n718), .Y(n1220) );
  INVX8 U187 ( .A(tempresult[27]), .Y(n723) );
  AOI222X4 U188 ( .A0(tempresult[27]), .A1(n353), .B0(tempresult[30]), .B1(
        n343), .C0(tempresult[26]), .C1(n824), .Y(n709) );
  NAND4X2 U189 ( .A(n711), .B(n710), .C(n709), .D(n708), .Y(n1218) );
  OA22X1 U190 ( .A0(n312), .A1(n712), .B0(n314), .B1(n707), .Y(n710) );
  OA22X2 U191 ( .A0(n366), .A1(n717), .B0(n338), .B1(n712), .Y(n690) );
  INVX6 U192 ( .A(tempresult[25]), .Y(n712) );
  OA22X2 U193 ( .A0(n367), .A1(n728), .B0(n337), .B1(n723), .Y(n702) );
  NAND2X1 U194 ( .A(n859), .B(n753), .Y(n754) );
  INVX12 U195 ( .A(n172), .Y(n314) );
  INVX4 U196 ( .A(tempresult[23]), .Y(n701) );
  OA22X4 U197 ( .A0(n312), .A1(n659), .B0(n315), .B1(n653), .Y(n656) );
  INVX4 U198 ( .A(tempresult[15]), .Y(n653) );
  NAND2X4 U199 ( .A(n860), .B(n729), .Y(n737) );
  OA22X2 U200 ( .A0(n365), .A1(n707), .B0(n339), .B1(n701), .Y(n678) );
  AND2X8 U201 ( .A(n1061), .B(n323), .Y(subaluinB[26]) );
  NAND4X2 U202 ( .A(n621), .B(n620), .C(n619), .D(n618), .Y(n1203) );
  OA22X1 U203 ( .A0(n366), .A1(n647), .B0(n337), .B1(n641), .Y(n618) );
  NAND4X2 U204 ( .A(n651), .B(n650), .C(n649), .D(n648), .Y(n1208) );
  OA22X2 U205 ( .A0(n313), .A1(n653), .B0(n315), .B1(n647), .Y(n650) );
  OA22X2 U206 ( .A0(n366), .A1(n659), .B0(n337), .B1(n653), .Y(n630) );
  INVX8 U207 ( .A(tempresult[22]), .Y(n695) );
  AOI222X4 U208 ( .A0(tempresult[19]), .A1(n353), .B0(tempresult[22]), .B1(
        n343), .C0(tempresult[18]), .C1(n824), .Y(n661) );
  AOI222X4 U209 ( .A0(tempresult[22]), .A1(n353), .B0(tempresult[25]), .B1(
        n343), .C0(tempresult[21]), .C1(n824), .Y(n679) );
  NAND4X2 U210 ( .A(n675), .B(n674), .C(n673), .D(n672), .Y(n1212) );
  NAND4X2 U211 ( .A(n669), .B(n668), .C(n667), .D(n666), .Y(n1211) );
  OA22X2 U212 ( .A0(n366), .A1(n653), .B0(n337), .B1(n647), .Y(n624) );
  INVX6 U213 ( .A(tempresult[14]), .Y(n647) );
  OA21X4 U214 ( .A0(n1463), .A1(n1447), .B0(n1445), .Y(n58) );
  NAND2X6 U215 ( .A(n58), .B(n1446), .Y(ALUout[23]) );
  INVX3 U216 ( .A(N1008), .Y(n1447) );
  NAND2X4 U217 ( .A(N976), .B(n1542), .Y(n1445) );
  AOI222X4 U218 ( .A0(N1072), .A1(n152), .B0(n1444), .B1(n394), .C0(N1104), 
        .C1(n1443), .Y(n1446) );
  NAND2X6 U219 ( .A(N1005), .B(n1541), .Y(n1402) );
  CLKINVX12 U220 ( .A(ALUinB[16]), .Y(n220) );
  CLKAND2X2 U221 ( .A(n213), .B(n263), .Y(n161) );
  NAND2BXL U222 ( .AN(n261), .B(n1306), .Y(n1308) );
  NOR3X6 U223 ( .A(n1554), .B(n16), .C(n1556), .Y(n1557) );
  AND3X1 U224 ( .A(n248), .B(n279), .C(n242), .Y(n1555) );
  INVX12 U225 ( .A(n210), .Y(n211) );
  NOR4BBX1 U226 ( .AN(n166), .BN(n909), .C(n911), .D(n910), .Y(n913) );
  INVX3 U227 ( .A(n419), .Y(n910) );
  INVX1 U228 ( .A(n378), .Y(n166) );
  BUFX20 U229 ( .A(n912), .Y(n378) );
  INVX8 U230 ( .A(n865), .Y(n912) );
  BUFX16 U231 ( .A(ALUinA[7]), .Y(n87) );
  INVX2 U232 ( .A(n74), .Y(n117) );
  INVX2 U233 ( .A(n96), .Y(n127) );
  CLKINVX6 U234 ( .A(n210), .Y(n212) );
  BUFX20 U235 ( .A(ALUinB[27]), .Y(n150) );
  CLKINVX20 U236 ( .A(n401), .Y(n400) );
  BUFX20 U237 ( .A(ALUinA[7]), .Y(n256) );
  BUFX16 U238 ( .A(ALUinA[9]), .Y(n86) );
  BUFX16 U239 ( .A(ALUinA[10]), .Y(n78) );
  BUFX8 U240 ( .A(ALUinA[3]), .Y(n252) );
  BUFX16 U241 ( .A(ALUinB[20]), .Y(n120) );
  INVX8 U242 ( .A(n273), .Y(n1449) );
  NAND2X8 U243 ( .A(n151), .B(n1434), .Y(ALUout[22]) );
  AOI2BB1X1 U244 ( .A0N(n392), .A1N(n165), .B0(n387), .Y(n1229) );
  AND2X2 U245 ( .A(n74), .B(n254), .Y(n165) );
  INVX16 U246 ( .A(ALUinB[8]), .Y(n217) );
  NAND2BX4 U247 ( .AN(n257), .B(n217), .Y(n1265) );
  MX2X2 U248 ( .A(n387), .B(n384), .S0(n1561), .Y(n1556) );
  CLKINVX8 U249 ( .A(N1009), .Y(n1462) );
  AND2X8 U250 ( .A(ALUinB[23]), .B(n272), .Y(n180) );
  AND3X8 U251 ( .A(n111), .B(n112), .C(n113), .Y(n1390) );
  NAND3X4 U252 ( .A(n59), .B(n27), .C(n60), .Y(n61) );
  NAND2X6 U253 ( .A(n61), .B(n952), .Y(n965) );
  INVXL U254 ( .A(n202), .Y(n59) );
  INVX3 U255 ( .A(n953), .Y(n60) );
  CLKAND2X8 U256 ( .A(ALUOp_regD[1]), .B(n954), .Y(n202) );
  OAI211X4 U257 ( .A0(n950), .A1(n970), .B0(n949), .C0(n948), .Y(n953) );
  INVX2 U258 ( .A(n951), .Y(n952) );
  NAND3X2 U259 ( .A(n239), .B(n397), .C(N995), .Y(n187) );
  NAND2X6 U260 ( .A(n121), .B(n122), .Y(n1282) );
  NAND2X6 U261 ( .A(N1058), .B(n152), .Y(n122) );
  NAND3X8 U262 ( .A(n1518), .B(n1520), .C(n1519), .Y(ALUout[28]) );
  CLKINVX2 U263 ( .A(N974), .Y(n1420) );
  AND2X4 U264 ( .A(N1067), .B(n152), .Y(n106) );
  NAND4BX4 U265 ( .AN(n1248), .B(n62), .C(n1247), .D(n1246), .Y(n1249) );
  NAND2X2 U266 ( .A(N959), .B(n1354), .Y(n62) );
  NAND3BX2 U267 ( .AN(n836), .B(state[5]), .C(n200), .Y(n417) );
  NAND2X4 U268 ( .A(\stateplus4[1] ), .B(n201), .Y(n413) );
  NAND2BX4 U269 ( .AN(n904), .B(n419), .Y(n416) );
  AND2X4 U270 ( .A(n1059), .B(n323), .Y(subaluinB[24]) );
  INVX4 U271 ( .A(N1088), .Y(n1263) );
  INVX6 U272 ( .A(n31), .Y(n64) );
  CLKINVX6 U273 ( .A(n628), .Y(n65) );
  INVX4 U274 ( .A(n65), .Y(n66) );
  INVX8 U275 ( .A(n65), .Y(n67) );
  CLKINVX6 U276 ( .A(n652), .Y(n68) );
  INVX4 U277 ( .A(n68), .Y(n69) );
  INVX8 U278 ( .A(n68), .Y(n70) );
  AOI2BB1X4 U279 ( .A0N(n186), .A1N(n391), .B0(n387), .Y(n1524) );
  BUFX20 U280 ( .A(n1559), .Y(n391) );
  NAND2X6 U281 ( .A(N1080), .B(n152), .Y(n1571) );
  OAI2BB2X4 U282 ( .B0(n154), .B1(n71), .A0N(n1541), .A1N(N1013), .Y(n72) );
  CLKINVX8 U283 ( .A(n72), .Y(n1518) );
  OAI2BB1X4 U284 ( .A0N(n1541), .A1N(N1007), .B0(n1435), .Y(n73) );
  CLKINVX8 U285 ( .A(n73), .Y(n151) );
  INVX12 U286 ( .A(ALUinB[15]), .Y(n114) );
  CLKINVX12 U287 ( .A(ALUinB[19]), .Y(n132) );
  BUFX20 U288 ( .A(ALUinB[5]), .Y(n74) );
  NAND2X6 U289 ( .A(N977), .B(n1542), .Y(n1460) );
  OAI211X2 U290 ( .A0(n1527), .A1(n1560), .B0(n1526), .C0(n1525), .Y(n1528) );
  INVX3 U291 ( .A(n117), .Y(n75) );
  AND2X1 U292 ( .A(n247), .B(n276), .Y(n1511) );
  BUFX3 U293 ( .A(N985), .Y(n76) );
  CLKINVX12 U294 ( .A(ALUinB[14]), .Y(n210) );
  INVX12 U295 ( .A(n135), .Y(n137) );
  BUFX20 U296 ( .A(ALUinA[4]), .Y(n88) );
  BUFX20 U297 ( .A(ALUinA[18]), .Y(n267) );
  BUFX16 U298 ( .A(ALUinA[21]), .Y(n270) );
  NOR2X4 U299 ( .A(n401), .B(n918), .Y(n79) );
  BUFX20 U300 ( .A(ALUinA[6]), .Y(n80) );
  NAND4X8 U301 ( .A(n1516), .B(n1515), .C(n1514), .D(n1513), .Y(n1517) );
  AOI2BB1X1 U302 ( .A0N(n391), .A1N(n181), .B0(n388), .Y(n1494) );
  NAND3X2 U303 ( .A(n1237), .B(n1236), .C(n1235), .Y(n138) );
  AOI2BB1X2 U304 ( .A0N(n391), .A1N(n179), .B0(n388), .Y(n1371) );
  CLKAND2X3 U305 ( .A(ALUinB[18]), .B(n93), .Y(n179) );
  BUFX20 U306 ( .A(ALUinA[20]), .Y(n81) );
  NAND2X4 U307 ( .A(N1082), .B(n1564), .Y(n997) );
  NAND2X2 U308 ( .A(n380), .B(n1240), .Y(n1243) );
  AO22X2 U309 ( .A0(n988), .A1(n240), .B0(n380), .B1(n987), .Y(n989) );
  NAND2X2 U310 ( .A(n380), .B(n1296), .Y(n1302) );
  NAND2X2 U311 ( .A(n380), .B(n1265), .Y(n1268) );
  BUFX12 U312 ( .A(n1510), .Y(n380) );
  BUFX8 U313 ( .A(ALUinA[5]), .Y(n82) );
  NAND3BX2 U314 ( .AN(funct_regD[3]), .B(n934), .C(n933), .Y(n983) );
  INVX6 U315 ( .A(funct_regD[2]), .Y(n934) );
  NAND2BX1 U316 ( .AN(n80), .B(n135), .Y(n1240) );
  INVX20 U317 ( .A(n871), .Y(n824) );
  NAND2X4 U318 ( .A(N985), .B(n921), .Y(n944) );
  BUFX12 U319 ( .A(ALUinB[27]), .Y(n149) );
  NAND3X8 U320 ( .A(n1529), .B(n1531), .C(n1530), .Y(ALUout[29]) );
  INVX2 U321 ( .A(n398), .Y(n123) );
  NAND2XL U322 ( .A(n398), .B(n250), .Y(n986) );
  OR4XL U323 ( .A(n959), .B(n962), .C(n919), .D(ALUOp_regD[0]), .Y(n972) );
  INVX3 U324 ( .A(ALUOp_regD[1]), .Y(n959) );
  INVX3 U325 ( .A(ALUOp_regD[2]), .Y(n962) );
  INVX3 U326 ( .A(n919), .Y(n958) );
  NAND2X2 U327 ( .A(ALUOp_regD[3]), .B(n920), .Y(n919) );
  INVX3 U328 ( .A(ALUOp_regD[0]), .Y(n954) );
  NAND2X1 U329 ( .A(n379), .B(n1492), .Y(n1496) );
  INVX3 U330 ( .A(ALUinB[21]), .Y(n1407) );
  INVX1 U331 ( .A(n1028), .Y(n1030) );
  CLKMX2X2 U332 ( .A(n385), .B(n1452), .S0(n1455), .Y(n1453) );
  NAND2BX4 U333 ( .AN(n1451), .B(n1450), .Y(n1452) );
  CLKINVX12 U334 ( .A(n265), .Y(n84) );
  INVX20 U335 ( .A(n84), .Y(n85) );
  AOI222X1 U336 ( .A0(subaluinA[9]), .A1(n241), .B0(n174), .B1(n242), .C0(n302), .C1(n390), .Y(n1278) );
  NAND2X4 U337 ( .A(N1068), .B(n152), .Y(n111) );
  BUFX12 U338 ( .A(n1547), .Y(n90) );
  CLKINVX1 U339 ( .A(n279), .Y(n1547) );
  BUFX12 U340 ( .A(ALUinB[29]), .Y(n147) );
  BUFX16 U341 ( .A(ALUinA[18]), .Y(n93) );
  INVX4 U342 ( .A(ALUinB[30]), .Y(n1532) );
  AND2X1 U343 ( .A(ALUinB[30]), .B(n278), .Y(n192) );
  NAND2X6 U344 ( .A(N1010), .B(n1541), .Y(n139) );
  NAND3X4 U345 ( .A(n177), .B(n1305), .C(n1304), .Y(ALUout[11]) );
  INVX12 U346 ( .A(n749), .Y(n734) );
  NOR3X6 U347 ( .A(n106), .B(n107), .C(n108), .Y(n1379) );
  CLKINVX8 U348 ( .A(N1057), .Y(n109) );
  NAND2X6 U349 ( .A(N971), .B(n1542), .Y(n1378) );
  INVX20 U350 ( .A(n403), .Y(n96) );
  INVX20 U351 ( .A(n217), .Y(n218) );
  NAND3X6 U352 ( .A(n394), .B(N1016), .C(n239), .Y(n1569) );
  NAND2X1 U353 ( .A(n96), .B(n251), .Y(n1001) );
  CLKINVX6 U354 ( .A(n235), .Y(n236) );
  OAI211X2 U355 ( .A0(n1503), .A1(n1138), .B0(n1457), .C0(n1456), .Y(n1459) );
  CLKAND2X8 U356 ( .A(n221), .B(n85), .Y(n156) );
  NAND2X6 U357 ( .A(n128), .B(n1460), .Y(ALUout[24]) );
  OA21X2 U358 ( .A0(n926), .A1(n925), .B0(n395), .Y(n144) );
  OA22X2 U359 ( .A0(n1506), .A1(n957), .B0(n956), .B1(n1560), .Y(n964) );
  BUFX20 U360 ( .A(ALUinA[15]), .Y(n264) );
  CLKINVX8 U361 ( .A(n92), .Y(n1509) );
  NAND2X4 U362 ( .A(N970), .B(n1542), .Y(n97) );
  NAND2X1 U363 ( .A(n1365), .B(n394), .Y(n98) );
  NAND2X2 U364 ( .A(N1098), .B(n1443), .Y(n99) );
  AND3X2 U365 ( .A(n97), .B(n98), .C(n99), .Y(n1367) );
  OA21X4 U366 ( .A0(n1463), .A1(n1368), .B0(n1366), .Y(n100) );
  NAND4X1 U367 ( .A(n1364), .B(n1363), .C(n1362), .D(n1361), .Y(n1365) );
  BUFX16 U368 ( .A(ALUinB[20]), .Y(n119) );
  INVXL U369 ( .A(n406), .Y(n101) );
  OR2X2 U370 ( .A(n102), .B(n29), .Y(n1514) );
  NAND3BX1 U371 ( .AN(n1509), .B(n247), .C(n1534), .Y(n1515) );
  OAI221X1 U372 ( .A0(n1566), .A1(n979), .B0(n1419), .B1(n979), .C0(n978), .Y(
        n995) );
  NAND3X8 U373 ( .A(n1502), .B(n1501), .C(n1500), .Y(ALUout[27]) );
  AOI32X2 U374 ( .A0(N1060), .A1(n394), .A2(n170), .B0(N1092), .B1(n1443), .Y(
        n1304) );
  BUFX20 U375 ( .A(ALUinA[26]), .Y(n275) );
  BUFX16 U376 ( .A(ALUinB[29]), .Y(n148) );
  INVX1 U377 ( .A(ALUinB[23]), .Y(n1436) );
  NAND4X4 U378 ( .A(n1403), .B(n1404), .C(n1402), .D(n1405), .Y(ALUout[20]) );
  CLKINVX12 U379 ( .A(ALUinB[7]), .Y(n103) );
  CLKAND2X8 U380 ( .A(N1099), .B(n1443), .Y(n108) );
  INVX1 U381 ( .A(n1029), .Y(n1032) );
  NAND2BX1 U382 ( .AN(n264), .B(n114), .Y(n1340) );
  AOI211X4 U383 ( .A0(N953), .A1(n969), .B0(n946), .C0(n945), .Y(n949) );
  NAND2X4 U384 ( .A(n918), .B(n118), .Y(n955) );
  NAND2X1 U385 ( .A(n379), .B(n1480), .Y(n1485) );
  NAND2X2 U386 ( .A(n104), .B(n256), .Y(n1256) );
  AOI222X4 U387 ( .A0(subaluinA[14]), .A1(n241), .B0(n161), .B1(n242), .C0(
        n297), .C1(n390), .Y(n1332) );
  NAND4X4 U388 ( .A(n1335), .B(n1334), .C(n1333), .D(n1332), .Y(n1336) );
  INVX4 U389 ( .A(N1004), .Y(n1391) );
  NAND2X4 U390 ( .A(N972), .B(n1542), .Y(n1389) );
  INVX4 U391 ( .A(n120), .Y(n1392) );
  NAND3X6 U392 ( .A(n1545), .B(n1544), .C(n1543), .Y(ALUout[30]) );
  NAND3BX4 U393 ( .AN(n995), .B(n994), .C(n993), .Y(n996) );
  AOI2BB1X4 U394 ( .A0N(n392), .A1N(n1253), .B0(n387), .Y(n1254) );
  AND2X2 U395 ( .A(n1377), .B(n394), .Y(n107) );
  NAND4X1 U396 ( .A(n1376), .B(n1375), .C(n1374), .D(n1373), .Y(n1377) );
  NAND2X2 U397 ( .A(N1077), .B(n152), .Y(n1520) );
  AOI32X2 U398 ( .A0(N1062), .A1(n394), .A2(n170), .B0(N1094), .B1(n1443), .Y(
        n1326) );
  INVX6 U399 ( .A(funct_regD[0]), .Y(n975) );
  NAND2X2 U400 ( .A(n985), .B(n984), .Y(n1503) );
  INVX4 U401 ( .A(n942), .Y(n985) );
  BUFX20 U402 ( .A(n1552), .Y(n241) );
  INVX8 U403 ( .A(n1503), .Y(n1552) );
  NAND2X8 U404 ( .A(n975), .B(n976), .Y(n941) );
  INVX16 U405 ( .A(n132), .Y(n133) );
  AOI211X2 U406 ( .A0(n379), .A1(n1321), .B0(n1320), .C0(n1319), .Y(n1322) );
  CLKMX2X3 U407 ( .A(n384), .B(n1318), .S0(n1321), .Y(n1319) );
  AOI2BB1X2 U408 ( .A0N(n1316), .A1N(n1315), .B0(n391), .Y(n1317) );
  INVX1 U409 ( .A(n262), .Y(n1316) );
  OAI2BB2X4 U410 ( .B0(n109), .B1(n110), .A0N(n1443), .A1N(N1089), .Y(n1270)
         );
  INVX3 U411 ( .A(n247), .Y(n1508) );
  NAND2BX1 U412 ( .AN(n274), .B(n1464), .Y(n1466) );
  INVX4 U413 ( .A(n245), .Y(n1464) );
  NAND4X4 U414 ( .A(n1387), .B(n1386), .C(n1385), .D(n1384), .Y(n1388) );
  AOI2BB1X1 U415 ( .A0N(n391), .A1N(n182), .B0(n388), .Y(n1382) );
  NAND2X8 U416 ( .A(n1475), .B(n1474), .Y(ALUout[25]) );
  NAND2X2 U417 ( .A(n1388), .B(n394), .Y(n112) );
  NAND2X2 U418 ( .A(N1100), .B(n1443), .Y(n113) );
  BUFX20 U419 ( .A(n393), .Y(n394) );
  OAI211X2 U420 ( .A0(n1463), .A1(n1391), .B0(n1390), .C0(n1389), .Y(
        ALUout[19]) );
  NAND2XL U421 ( .A(n379), .B(n1466), .Y(n1472) );
  AOI2BB2X4 U422 ( .B0(n1401), .B1(n394), .A0N(n280), .A1N(n1400), .Y(n1405)
         );
  AND2X8 U423 ( .A(n911), .B(n729), .Y(n172) );
  INVX12 U424 ( .A(tempresult[31]), .Y(n729) );
  INVX6 U425 ( .A(n150), .Y(n1491) );
  NAND2BX4 U426 ( .AN(n1567), .B(N984), .Y(n1570) );
  INVX12 U427 ( .A(n114), .Y(n115) );
  CLKINVX8 U428 ( .A(n114), .Y(n116) );
  INVXL U429 ( .A(n400), .Y(n118) );
  NAND2BX4 U430 ( .AN(n93), .B(n1369), .Y(n1372) );
  AOI2BB1X2 U431 ( .A0N(n1449), .A1N(n1448), .B0(n391), .Y(n1451) );
  OR2X4 U432 ( .A(n1273), .B(n1272), .Y(n143) );
  AND2X4 U433 ( .A(n149), .B(n146), .Y(n181) );
  CLKAND2X12 U434 ( .A(n971), .B(n984), .Y(n178) );
  INVX6 U435 ( .A(n982), .Y(n984) );
  OAI2BB1X1 U436 ( .A0N(n973), .A1N(n178), .B0(n972), .Y(n974) );
  INVX16 U437 ( .A(n132), .Y(n134) );
  MX2X1 U438 ( .A(n381), .B(n1524), .S0(n1523), .Y(n1525) );
  NAND2X1 U439 ( .A(n1522), .B(n1521), .Y(n1523) );
  CLKAND2X8 U440 ( .A(n120), .B(n81), .Y(n185) );
  NAND2X1 U441 ( .A(N957), .B(n1354), .Y(n1033) );
  NAND2X6 U442 ( .A(N975), .B(n1542), .Y(n1434) );
  AND2X1 U443 ( .A(n137), .B(n80), .Y(n184) );
  NAND2X1 U444 ( .A(n1449), .B(n1448), .Y(n1455) );
  NAND2X4 U445 ( .A(N1083), .B(n1564), .Y(n1012) );
  MX2X2 U446 ( .A(n381), .B(n977), .S0(n987), .Y(n978) );
  AOI2BB1X2 U447 ( .A0N(n391), .A1N(n158), .B0(n388), .Y(n1359) );
  AND2X1 U448 ( .A(n237), .B(n266), .Y(n158) );
  INVXL U449 ( .A(n1523), .Y(n1527) );
  CLKINVX6 U450 ( .A(n1546), .Y(n1561) );
  NAND2X6 U451 ( .A(n90), .B(n859), .Y(n1546) );
  MX2X1 U452 ( .A(n382), .B(n1254), .S0(n1252), .Y(n1255) );
  NAND2BX1 U453 ( .AN(n256), .B(n103), .Y(n1252) );
  AOI22X2 U454 ( .A0(N1063), .A1(n152), .B0(N1095), .B1(n1443), .Y(n164) );
  NAND2X2 U455 ( .A(N1076), .B(n152), .Y(n1501) );
  INVX12 U456 ( .A(ALUinB[12]), .Y(n207) );
  INVX6 U457 ( .A(n246), .Y(n1477) );
  CLKINVX12 U458 ( .A(ALUinB[10]), .Y(n124) );
  NAND4X2 U459 ( .A(n1432), .B(n1431), .C(n1430), .D(n1429), .Y(n1433) );
  MX2X1 U460 ( .A(n1427), .B(n381), .S0(n1426), .Y(n1432) );
  INVX3 U461 ( .A(n131), .Y(n1425) );
  NAND2BX4 U462 ( .AN(n268), .B(n132), .Y(n1383) );
  AND4X2 U463 ( .A(n1269), .B(n1268), .C(n1267), .D(n1266), .Y(n1274) );
  CLKMX2X2 U464 ( .A(n382), .B(n1264), .S0(n1265), .Y(n1269) );
  AOI222XL U465 ( .A0(subaluinA[8]), .A1(n241), .B0(n157), .B1(n242), .C0(n303), .C1(n390), .Y(n1266) );
  AND2X2 U466 ( .A(n219), .B(n257), .Y(n157) );
  OAI221X1 U467 ( .A0(n1413), .A1(n1560), .B0(n1506), .B1(n1412), .C0(n1411), 
        .Y(n1414) );
  INVX4 U468 ( .A(n148), .Y(n1521) );
  INVX8 U469 ( .A(n244), .Y(n1448) );
  OAI2BB2X4 U470 ( .B0(n280), .B1(n1012), .A0N(n1011), .A1N(n397), .Y(
        ALUout[2]) );
  NAND2X2 U471 ( .A(N1079), .B(n152), .Y(n1544) );
  BUFX20 U472 ( .A(n1559), .Y(n392) );
  CLKINVX4 U473 ( .A(n974), .Y(n1559) );
  NAND4X2 U474 ( .A(funct_regD[5]), .B(funct_regD[2]), .C(n933), .D(n939), .Y(
        n970) );
  INVX8 U475 ( .A(funct_regD[3]), .Y(n939) );
  INVX4 U476 ( .A(funct_regD[4]), .Y(n933) );
  INVX12 U477 ( .A(ALUinB[4]), .Y(n407) );
  NAND4X4 U478 ( .A(n1486), .B(n1485), .C(n1484), .D(n1483), .Y(n1487) );
  OA21X4 U479 ( .A0(n1463), .A1(n1462), .B0(n1461), .Y(n128) );
  NAND2BX4 U480 ( .AN(n278), .B(n1532), .Y(n1533) );
  OAI211X2 U481 ( .A0(n1463), .A1(n1380), .B0(n1378), .C0(n1379), .Y(
        ALUout[18]) );
  INVX3 U482 ( .A(N1003), .Y(n1380) );
  INVX20 U483 ( .A(n407), .Y(n406) );
  NAND2X6 U484 ( .A(N978), .B(n1542), .Y(n140) );
  BUFX20 U485 ( .A(n737), .Y(n313) );
  NAND3X4 U486 ( .A(n142), .B(n143), .C(n1271), .Y(ALUout[8]) );
  NAND2X1 U487 ( .A(n406), .B(n88), .Y(n1028) );
  AO22X4 U488 ( .A0(subaluinA[31]), .A1(n241), .B0(reg_lo[31]), .B1(n390), .Y(
        n1553) );
  AOI32X2 U489 ( .A0(n244), .A1(n273), .A2(n242), .B0(n287), .B1(n390), .Y(
        n1457) );
  AOI222X4 U490 ( .A0(subaluinA[5]), .A1(n241), .B0(n165), .B1(n242), .C0(n306), .C1(n390), .Y(n1230) );
  AOI222X4 U491 ( .A0(subaluinA[10]), .A1(n241), .B0(n175), .B1(n242), .C0(
        n301), .C1(n390), .Y(n1290) );
  AOI222X1 U492 ( .A0(subaluinA[12]), .A1(n241), .B0(n159), .B1(n242), .C0(
        n299), .C1(n390), .Y(n1309) );
  BUFX16 U493 ( .A(n1551), .Y(n390) );
  AND2X1 U494 ( .A(n134), .B(n268), .Y(n182) );
  CLKMX2X4 U495 ( .A(n382), .B(n1536), .S0(n1533), .Y(n1537) );
  INVX8 U496 ( .A(n214), .Y(n215) );
  OAI221X4 U497 ( .A0(n1564), .A1(n1563), .B0(N1112), .B1(n1563), .C0(n395), 
        .Y(n1572) );
  AOI222X4 U498 ( .A0(n192), .A1(n1534), .B0(n281), .B1(n389), .C0(
        subaluinA[30]), .C1(n241), .Y(n1538) );
  AOI2BB1X1 U499 ( .A0N(n391), .A1N(n192), .B0(n387), .Y(n1536) );
  CLKMX2X4 U500 ( .A(n1382), .B(n381), .S0(n1381), .Y(n1387) );
  AOI31X2 U501 ( .A0(N993), .A1(n394), .A2(n239), .B0(n1270), .Y(n1271) );
  BUFX20 U502 ( .A(ALUinA[27]), .Y(n145) );
  BUFX20 U503 ( .A(ALUinA[13]), .Y(n262) );
  NAND4X1 U504 ( .A(n1399), .B(n1398), .C(n1397), .D(n1396), .Y(n1401) );
  CLKINVX8 U505 ( .A(N1014), .Y(n129) );
  AOI2BB2X4 U506 ( .B0(N982), .B1(n1542), .A0N(n129), .A1N(n1463), .Y(n1529)
         );
  INVX3 U507 ( .A(N962), .Y(n1284) );
  AND3X4 U508 ( .A(n973), .B(n940), .C(n939), .Y(n191) );
  NAND3BX1 U509 ( .AN(n939), .B(n198), .C(n940), .Y(n756) );
  INVX6 U510 ( .A(n414), .Y(n940) );
  NAND2X2 U511 ( .A(n379), .B(n1383), .Y(n1386) );
  CLKINVX4 U512 ( .A(n1428), .Y(n1426) );
  NAND2X2 U513 ( .A(n379), .B(n1428), .Y(n1431) );
  NAND2BX2 U514 ( .AN(n271), .B(n1425), .Y(n1428) );
  AOI2BB2X4 U515 ( .B0(N1055), .B1(n170), .A0N(n1419), .A1N(n1245), .Y(n1246)
         );
  NAND3BX4 U516 ( .AN(n975), .B(n178), .C(n976), .Y(n1450) );
  BUFX20 U517 ( .A(n1548), .Y(n387) );
  INVX8 U518 ( .A(n1450), .Y(n1548) );
  OAI221X4 U519 ( .A0(n1257), .A1(n1560), .B0(n1506), .B1(n1256), .C0(n1255), 
        .Y(n1258) );
  OAI2BB2X4 U520 ( .B0(n280), .B1(n997), .A0N(n996), .A1N(n397), .Y(ALUout[1])
         );
  AND2X2 U521 ( .A(n147), .B(n277), .Y(n186) );
  OAI221X2 U522 ( .A0(N1110), .A1(n1528), .B0(n1564), .B1(n1528), .C0(n395), 
        .Y(n1530) );
  OAI211X4 U523 ( .A0(n930), .A1(n972), .B0(n944), .C0(n982), .Y(n925) );
  NAND2X2 U524 ( .A(n957), .B(n955), .Y(n930) );
  NAND3X8 U525 ( .A(n193), .B(n194), .C(n195), .Y(ALUout[12]) );
  CLKINVX6 U526 ( .A(n248), .Y(n859) );
  AOI22X4 U527 ( .A0(N1061), .A1(n152), .B0(N1093), .B1(n1443), .Y(n195) );
  AOI222X1 U528 ( .A0(subaluinA[18]), .A1(n241), .B0(n179), .B1(n242), .C0(
        n293), .C1(n389), .Y(n1373) );
  BUFX20 U529 ( .A(n1551), .Y(n389) );
  OAI32X2 U530 ( .A0(n1263), .A1(n1416), .A2(n280), .B0(n1262), .B1(n280), .Y(
        ALUout[7]) );
  AOI22X4 U531 ( .A0(N979), .A1(n1542), .B0(N1011), .B1(n1541), .Y(n1488) );
  OAI2BB2X4 U532 ( .B0(n280), .B1(n1250), .A0N(n1249), .A1N(n397), .Y(
        ALUout[6]) );
  BUFX20 U533 ( .A(ALUinA[27]), .Y(n146) );
  AOI222X4 U534 ( .A0(subaluinA[19]), .A1(n241), .B0(n182), .B1(n242), .C0(
        n292), .C1(n389), .Y(n1384) );
  AOI32X2 U535 ( .A0(N1070), .A1(n394), .A2(n170), .B0(N974), .B1(n1418), .Y(
        n1422) );
  AOI31X2 U536 ( .A0(N994), .A1(n239), .A2(n394), .B0(n1282), .Y(n1283) );
  AOI222X4 U537 ( .A0(n181), .A1(n242), .B0(n284), .B1(n389), .C0(n64), .C1(
        n241), .Y(n1498) );
  BUFX20 U538 ( .A(ALUinB[24]), .Y(n244) );
  BUFX20 U539 ( .A(ALUinB[25]), .Y(n245) );
  AOI2BB2X4 U540 ( .B0(N1006), .B1(n1541), .A0N(n1420), .A1N(n1419), .Y(n1421)
         );
  BUFX20 U541 ( .A(ALUinA[29]), .Y(n277) );
  BUFX20 U542 ( .A(ALUinB[28]), .Y(n247) );
  OAI2BB2X4 U543 ( .B0(n280), .B1(n1027), .A0N(n1026), .A1N(n397), .Y(
        ALUout[3]) );
  AOI222X2 U544 ( .A0(N1071), .A1(n152), .B0(N1103), .B1(n1443), .C0(n1433), 
        .C1(n394), .Y(n1435) );
  NAND4BX4 U545 ( .AN(n1424), .B(n1422), .C(n1423), .D(n1421), .Y(ALUout[21])
         );
  BUFX20 U546 ( .A(ALUinA[23]), .Y(n272) );
  BUFX20 U547 ( .A(ALUinA[22]), .Y(n271) );
  BUFX20 U548 ( .A(ALUinA[2]), .Y(n251) );
  BUFX20 U549 ( .A(ALUinA[30]), .Y(n278) );
  AND2X8 U550 ( .A(n138), .B(n394), .Y(ALUout[5]) );
  BUFX20 U551 ( .A(ALUinA[17]), .Y(n266) );
  NAND2X6 U552 ( .A(N1074), .B(n152), .Y(n141) );
  AND3X8 U553 ( .A(n139), .B(n140), .C(n141), .Y(n1475) );
  OR2X2 U554 ( .A(n280), .B(n1274), .Y(n142) );
  CLKINVX1 U555 ( .A(N961), .Y(n1272) );
  BUFX20 U556 ( .A(n393), .Y(n395) );
  NAND3BX4 U557 ( .AN(n923), .B(n922), .C(n929), .Y(n924) );
  BUFX20 U558 ( .A(ALUinA[0]), .Y(n249) );
  BUFX20 U559 ( .A(ALUinA[1]), .Y(n250) );
  BUFX12 U560 ( .A(n737), .Y(n312) );
  BUFX8 U561 ( .A(n825), .Y(n330) );
  BUFX3 U562 ( .A(n823), .Y(n325) );
  CLKBUFX2 U563 ( .A(n823), .Y(n326) );
  CLKBUFX2 U564 ( .A(n825), .Y(n329) );
  BUFX8 U565 ( .A(n868), .Y(n343) );
  BUFX8 U566 ( .A(n874), .Y(n351) );
  CLKBUFX2 U567 ( .A(n868), .Y(n344) );
  CLKBUFX3 U568 ( .A(n874), .Y(n352) );
  INVX2 U569 ( .A(n359), .Y(n353) );
  INVX8 U570 ( .A(n357), .Y(n356) );
  NAND3BX2 U571 ( .AN(n172), .B(n312), .C(n871), .Y(n502) );
  INVX1 U572 ( .A(n1408), .Y(n1413) );
  CLKAND2X8 U573 ( .A(n959), .B(n395), .Y(n197) );
  NAND3BX2 U574 ( .AN(n941), .B(n940), .C(n939), .Y(n942) );
  INVXL U575 ( .A(n930), .Y(n932) );
  AOI222XL U576 ( .A0(n824), .A1(n291), .B0(n293), .B1(n348), .C0(
        ALUinA_com[19]), .C1(n325), .Y(n439) );
  BUFX2 U577 ( .A(n868), .Y(n345) );
  INVX2 U578 ( .A(n907), .Y(n906) );
  INVX3 U579 ( .A(n558), .Y(n868) );
  INVX2 U580 ( .A(n413), .Y(n905) );
  AOI222XL U581 ( .A0(n824), .A1(n286), .B0(n288), .B1(n346), .C0(
        ALUinA_com[24]), .C1(n325), .Y(n424) );
  XOR2XL U582 ( .A(n955), .B(funct_regD[1]), .Y(n931) );
  NAND4X8 U583 ( .A(ALUOp_regD[2]), .B(ALUOp_regD[0]), .C(n958), .D(n197), .Y(
        n1560) );
  AOI2BB1X2 U584 ( .A0N(n392), .A1N(n1030), .B0(n387), .Y(n1031) );
  CLKBUFX2 U585 ( .A(n394), .Y(n397) );
  CLKMX2X4 U586 ( .A(n382), .B(n1288), .S0(n1289), .Y(n1293) );
  INVX3 U587 ( .A(n1018), .Y(n1015) );
  NAND2X8 U588 ( .A(n239), .B(n395), .Y(n1463) );
  CLKINVX4 U589 ( .A(n206), .Y(n199) );
  CLKMX2X2 U590 ( .A(n426), .B(n287), .S0(n374), .Y(n1170) );
  CLKINVX4 U591 ( .A(n875), .Y(n360) );
  INVX6 U592 ( .A(n842), .Y(n894) );
  CLKINVX1 U593 ( .A(n1492), .Y(n1493) );
  CLKMX2X2 U594 ( .A(n382), .B(n1307), .S0(n1308), .Y(n1312) );
  NAND2X1 U595 ( .A(n380), .B(n1277), .Y(n1280) );
  CLKINVX3 U596 ( .A(n1360), .Y(n1358) );
  BUFX16 U597 ( .A(n394), .Y(n396) );
  NAND3X4 U598 ( .A(n162), .B(n163), .C(n164), .Y(ALUout[14]) );
  AND2XL U599 ( .A(n96), .B(n251), .Y(n998) );
  NAND2BXL U600 ( .AN(n263), .B(n1328), .Y(n1331) );
  NAND2BXL U601 ( .AN(n81), .B(n1392), .Y(n1395) );
  INVX6 U602 ( .A(n385), .Y(n382) );
  NAND2X1 U603 ( .A(n1465), .B(n240), .Y(n1470) );
  AOI2BB1X1 U604 ( .A0N(n392), .A1N(n184), .B0(n387), .Y(n1239) );
  INVX1 U605 ( .A(n1256), .Y(n1253) );
  CLKAND2X8 U606 ( .A(n373), .B(n748), .Y(n171) );
  INVXL U607 ( .A(n856), .Y(n857) );
  BUFX12 U608 ( .A(n878), .Y(n373) );
  BUFX20 U609 ( .A(ALUinA[10]), .Y(n259) );
  BUFX20 U610 ( .A(ALUinA[12]), .Y(n261) );
  BUFX20 U611 ( .A(ALUinA[9]), .Y(n258) );
  NAND3X4 U612 ( .A(n187), .B(n188), .C(n189), .Y(ALUout[10]) );
  INVXL U613 ( .A(n396), .Y(n153) );
  AND2XL U614 ( .A(ALUinB[9]), .B(n86), .Y(n174) );
  CLKINVX1 U615 ( .A(n1252), .Y(n1257) );
  MX2X2 U616 ( .A(n1371), .B(n381), .S0(n1370), .Y(n1376) );
  NAND2X1 U617 ( .A(n379), .B(n1360), .Y(n1363) );
  INVXL U618 ( .A(n981), .Y(n917) );
  INVXL U619 ( .A(n980), .Y(n921) );
  MX2XL U620 ( .A(n806), .B(n289), .S0(n374), .Y(n1172) );
  AOI222XL U621 ( .A0(n352), .A1(n283), .B0(ALUinA_com[26]), .B1(n329), .C0(
        n281), .C1(n355), .Y(n518) );
  AOI222XL U622 ( .A0(n351), .A1(n289), .B0(ALUinA_com[20]), .B1(n329), .C0(
        n287), .C1(n356), .Y(n803) );
  AOI222XL U623 ( .A0(n824), .A1(n289), .B0(n291), .B1(n347), .C0(
        ALUinA_com[21]), .C1(n326), .Y(n449) );
  AOI222XL U624 ( .A0(n824), .A1(n290), .B0(n292), .B1(n348), .C0(
        ALUinA_com[20]), .C1(n325), .Y(n444) );
  AOI222XL U625 ( .A0(n351), .A1(n286), .B0(ALUinA_com[23]), .B1(n330), .C0(
        n284), .C1(n356), .Y(n428) );
  MX2XL U626 ( .A(n441), .B(n292), .S0(n375), .Y(n1175) );
  MX2XL U627 ( .A(n456), .B(n297), .S0(n375), .Y(n1180) );
  AOI222XL U628 ( .A0(n824), .A1(n296), .B0(n298), .B1(n347), .C0(
        ALUinA_com[14]), .C1(n325), .Y(n454) );
  AOI222X1 U629 ( .A0(n70), .A1(n241), .B0(n183), .B1(n242), .C0(n296), .C1(
        n389), .Y(n1341) );
  INVX1 U630 ( .A(n1533), .Y(n1539) );
  AOI222X1 U631 ( .A0(subaluinA[16]), .A1(n241), .B0(n156), .B1(n242), .C0(
        n295), .C1(n389), .Y(n1350) );
  CLKAND2X12 U632 ( .A(\stateplus2[0] ), .B(n411), .Y(n201) );
  NAND2X1 U633 ( .A(ALUinB_com[7]), .B(n320), .Y(n784) );
  NAND2X1 U634 ( .A(ALUinB_com[10]), .B(n320), .Y(n781) );
  NAND2X1 U635 ( .A(ALUinB_com[9]), .B(n320), .Y(n782) );
  NAND2X1 U636 ( .A(ALUinB_com[12]), .B(n791), .Y(n779) );
  OAI221XL U637 ( .A0(n1369), .A1(n321), .B0(n377), .B1(n33), .C0(n773), .Y(
        n1085) );
  AND2XL U638 ( .A(n1043), .B(n324), .Y(subaluinB[8]) );
  INVX8 U639 ( .A(n363), .Y(n362) );
  BUFX4 U640 ( .A(n369), .Y(n364) );
  INVX1 U641 ( .A(n310), .Y(n309) );
  AOI2BB1X2 U642 ( .A0N(n391), .A1N(n988), .B0(n387), .Y(n977) );
  INVX8 U643 ( .A(n1507), .Y(n1549) );
  INVX6 U644 ( .A(n349), .Y(n348) );
  OA22XL U645 ( .A0(n359), .A1(n729), .B0(n336), .B1(n744), .Y(n730) );
  INVX1 U646 ( .A(ALUinA_com[29]), .Y(n547) );
  BUFX4 U647 ( .A(n341), .Y(n335) );
  BUFX4 U648 ( .A(n342), .Y(n334) );
  CLKBUFX2 U649 ( .A(n340), .Y(n338) );
  CLKBUFX2 U650 ( .A(n341), .Y(n336) );
  CLKBUFX2 U651 ( .A(n340), .Y(n337) );
  INVXL U652 ( .A(ALUinA_com[1]), .Y(n872) );
  NAND3X4 U653 ( .A(n239), .B(n397), .C(N1000), .Y(n167) );
  AOI22X2 U654 ( .A0(N1064), .A1(n152), .B0(N1096), .B1(n1443), .Y(n169) );
  BUFX12 U655 ( .A(n1510), .Y(n379) );
  AOI2BB1X2 U656 ( .A0N(n392), .A1N(n183), .B0(n388), .Y(n1339) );
  NAND2BXL U657 ( .AN(n83), .B(n1407), .Y(n1408) );
  NAND2BX2 U658 ( .AN(n78), .B(n1287), .Y(n1289) );
  NAND2BX2 U659 ( .AN(n94), .B(n214), .Y(n1296) );
  NAND2XL U660 ( .A(n174), .B(n240), .Y(n1279) );
  CLKMX2X4 U661 ( .A(n383), .B(n999), .S0(n1000), .Y(n1006) );
  CLKMX2X4 U662 ( .A(n1016), .B(n383), .S0(n1019), .Y(n1017) );
  AOI2BB1X2 U663 ( .A0N(n392), .A1N(n1015), .B0(n387), .Y(n1016) );
  CLKMX2X3 U664 ( .A(n382), .B(n1276), .S0(n1277), .Y(n1281) );
  BUFX8 U665 ( .A(n1562), .Y(n393) );
  CLKINVX8 U666 ( .A(n386), .Y(n381) );
  INVX4 U667 ( .A(n410), .Y(n411) );
  INVX8 U668 ( .A(n941), .Y(n991) );
  CLKINVX3 U669 ( .A(n384), .Y(n383) );
  BUFX12 U670 ( .A(n796), .Y(n324) );
  INVX3 U671 ( .A(tempresult[18]), .Y(n671) );
  INVX3 U672 ( .A(tempresult[28]), .Y(n728) );
  INVX3 U673 ( .A(tempresult[17]), .Y(n665) );
  INVX3 U674 ( .A(tempresult[26]), .Y(n717) );
  INVX3 U675 ( .A(tempresult[24]), .Y(n707) );
  INVX3 U676 ( .A(tempresult[21]), .Y(n689) );
  INVX3 U677 ( .A(tempresult[20]), .Y(n683) );
  INVX3 U678 ( .A(tempresult[19]), .Y(n677) );
  INVX3 U679 ( .A(tempresult[29]), .Y(n736) );
  INVX3 U680 ( .A(tempresult[4]), .Y(n587) );
  INVX3 U681 ( .A(tempresult[5]), .Y(n593) );
  AND2X4 U682 ( .A(n748), .B(n743), .Y(n173) );
  INVX3 U683 ( .A(tempresult[16]), .Y(n659) );
  INVX3 U684 ( .A(tempresult[6]), .Y(n599) );
  INVX3 U685 ( .A(tempresult[8]), .Y(n611) );
  INVX3 U686 ( .A(tempresult[7]), .Y(n605) );
  INVX3 U687 ( .A(tempresult[13]), .Y(n641) );
  INVX3 U688 ( .A(tempresult[12]), .Y(n635) );
  INVX3 U689 ( .A(tempresult[10]), .Y(n623) );
  INVX3 U690 ( .A(tempresult[9]), .Y(n617) );
  INVX3 U691 ( .A(tempresult[11]), .Y(n629) );
  NAND2X2 U692 ( .A(n855), .B(n845), .Y(n876) );
  INVX1 U693 ( .A(n845), .Y(n897) );
  INVXL U694 ( .A(n902), .Y(n420) );
  NAND2BXL U695 ( .AN(n418), .B(n420), .Y(n855) );
  INVXL U696 ( .A(n748), .Y(n735) );
  INVX4 U697 ( .A(n743), .Y(n874) );
  CLKBUFX2 U698 ( .A(n878), .Y(n371) );
  CLKBUFX2 U699 ( .A(n878), .Y(n372) );
  BUFX20 U700 ( .A(ALUinA[25]), .Y(n274) );
  BUFX20 U701 ( .A(ALUinA[14]), .Y(n263) );
  AOI2BB2X4 U702 ( .B0(N964), .B1(n1303), .A0N(n28), .A1N(n153), .Y(n177) );
  AOI32X2 U703 ( .A0(N1049), .A1(n991), .A2(n967), .B0(n76), .B1(n917), .Y(
        n928) );
  NAND4X2 U704 ( .A(n1344), .B(n1343), .C(n1342), .D(n1341), .Y(n1345) );
  CLKINVX4 U705 ( .A(N954), .Y(n979) );
  NAND2XL U706 ( .A(n379), .B(n1372), .Y(n1375) );
  AOI33XL U707 ( .A0(n246), .A1(n275), .A2(n240), .B0(n246), .B1(n275), .B2(
        n242), .Y(n1484) );
  NAND2XL U708 ( .A(n181), .B(n240), .Y(n1497) );
  NAND2XL U709 ( .A(n185), .B(n240), .Y(n1397) );
  NAND2XL U710 ( .A(n379), .B(n1395), .Y(n1398) );
  NAND3BX4 U711 ( .AN(n836), .B(n200), .C(n25), .Y(n409) );
  BUFX12 U712 ( .A(n1568), .Y(n239) );
  OAI31XL U713 ( .A0(n983), .A1(n982), .A2(n981), .B0(n980), .Y(n1568) );
  NAND2BXL U714 ( .AN(n254), .B(n117), .Y(n1228) );
  NAND2XL U715 ( .A(n196), .B(n201), .Y(n418) );
  CLKMX2X2 U716 ( .A(n811), .B(n294), .S0(n374), .Y(n1177) );
  CLKMX2X2 U717 ( .A(n531), .B(n293), .S0(n374), .Y(n1176) );
  CLKMX2X2 U718 ( .A(n431), .B(n286), .S0(n375), .Y(n1169) );
  CLKMX2X2 U719 ( .A(n446), .B(n291), .S0(n375), .Y(n1174) );
  OA22XL U720 ( .A0(n313), .A1(n647), .B0(n315), .B1(n641), .Y(n644) );
  OA22XL U721 ( .A0(n365), .A1(n671), .B0(n338), .B1(n665), .Y(n642) );
  OA22XL U722 ( .A0(n563), .A1(n313), .B0(n558), .B1(n593), .Y(n561) );
  CLKMX2X2 U723 ( .A(n536), .B(n298), .S0(n374), .Y(n1181) );
  NAND2X2 U724 ( .A(n856), .B(n886), .Y(n155) );
  INVX1 U725 ( .A(n891), .Y(n893) );
  INVXL U726 ( .A(n944), .Y(n945) );
  NAND2X1 U727 ( .A(n159), .B(n240), .Y(n1310) );
  NAND2X1 U728 ( .A(n180), .B(n240), .Y(n1440) );
  NAND3BXL U729 ( .AN(n905), .B(state[6]), .C(n417), .Y(n831) );
  NAND2XL U730 ( .A(n973), .B(funct_regD[5]), .Y(n981) );
  INVX3 U731 ( .A(n1535), .Y(n386) );
  BUFX8 U732 ( .A(reg_lo[29]), .Y(n282) );
  BUFX8 U733 ( .A(reg_lo[23]), .Y(n288) );
  BUFX8 U734 ( .A(reg_lo[25]), .Y(n286) );
  BUFX8 U735 ( .A(reg_lo[27]), .Y(n284) );
  BUFX8 U736 ( .A(reg_lo[19]), .Y(n292) );
  BUFX8 U737 ( .A(reg_lo[20]), .Y(n291) );
  BUFX8 U738 ( .A(reg_lo[28]), .Y(n283) );
  BUFX8 U739 ( .A(reg_lo[22]), .Y(n289) );
  BUFX8 U740 ( .A(reg_lo[13]), .Y(n298) );
  BUFX8 U741 ( .A(reg_lo[7]), .Y(n304) );
  BUFX8 U742 ( .A(reg_lo[24]), .Y(n287) );
  NAND2X1 U743 ( .A(ALUinB_com[25]), .B(n320), .Y(n766) );
  NAND2X1 U744 ( .A(ALUinB_com[24]), .B(n320), .Y(n767) );
  NAND2X1 U745 ( .A(ALUinB_com[26]), .B(n320), .Y(n765) );
  NAND2X1 U746 ( .A(ALUinB_com[28]), .B(n320), .Y(n763) );
  NAND2X1 U747 ( .A(ALUinB_com[30]), .B(n320), .Y(n761) );
  NAND2X1 U748 ( .A(ALUinB_com[20]), .B(n320), .Y(n771) );
  NAND2X1 U749 ( .A(ALUinB_com[29]), .B(n320), .Y(n762) );
  NAND2X1 U750 ( .A(ALUinB_com[21]), .B(n320), .Y(n770) );
  NAND2X1 U751 ( .A(ALUinB_com[22]), .B(n320), .Y(n769) );
  NAND2X1 U752 ( .A(ALUinB_com[17]), .B(n791), .Y(n774) );
  NAND2X1 U753 ( .A(ALUinB_com[19]), .B(n320), .Y(n772) );
  NAND2X1 U754 ( .A(ALUinB_com[14]), .B(n791), .Y(n777) );
  INVX3 U755 ( .A(n1162), .Y(n943) );
  NAND2X1 U756 ( .A(ALUinB_com[18]), .B(n791), .Y(n773) );
  BUFX8 U757 ( .A(reg_lo[10]), .Y(n301) );
  BUFX8 U758 ( .A(reg_lo[12]), .Y(n299) );
  BUFX8 U759 ( .A(reg_lo[30]), .Y(n281) );
  BUFX8 U760 ( .A(reg_lo[11]), .Y(n300) );
  BUFX8 U761 ( .A(reg_lo[21]), .Y(n290) );
  BUFX8 U762 ( .A(reg_lo[15]), .Y(n296) );
  BUFX8 U763 ( .A(reg_lo[17]), .Y(n294) );
  BUFX8 U764 ( .A(reg_lo[9]), .Y(n302) );
  BUFX8 U765 ( .A(reg_lo[16]), .Y(n295) );
  BUFX8 U766 ( .A(reg_lo[14]), .Y(n297) );
  BUFX8 U767 ( .A(reg_lo[18]), .Y(n293) );
  BUFX8 U768 ( .A(reg_lo[26]), .Y(n285) );
  BUFX8 U769 ( .A(reg_lo[5]), .Y(n306) );
  BUFX8 U770 ( .A(reg_lo[8]), .Y(n303) );
  BUFX8 U771 ( .A(reg_lo[6]), .Y(n305) );
  AND2XL U772 ( .A(n1049), .B(n324), .Y(subaluinB[14]) );
  AND2XL U773 ( .A(n1041), .B(n324), .Y(subaluinB[6]) );
  AND2XL U774 ( .A(n1035), .B(n324), .Y(subaluinB[0]) );
  NAND2X1 U775 ( .A(ALUinB_com[13]), .B(n791), .Y(n778) );
  NAND2X1 U776 ( .A(ALUinB_com[16]), .B(n791), .Y(n775) );
  AOI222XL U777 ( .A0(lo_com[8]), .A1(n371), .B0(n299), .B1(n361), .C0(n300), 
        .C1(n331), .Y(n537) );
  AOI222XL U778 ( .A0(lo_com[17]), .A1(n371), .B0(n290), .B1(n361), .C0(n291), 
        .C1(n332), .Y(n807) );
  AOI222XL U779 ( .A0(lo_com[23]), .A1(n371), .B0(n284), .B1(n361), .C0(n285), 
        .C1(n331), .Y(n522) );
  AOI222XL U780 ( .A0(lo_com[15]), .A1(n372), .B0(n292), .B1(n362), .C0(n293), 
        .C1(n332), .Y(n457) );
  AOI222XL U781 ( .A0(lo_com[11]), .A1(n372), .B0(n296), .B1(n362), .C0(n297), 
        .C1(n332), .Y(n477) );
  AOI222XL U782 ( .A0(lo_com[25]), .A1(n373), .B0(n282), .B1(n362), .C0(n283), 
        .C1(n332), .Y(n427) );
  AND2XL U783 ( .A(n1063), .B(n323), .Y(subaluinB[28]) );
  NAND2X1 U784 ( .A(ALUinB_com[15]), .B(n791), .Y(n776) );
  AND2XL U785 ( .A(n1057), .B(n323), .Y(subaluinB[22]) );
  NAND2XL U786 ( .A(state[2]), .B(n836), .Y(n844) );
  CLKINVX1 U787 ( .A(N955), .Y(n1010) );
  CLKBUFX3 U788 ( .A(n370), .Y(n363) );
  CLKBUFX2 U789 ( .A(n912), .Y(n376) );
  CLKBUFX2 U790 ( .A(n912), .Y(n377) );
  CLKBUFX3 U791 ( .A(n234), .Y(n227) );
  CLKBUFX3 U792 ( .A(n232), .Y(n228) );
  CLKBUFX3 U793 ( .A(n232), .Y(n230) );
  CLKBUFX3 U794 ( .A(n233), .Y(n229) );
  CLKBUFX3 U795 ( .A(n233), .Y(n224) );
  CLKBUFX3 U796 ( .A(n233), .Y(n225) );
  CLKBUFX3 U797 ( .A(n234), .Y(n226) );
  CLKBUFX3 U798 ( .A(n232), .Y(n231) );
  AOI2BB1X1 U799 ( .A0N(n392), .A1N(n160), .B0(n387), .Y(n1298) );
  AOI2BB1X1 U800 ( .A0N(n392), .A1N(n161), .B0(n387), .Y(n1330) );
  BUFX20 U801 ( .A(n1549), .Y(n242) );
  NAND2X1 U802 ( .A(n379), .B(n1349), .Y(n1352) );
  CLKINVX1 U803 ( .A(n1340), .Y(n1338) );
  CLKINVX1 U804 ( .A(n1240), .Y(n1238) );
  CLKINVX1 U805 ( .A(n1372), .Y(n1370) );
  CLKINVX1 U806 ( .A(n1395), .Y(n1393) );
  CLKINVX1 U807 ( .A(n1331), .Y(n1329) );
  CLKINVX1 U808 ( .A(n1296), .Y(n1297) );
  BUFX12 U809 ( .A(n1548), .Y(n388) );
  CLKBUFX3 U810 ( .A(n171), .Y(n317) );
  CLKBUFX3 U811 ( .A(n171), .Y(n318) );
  CLKBUFX3 U812 ( .A(n171), .Y(n319) );
  CLKBUFX3 U813 ( .A(n340), .Y(n339) );
  CLKINVX1 U814 ( .A(n876), .Y(n369) );
  CLKINVX1 U815 ( .A(n876), .Y(n370) );
  CLKINVX1 U816 ( .A(tempresult[32]), .Y(n744) );
  NAND2BXL U817 ( .AN(n901), .B(n90), .Y(n549) );
  CLKINVX1 U818 ( .A(n855), .Y(n858) );
  CLKBUFX3 U819 ( .A(n173), .Y(n310) );
  INVX3 U820 ( .A(n173), .Y(n307) );
  INVX3 U821 ( .A(n311), .Y(n308) );
  CLKBUFX3 U822 ( .A(n173), .Y(n311) );
  CLKBUFX3 U823 ( .A(n234), .Y(n223) );
  NAND2X1 U824 ( .A(n404), .B(n89), .Y(n1018) );
  NAND2XL U825 ( .A(n860), .B(n1546), .Y(n909) );
  NAND2BX1 U826 ( .AN(n272), .B(n1436), .Y(n1438) );
  NAND2X1 U827 ( .A(n1316), .B(n1315), .Y(n1321) );
  NAND2BX1 U828 ( .AN(n266), .B(n235), .Y(n1360) );
  NAND2BX1 U829 ( .AN(n146), .B(n1491), .Y(n1492) );
  AND2X2 U830 ( .A(n216), .B(n94), .Y(n160) );
  AOI2BB1XL U831 ( .A0N(n391), .A1N(n185), .B0(n388), .Y(n1394) );
  CLKINVX1 U832 ( .A(n277), .Y(n1522) );
  NAND3X6 U833 ( .A(n239), .B(n396), .C(N999), .Y(n162) );
  AOI22X4 U834 ( .A0(N967), .A1(n1337), .B0(n1336), .B1(n396), .Y(n163) );
  NAND2X1 U835 ( .A(N956), .B(n238), .Y(n1023) );
  NAND2XL U836 ( .A(n157), .B(n240), .Y(n1267) );
  NAND2XL U837 ( .A(n156), .B(n240), .Y(n1351) );
  CLKMX2X2 U838 ( .A(n382), .B(n1229), .S0(n1228), .Y(n1232) );
  CLKMX2X2 U839 ( .A(n381), .B(n1437), .S0(n1438), .Y(n1442) );
  AOI22X4 U840 ( .A0(N968), .A1(n1346), .B0(n1345), .B1(n396), .Y(n168) );
  NAND2X1 U841 ( .A(n902), .B(n904), .Y(n916) );
  INVXL U842 ( .A(n955), .Y(n956) );
  AO21XL U843 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1303) );
  AO21XL U844 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1337) );
  AO21XL U845 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1346) );
  AO21XL U846 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1295) );
  AO21XL U847 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1314) );
  AO21XL U848 ( .A0(n1354), .A1(n396), .B0(n238), .Y(n1325) );
  NAND3BXL U849 ( .AN(n941), .B(n760), .C(n90), .Y(n408) );
  NAND3BXL U850 ( .AN(n90), .B(n973), .C(n760), .Y(n746) );
  AOI222XL U851 ( .A0(tempresult[4]), .A1(n355), .B0(tempresult[7]), .B1(n344), 
        .C0(tempresult[3]), .C1(n824), .Y(n571) );
  AOI222XL U852 ( .A0(tempresult[16]), .A1(n354), .B0(tempresult[19]), .B1(
        n344), .C0(tempresult[15]), .C1(n824), .Y(n643) );
  AOI222XL U853 ( .A0(tempresult[15]), .A1(n354), .B0(tempresult[18]), .B1(
        n344), .C0(tempresult[14]), .C1(n824), .Y(n637) );
  AOI222XL U854 ( .A0(tempresult[14]), .A1(n354), .B0(tempresult[17]), .B1(
        n344), .C0(tempresult[13]), .C1(n824), .Y(n631) );
  AOI222XL U855 ( .A0(tempresult[13]), .A1(n354), .B0(tempresult[16]), .B1(
        n344), .C0(tempresult[12]), .C1(n824), .Y(n625) );
  AOI222XL U856 ( .A0(tempresult[11]), .A1(n354), .B0(tempresult[14]), .B1(
        n344), .C0(tempresult[10]), .C1(n327), .Y(n613) );
  AOI222XL U857 ( .A0(tempresult[10]), .A1(n354), .B0(tempresult[13]), .B1(
        n344), .C0(tempresult[9]), .C1(n824), .Y(n607) );
  AOI222XL U858 ( .A0(tempresult[5]), .A1(n355), .B0(tempresult[8]), .B1(n344), 
        .C0(tempresult[4]), .C1(n824), .Y(n577) );
  AOI222XL U859 ( .A0(tempresult[17]), .A1(n354), .B0(tempresult[20]), .B1(
        n344), .C0(tempresult[16]), .C1(n824), .Y(n649) );
  AOI222XL U860 ( .A0(tempresult[9]), .A1(n354), .B0(tempresult[12]), .B1(n344), .C0(tempresult[8]), .C1(n824), .Y(n601) );
  AOI222XL U861 ( .A0(tempresult[8]), .A1(n354), .B0(tempresult[11]), .B1(n344), .C0(tempresult[7]), .C1(n824), .Y(n595) );
  AOI222XL U862 ( .A0(tempresult[7]), .A1(n354), .B0(tempresult[10]), .B1(n345), .C0(tempresult[6]), .C1(n824), .Y(n589) );
  AOI222XL U863 ( .A0(tempresult[6]), .A1(n354), .B0(tempresult[9]), .B1(n345), 
        .C0(tempresult[5]), .C1(n824), .Y(n583) );
  AOI222XL U864 ( .A0(tempresult[24]), .A1(n353), .B0(tempresult[27]), .B1(
        n343), .C0(tempresult[23]), .C1(n824), .Y(n691) );
  AOI222XL U865 ( .A0(tempresult[21]), .A1(n353), .B0(tempresult[24]), .B1(
        n343), .C0(tempresult[20]), .C1(n824), .Y(n673) );
  AOI222XL U866 ( .A0(tempresult[20]), .A1(n353), .B0(tempresult[23]), .B1(
        n343), .C0(tempresult[19]), .C1(n824), .Y(n667) );
  AOI222XL U867 ( .A0(tempresult[3]), .A1(n355), .B0(tempresult[6]), .B1(n344), 
        .C0(tempresult[2]), .C1(n824), .Y(n565) );
  AOI222XL U868 ( .A0(tempresult[29]), .A1(n353), .B0(tempresult[32]), .B1(
        n343), .C0(tempresult[28]), .C1(n824), .Y(n719) );
  AOI222XL U869 ( .A0(tempresult[26]), .A1(n353), .B0(tempresult[29]), .B1(
        n343), .C0(tempresult[25]), .C1(n824), .Y(n703) );
  AOI222XL U870 ( .A0(tempresult[25]), .A1(n353), .B0(tempresult[28]), .B1(
        n343), .C0(tempresult[24]), .C1(n824), .Y(n697) );
  AOI222XL U871 ( .A0(tempresult[18]), .A1(n353), .B0(tempresult[21]), .B1(
        n343), .C0(tempresult[17]), .C1(n824), .Y(n655) );
  CLKBUFX3 U872 ( .A(n360), .Y(n358) );
  CLKBUFX3 U873 ( .A(n360), .Y(n357) );
  CLKBUFX3 U874 ( .A(n360), .Y(n359) );
  CLKINVX1 U875 ( .A(ALUinA_com[31]), .Y(n745) );
  CLKINVX1 U876 ( .A(n155), .Y(n341) );
  CLKINVX1 U877 ( .A(n155), .Y(n340) );
  CLKINVX1 U878 ( .A(n155), .Y(n342) );
  NAND3BXL U879 ( .AN(n941), .B(n279), .C(n760), .Y(n873) );
  CLKINVX1 U880 ( .A(tempresult[3]), .Y(n581) );
  NAND2XL U881 ( .A(n760), .B(n973), .Y(n901) );
  CLKINVX1 U882 ( .A(tempresult[1]), .Y(n569) );
  CLKINVX1 U883 ( .A(tempresult[2]), .Y(n575) );
  INVX3 U884 ( .A(n350), .Y(n346) );
  INVX3 U885 ( .A(n349), .Y(n347) );
  AOI2BB1XL U886 ( .A0N(n280), .A1N(n1566), .B0(n238), .Y(n1285) );
  AOI2BB1XL U887 ( .A0N(n280), .A1N(n1566), .B0(n238), .Y(n1273) );
  AND3XL U888 ( .A(n920), .B(n962), .C(n202), .Y(n926) );
  CLKINVX1 U889 ( .A(n925), .Y(n922) );
  AND2XL U890 ( .A(n126), .B(n78), .Y(n175) );
  NAND2X1 U891 ( .A(n1507), .B(n1506), .Y(n1534) );
  AOI22X4 U892 ( .A0(N966), .A1(n1325), .B0(n1324), .B1(n396), .Y(n176) );
  OA22XL U893 ( .A0(n1505), .A1(n1482), .B0(n1503), .B1(n1481), .Y(n1483) );
  OA22XL U894 ( .A0(n1505), .A1(n1504), .B0(n1503), .B1(n1134), .Y(n1516) );
  OA22XL U895 ( .A0(n1505), .A1(n1002), .B0(n1503), .B1(n1160), .Y(n1003) );
  AOI2BB1XL U896 ( .A0N(n280), .A1N(n1566), .B0(n238), .Y(n1567) );
  OA22XL U897 ( .A0(n1506), .A1(n1001), .B0(n1507), .B1(n1001), .Y(n1004) );
  NAND2XL U898 ( .A(n182), .B(n240), .Y(n1385) );
  NAND2XL U899 ( .A(n179), .B(n240), .Y(n1374) );
  NAND2XL U900 ( .A(n15), .B(n240), .Y(n1430) );
  AND2XL U901 ( .A(n115), .B(n264), .Y(n183) );
  NAND2XL U902 ( .A(n160), .B(n240), .Y(n1300) );
  NAND2XL U903 ( .A(n379), .B(n1340), .Y(n1343) );
  NAND2XL U904 ( .A(n183), .B(n240), .Y(n1342) );
  NAND2X1 U905 ( .A(n380), .B(n1331), .Y(n1334) );
  NAND2XL U906 ( .A(n161), .B(n240), .Y(n1333) );
  NAND4X1 U907 ( .A(n1244), .B(n1243), .C(n1242), .D(n1241), .Y(n1248) );
  NAND2XL U908 ( .A(n184), .B(n240), .Y(n1242) );
  AOI22X4 U909 ( .A0(N963), .A1(n1295), .B0(n1294), .B1(n396), .Y(n188) );
  AND4X4 U910 ( .A(n954), .B(n920), .C(n959), .D(n923), .Y(n190) );
  NAND3BXL U911 ( .AN(n983), .B(n984), .C(n967), .Y(n968) );
  BUFX20 U912 ( .A(ALUinA[24]), .Y(n273) );
  BUFX20 U913 ( .A(ALUinA[4]), .Y(n253) );
  BUFX20 U914 ( .A(ALUinA[16]), .Y(n265) );
  INVX20 U915 ( .A(n399), .Y(n398) );
  BUFX20 U916 ( .A(ALUinA[31]), .Y(n279) );
  CLKBUFX3 U917 ( .A(n386), .Y(n385) );
  CLKBUFX3 U918 ( .A(n386), .Y(n384) );
  INVX1 U919 ( .A(n1466), .Y(n1467) );
  CLKMX2X2 U920 ( .A(n1479), .B(n381), .S0(n1478), .Y(n1486) );
  AND2XL U921 ( .A(n246), .B(n275), .Y(n1476) );
  OAI222XL U922 ( .A0(n1505), .A1(n1129), .B0(n1507), .B1(n986), .C0(n1503), 
        .C1(n1161), .Y(n990) );
  AND3XL U923 ( .A(n240), .B(n279), .C(n248), .Y(n1554) );
  NAND2BXL U924 ( .AN(n89), .B(n405), .Y(n1014) );
  AND3XL U925 ( .A(n244), .B(n273), .C(n240), .Y(n1454) );
  AND3XL U926 ( .A(n243), .B(n262), .C(n240), .Y(n1320) );
  NAND3X6 U927 ( .A(n239), .B(n397), .C(N997), .Y(n193) );
  AOI22X4 U928 ( .A0(N965), .A1(n1314), .B0(n1313), .B1(n396), .Y(n194) );
  NAND3BXL U929 ( .AN(n19), .B(n196), .C(n411), .Y(n907) );
  NAND2XL U930 ( .A(n938), .B(n941), .Y(n755) );
  CLKINVX1 U931 ( .A(n831), .Y(n911) );
  NOR2X2 U932 ( .A(n409), .B(n199), .Y(n198) );
  BUFX20 U933 ( .A(n1550), .Y(n240) );
  BUFX20 U934 ( .A(n1565), .Y(n238) );
  NAND2X1 U935 ( .A(n871), .B(n831), .Y(n898) );
  NAND3BX1 U936 ( .AN(n902), .B(n910), .C(n1013), .Y(n845) );
  OAI222XL U937 ( .A0(n556), .A1(n743), .B0(n359), .B1(n569), .C0(n363), .C1(
        n581), .Y(n550) );
  NAND2X1 U938 ( .A(n205), .B(n90), .Y(n748) );
  NAND2X1 U939 ( .A(n1129), .B(n1002), .Y(n902) );
  AOI222XL U940 ( .A0(lo_com[24]), .A1(n372), .B0(n283), .B1(n362), .C0(n284), 
        .C1(n331), .Y(n422) );
  AOI222XL U941 ( .A0(lo_com[18]), .A1(n371), .B0(n289), .B1(n361), .C0(n290), 
        .C1(n331), .Y(n527) );
  AOI222XL U942 ( .A0(lo_com[12]), .A1(n371), .B0(n295), .B1(n361), .C0(n296), 
        .C1(n331), .Y(n812) );
  AOI222XL U943 ( .A0(lo_com[4]), .A1(n372), .B0(n303), .B1(n362), .C0(n304), 
        .C1(n332), .Y(n482) );
  AOI222XL U944 ( .A0(lo_com[10]), .A1(n372), .B0(n297), .B1(n362), .C0(n298), 
        .C1(n332), .Y(n472) );
  AOI222XL U945 ( .A0(n352), .A1(n281), .B0(ALUinA_com[28]), .B1(n330), .C0(
        tempresult[0]), .C1(n355), .Y(n508) );
  AOI222XL U946 ( .A0(n351), .A1(n288), .B0(ALUinA_com[21]), .B1(n329), .C0(
        n286), .C1(n355), .Y(n523) );
  AOI222XL U947 ( .A0(n351), .A1(n293), .B0(ALUinA_com[16]), .B1(n329), .C0(
        n291), .C1(n355), .Y(n528) );
  AOI222XL U948 ( .A0(n351), .A1(n298), .B0(ALUinA_com[11]), .B1(n329), .C0(
        n296), .C1(n355), .Y(n533) );
  AOI222XL U949 ( .A0(n351), .A1(n303), .B0(ALUinA_com[6]), .B1(n329), .C0(
        n301), .C1(n355), .Y(n538) );
  AOI222XL U950 ( .A0(n351), .A1(n285), .B0(ALUinA_com[24]), .B1(n330), .C0(
        n283), .C1(n356), .Y(n433) );
  AOI222XL U951 ( .A0(n351), .A1(n290), .B0(ALUinA_com[19]), .B1(n330), .C0(
        n288), .C1(n356), .Y(n448) );
  AOI222XL U952 ( .A0(n351), .A1(n291), .B0(ALUinA_com[18]), .B1(n330), .C0(
        n289), .C1(n356), .Y(n443) );
  AOI222XL U953 ( .A0(n351), .A1(n292), .B0(ALUinA_com[17]), .B1(n330), .C0(
        n290), .C1(n356), .Y(n438) );
  AOI222XL U954 ( .A0(n352), .A1(n297), .B0(ALUinA_com[12]), .B1(n330), .C0(
        n295), .C1(n356), .Y(n453) );
  AOI222XL U955 ( .A0(n352), .A1(n295), .B0(ALUinA_com[14]), .B1(n330), .C0(
        n293), .C1(n356), .Y(n463) );
  AOI222XL U956 ( .A0(n352), .A1(n296), .B0(ALUinA_com[13]), .B1(n330), .C0(
        n294), .C1(n356), .Y(n458) );
  AOI222XL U957 ( .A0(n352), .A1(n300), .B0(ALUinA_com[9]), .B1(n330), .C0(
        n298), .C1(n356), .Y(n478) );
  AOI222XL U958 ( .A0(n352), .A1(n301), .B0(ALUinA_com[8]), .B1(n330), .C0(
        n299), .C1(n356), .Y(n473) );
  AOI222XL U959 ( .A0(n352), .A1(n302), .B0(ALUinA_com[7]), .B1(n330), .C0(
        n300), .C1(n356), .Y(n468) );
  AOI222XL U960 ( .A0(n352), .A1(n305), .B0(ALUinA_com[4]), .B1(n330), .C0(
        n303), .C1(n356), .Y(n493) );
  AOI222XL U961 ( .A0(n352), .A1(n306), .B0(ALUinA_com[3]), .B1(n330), .C0(
        n304), .C1(n356), .Y(n488) );
  AOI222XL U962 ( .A0(n351), .A1(n284), .B0(ALUinA_com[25]), .B1(n329), .C0(
        n282), .C1(n356), .Y(n798) );
  AOI222XL U963 ( .A0(n351), .A1(n287), .B0(ALUinA_com[22]), .B1(n329), .C0(
        n285), .C1(n356), .Y(n423) );
  AOI222XL U964 ( .A0(n352), .A1(n294), .B0(ALUinA_com[15]), .B1(n329), .C0(
        n292), .C1(n356), .Y(n808) );
  AOI222XL U965 ( .A0(n351), .A1(n299), .B0(ALUinA_com[10]), .B1(n329), .C0(
        n297), .C1(n356), .Y(n813) );
  AOI222XL U966 ( .A0(n351), .A1(n304), .B0(ALUinA_com[5]), .B1(n329), .C0(
        n302), .C1(n356), .Y(n818) );
  NAND2XL U967 ( .A(n845), .B(n842), .Y(n864) );
  NAND2XL U968 ( .A(n205), .B(n1558), .Y(n504) );
  NAND2X1 U969 ( .A(n934), .B(n933), .Y(n947) );
  AOI2BB1XL U970 ( .A0N(n906), .A1N(n892), .B0(n1013), .Y(n501) );
  AOI2BB1XL U971 ( .A0N(n734), .A1N(n316), .B0(n556), .Y(n557) );
  NAND4X1 U972 ( .A(n562), .B(n561), .C(n560), .D(n559), .Y(n1226) );
  OA22XL U973 ( .A0(n366), .A1(n587), .B0(n336), .B1(n581), .Y(n559) );
  NAND4X1 U974 ( .A(n727), .B(n726), .C(n725), .D(n724), .Y(n1221) );
  OA22XL U975 ( .A0(n312), .A1(n728), .B0(n314), .B1(n723), .Y(n726) );
  OA22XL U976 ( .A0(n366), .A1(n744), .B0(n336), .B1(n729), .Y(n724) );
  AOI222XL U977 ( .A0(n735), .A1(n722), .B0(n734), .B1(n64), .C0(hi_com[28]), 
        .C1(n319), .Y(n727) );
  NAND4X1 U978 ( .A(n573), .B(n572), .C(n571), .D(n570), .Y(n1195) );
  OA22XL U979 ( .A0(n313), .A1(n575), .B0(n314), .B1(n569), .Y(n572) );
  AOI222XL U980 ( .A0(hi_com[2]), .A1(n319), .B0(n307), .B1(n574), .C0(n734), 
        .C1(n568), .Y(n573) );
  OA22XL U981 ( .A0(n367), .A1(n599), .B0(n336), .B1(n593), .Y(n570) );
  NAND4X1 U982 ( .A(n645), .B(n644), .C(n643), .D(n642), .Y(n1207) );
  AOI222XL U983 ( .A0(hi_com[14]), .A1(n318), .B0(n308), .B1(n646), .C0(n734), 
        .C1(n640), .Y(n645) );
  NAND4X1 U984 ( .A(n639), .B(n638), .C(n637), .D(n636), .Y(n1206) );
  OA22XL U985 ( .A0(n313), .A1(n641), .B0(n315), .B1(n635), .Y(n638) );
  OA22XL U986 ( .A0(n366), .A1(n665), .B0(n337), .B1(n659), .Y(n636) );
  AOI222XL U987 ( .A0(hi_com[13]), .A1(n318), .B0(n307), .B1(n640), .C0(n734), 
        .C1(n634), .Y(n639) );
  NAND4X1 U988 ( .A(n633), .B(n632), .C(n631), .D(n630), .Y(n1205) );
  OA22XL U989 ( .A0(n313), .A1(n635), .B0(n315), .B1(n629), .Y(n632) );
  AOI222XL U990 ( .A0(hi_com[12]), .A1(n318), .B0(n307), .B1(n634), .C0(n734), 
        .C1(n67), .Y(n633) );
  NAND4X1 U991 ( .A(n627), .B(n626), .C(n625), .D(n624), .Y(n1204) );
  OA22XL U992 ( .A0(n313), .A1(n629), .B0(n315), .B1(n623), .Y(n626) );
  AOI222XL U993 ( .A0(hi_com[11]), .A1(n318), .B0(n307), .B1(n67), .C0(n734), 
        .C1(n622), .Y(n627) );
  AOI222XL U994 ( .A0(hi_com[10]), .A1(n318), .B0(n307), .B1(n622), .C0(n734), 
        .C1(n616), .Y(n621) );
  NAND4X1 U995 ( .A(n615), .B(n614), .C(n613), .D(n612), .Y(n1202) );
  OA22XL U996 ( .A0(n313), .A1(n617), .B0(n315), .B1(n611), .Y(n614) );
  OA22XL U997 ( .A0(n366), .A1(n641), .B0(n337), .B1(n635), .Y(n612) );
  AOI222XL U998 ( .A0(hi_com[9]), .A1(n318), .B0(n307), .B1(n616), .C0(n734), 
        .C1(n610), .Y(n615) );
  NAND4X1 U999 ( .A(n609), .B(n608), .C(n607), .D(n606), .Y(n1201) );
  OA22XL U1000 ( .A0(n313), .A1(n611), .B0(n315), .B1(n605), .Y(n608) );
  OA22XL U1001 ( .A0(n367), .A1(n635), .B0(n338), .B1(n629), .Y(n606) );
  AOI222XL U1002 ( .A0(hi_com[8]), .A1(n318), .B0(n307), .B1(n610), .C0(n734), 
        .C1(n604), .Y(n609) );
  NAND4X1 U1003 ( .A(n579), .B(n578), .C(n577), .D(n576), .Y(n1196) );
  OA22XL U1004 ( .A0(n313), .A1(n581), .B0(n314), .B1(n575), .Y(n578) );
  AOI222XL U1005 ( .A0(hi_com[3]), .A1(n319), .B0(n307), .B1(n580), .C0(n734), 
        .C1(n574), .Y(n579) );
  OA22XL U1006 ( .A0(n367), .A1(n605), .B0(n336), .B1(n599), .Y(n576) );
  OA22XL U1007 ( .A0(n365), .A1(n677), .B0(n338), .B1(n671), .Y(n648) );
  AOI222XL U1008 ( .A0(hi_com[15]), .A1(n317), .B0(n308), .B1(n70), .C0(n734), 
        .C1(n646), .Y(n651) );
  NAND4X1 U1009 ( .A(n603), .B(n602), .C(n601), .D(n600), .Y(n1200) );
  OA22XL U1010 ( .A0(n313), .A1(n605), .B0(n315), .B1(n599), .Y(n602) );
  OA22XL U1011 ( .A0(n367), .A1(n629), .B0(n336), .B1(n623), .Y(n600) );
  AOI222XL U1012 ( .A0(hi_com[7]), .A1(n318), .B0(n307), .B1(n604), .C0(n734), 
        .C1(n598), .Y(n603) );
  NAND4X1 U1013 ( .A(n597), .B(n596), .C(n595), .D(n594), .Y(n1199) );
  OA22XL U1014 ( .A0(n313), .A1(n599), .B0(n315), .B1(n593), .Y(n596) );
  OA22XL U1015 ( .A0(n367), .A1(n623), .B0(n336), .B1(n617), .Y(n594) );
  AOI222XL U1016 ( .A0(hi_com[6]), .A1(n318), .B0(n307), .B1(n598), .C0(n734), 
        .C1(n592), .Y(n597) );
  NAND4X1 U1017 ( .A(n591), .B(n590), .C(n589), .D(n588), .Y(n1198) );
  OA22XL U1018 ( .A0(n313), .A1(n593), .B0(n314), .B1(n587), .Y(n590) );
  OA22XL U1019 ( .A0(n367), .A1(n617), .B0(n339), .B1(n611), .Y(n588) );
  AOI222XL U1020 ( .A0(hi_com[5]), .A1(n318), .B0(n307), .B1(n592), .C0(n734), 
        .C1(n586), .Y(n591) );
  NAND4X1 U1021 ( .A(n585), .B(n584), .C(n583), .D(n582), .Y(n1197) );
  OA22XL U1022 ( .A0(n313), .A1(n587), .B0(n314), .B1(n581), .Y(n584) );
  OA22XL U1023 ( .A0(n367), .A1(n611), .B0(n339), .B1(n605), .Y(n582) );
  AOI222XL U1024 ( .A0(hi_com[4]), .A1(n318), .B0(n307), .B1(n586), .C0(n734), 
        .C1(n580), .Y(n585) );
  OA22XL U1025 ( .A0(n312), .A1(n723), .B0(n314), .B1(n717), .Y(n720) );
  OA22XL U1026 ( .A0(n367), .A1(n729), .B0(n336), .B1(n747), .Y(n718) );
  AOI222XL U1027 ( .A0(hi_com[27]), .A1(n317), .B0(n309), .B1(n64), .C0(n734), 
        .C1(subaluinA[26]), .Y(n721) );
  NAND4X1 U1028 ( .A(n716), .B(n715), .C(n714), .D(n713), .Y(n1219) );
  OA22XL U1029 ( .A0(n312), .A1(n717), .B0(n314), .B1(n712), .Y(n715) );
  OA22XL U1030 ( .A0(n364), .A1(n747), .B0(n335), .B1(n736), .Y(n713) );
  AOI222XL U1031 ( .A0(hi_com[26]), .A1(n317), .B0(n308), .B1(subaluinA[26]), 
        .C0(n734), .C1(n63), .Y(n716) );
  OA22XL U1032 ( .A0(n366), .A1(n736), .B0(n337), .B1(n728), .Y(n708) );
  AOI222XL U1033 ( .A0(hi_com[25]), .A1(n317), .B0(n308), .B1(n63), .C0(n734), 
        .C1(n706), .Y(n711) );
  NAND4X1 U1034 ( .A(n705), .B(n704), .C(n703), .D(n702), .Y(n1217) );
  AOI222XL U1035 ( .A0(hi_com[24]), .A1(n317), .B0(n308), .B1(n706), .C0(n734), 
        .C1(n700), .Y(n705) );
  NAND4X1 U1036 ( .A(n699), .B(n698), .C(n697), .D(n696), .Y(n1216) );
  OA22XL U1037 ( .A0(n312), .A1(n701), .B0(n314), .B1(n695), .Y(n698) );
  OA22XL U1038 ( .A0(n366), .A1(n723), .B0(n334), .B1(n717), .Y(n696) );
  AOI222XL U1039 ( .A0(hi_com[23]), .A1(n318), .B0(n308), .B1(n700), .C0(n734), 
        .C1(n694), .Y(n699) );
  NAND4X1 U1040 ( .A(n693), .B(n692), .C(n691), .D(n690), .Y(n1215) );
  OA22XL U1041 ( .A0(n313), .A1(n695), .B0(n314), .B1(n689), .Y(n692) );
  AOI222XL U1042 ( .A0(hi_com[22]), .A1(n317), .B0(n308), .B1(n694), .C0(n734), 
        .C1(n688), .Y(n693) );
  NAND4X1 U1043 ( .A(n687), .B(n686), .C(n685), .D(n684), .Y(n1214) );
  OA22XL U1044 ( .A0(n312), .A1(n689), .B0(n314), .B1(n683), .Y(n686) );
  OA22XL U1045 ( .A0(n367), .A1(n712), .B0(n339), .B1(n707), .Y(n684) );
  AOI222XL U1046 ( .A0(hi_com[21]), .A1(n317), .B0(n308), .B1(n688), .C0(n734), 
        .C1(n682), .Y(n687) );
  NAND4X1 U1047 ( .A(n681), .B(n680), .C(n679), .D(n678), .Y(n1213) );
  OA22XL U1048 ( .A0(n312), .A1(n683), .B0(n314), .B1(n677), .Y(n680) );
  AOI222XL U1049 ( .A0(hi_com[20]), .A1(n317), .B0(n308), .B1(n682), .C0(n734), 
        .C1(n676), .Y(n681) );
  OA22XL U1050 ( .A0(n312), .A1(n677), .B0(n314), .B1(n671), .Y(n674) );
  OA22XL U1051 ( .A0(n365), .A1(n701), .B0(n339), .B1(n695), .Y(n672) );
  AOI222XL U1052 ( .A0(hi_com[19]), .A1(n317), .B0(n308), .B1(n676), .C0(n734), 
        .C1(n670), .Y(n675) );
  OA22XL U1053 ( .A0(n312), .A1(n671), .B0(n314), .B1(n665), .Y(n668) );
  OA22XL U1054 ( .A0(n365), .A1(n695), .B0(n338), .B1(n689), .Y(n666) );
  AOI222XL U1055 ( .A0(hi_com[18]), .A1(n317), .B0(n308), .B1(n670), .C0(n734), 
        .C1(n664), .Y(n669) );
  NAND4X1 U1056 ( .A(n663), .B(n662), .C(n661), .D(n660), .Y(n1210) );
  OA22XL U1057 ( .A0(n312), .A1(n665), .B0(n315), .B1(n659), .Y(n662) );
  OA22XL U1058 ( .A0(n365), .A1(n689), .B0(n338), .B1(n683), .Y(n660) );
  AOI222XL U1059 ( .A0(hi_com[17]), .A1(n317), .B0(n308), .B1(n664), .C0(n734), 
        .C1(n658), .Y(n663) );
  NAND4X1 U1060 ( .A(n657), .B(n656), .C(n655), .D(n654), .Y(n1209) );
  OA22XL U1061 ( .A0(n365), .A1(n683), .B0(n338), .B1(n677), .Y(n654) );
  AOI222XL U1062 ( .A0(hi_com[16]), .A1(n317), .B0(n308), .B1(n658), .C0(n734), 
        .C1(n70), .Y(n657) );
  NAND4X1 U1063 ( .A(n567), .B(n566), .C(n565), .D(n564), .Y(n1194) );
  OA22XL U1064 ( .A0(n313), .A1(n569), .B0(n563), .B1(n314), .Y(n566) );
  AOI222XL U1065 ( .A0(hi_com[1]), .A1(n319), .B0(n307), .B1(n568), .C0(n734), 
        .C1(n943), .Y(n567) );
  OA22XL U1066 ( .A0(n365), .A1(n593), .B0(n336), .B1(n587), .Y(n564) );
  NAND4XL U1067 ( .A(n901), .B(n909), .C(n900), .D(n899), .Y(state_next[6]) );
  AOI222XL U1068 ( .A0(n897), .A1(n896), .B0(n895), .B1(n894), .C0(n893), .C1(
        n892), .Y(n900) );
  NAND2X1 U1069 ( .A(stateplus1[6]), .B(n898), .Y(n899) );
  CLKINVX1 U1070 ( .A(n890), .Y(n895) );
  AO21XL U1071 ( .A0(n892), .A1(n26), .B0(n894), .Y(n885) );
  NAND2XL U1072 ( .A(n499), .B(n831), .Y(n870) );
  INVXL U1073 ( .A(n416), .Y(n412) );
  CLKMX2X2 U1074 ( .A(n451), .B(n290), .S0(n375), .Y(n1173) );
  NAND4X1 U1075 ( .A(n450), .B(n449), .C(n448), .D(n447), .Y(n451) );
  AOI222XL U1076 ( .A0(n822), .A1(n268), .B0(n869), .B1(n83), .C0(n343), .C1(
        n285), .Y(n450) );
  AOI222XL U1077 ( .A0(lo_com[21]), .A1(n373), .B0(n286), .B1(n362), .C0(n287), 
        .C1(n333), .Y(n447) );
  NAND4X1 U1078 ( .A(n445), .B(n444), .C(n443), .D(n442), .Y(n446) );
  AOI222XL U1079 ( .A0(n822), .A1(n93), .B0(n869), .B1(n81), .C0(n343), .C1(
        n286), .Y(n445) );
  AOI222XL U1080 ( .A0(lo_com[20]), .A1(n373), .B0(n287), .B1(n362), .C0(n288), 
        .C1(n333), .Y(n442) );
  NAND4X1 U1081 ( .A(n440), .B(n439), .C(n438), .D(n437), .Y(n441) );
  AOI222XL U1082 ( .A0(n822), .A1(n266), .B0(n869), .B1(n268), .C0(n343), .C1(
        n287), .Y(n440) );
  AOI222XL U1083 ( .A0(lo_com[19]), .A1(n373), .B0(n288), .B1(n362), .C0(n289), 
        .C1(n333), .Y(n437) );
  NAND4X1 U1084 ( .A(n455), .B(n454), .C(n453), .D(n452), .Y(n456) );
  AOI222XL U1085 ( .A0(n822), .A1(n261), .B0(n869), .B1(n263), .C0(n343), .C1(
        n292), .Y(n455) );
  NAND4X1 U1086 ( .A(n430), .B(n429), .C(n428), .D(n427), .Y(n431) );
  AOI222XL U1087 ( .A0(n822), .A1(n272), .B0(n869), .B1(n274), .C0(n343), .C1(
        n281), .Y(n430) );
  AOI222XL U1088 ( .A0(n824), .A1(n285), .B0(n287), .B1(n348), .C0(
        ALUinA_com[25]), .C1(n325), .Y(n429) );
  CLKMX2X2 U1089 ( .A(n516), .B(n282), .S0(n883), .Y(n1165) );
  NAND4X1 U1090 ( .A(n515), .B(n514), .C(n513), .D(n512), .Y(n516) );
  AOI222XL U1091 ( .A0(n822), .A1(n146), .B0(n869), .B1(n277), .C0(
        tempresult[2]), .C1(n345), .Y(n515) );
  AOI222XL U1092 ( .A0(n824), .A1(n281), .B0(n283), .B1(n347), .C0(
        ALUinA_com[29]), .C1(n326), .Y(n514) );
  MX2XL U1093 ( .A(n521), .B(n283), .S0(n375), .Y(n1166) );
  NAND4X1 U1094 ( .A(n520), .B(n519), .C(n518), .D(n517), .Y(n521) );
  AOI222XL U1095 ( .A0(n822), .A1(n275), .B0(n869), .B1(ALUinA[28]), .C0(
        tempresult[1]), .C1(n345), .Y(n520) );
  AOI222XL U1096 ( .A0(n824), .A1(n282), .B0(n284), .B1(n346), .C0(
        ALUinA_com[28]), .C1(n325), .Y(n519) );
  CLKMX2X2 U1097 ( .A(n526), .B(n288), .S0(n374), .Y(n1171) );
  NAND4X1 U1098 ( .A(n525), .B(n524), .C(n523), .D(n522), .Y(n526) );
  AOI222XL U1099 ( .A0(n822), .A1(n83), .B0(n869), .B1(n272), .C0(n345), .C1(
        n283), .Y(n525) );
  AOI222XL U1100 ( .A0(n824), .A1(n287), .B0(n289), .B1(n346), .C0(
        ALUinA_com[23]), .C1(n325), .Y(n524) );
  NAND4X1 U1101 ( .A(n530), .B(n529), .C(n528), .D(n527), .Y(n531) );
  AOI222XL U1102 ( .A0(n822), .A1(n85), .B0(n869), .B1(n267), .C0(n345), .C1(
        n288), .Y(n530) );
  AOI222XL U1103 ( .A0(n824), .A1(n292), .B0(n294), .B1(n346), .C0(
        ALUinA_com[18]), .C1(n325), .Y(n529) );
  NAND4X1 U1104 ( .A(n535), .B(n534), .C(n533), .D(n532), .Y(n536) );
  AOI222XL U1105 ( .A0(n822), .A1(n94), .B0(n869), .B1(n262), .C0(n345), .C1(
        n293), .Y(n535) );
  AOI222XL U1106 ( .A0(n824), .A1(n297), .B0(n299), .B1(n346), .C0(
        ALUinA_com[13]), .C1(n325), .Y(n534) );
  MX2XL U1107 ( .A(n541), .B(n303), .S0(n375), .Y(n1186) );
  NAND4X1 U1108 ( .A(n540), .B(n539), .C(n538), .D(n537), .Y(n541) );
  AOI222XL U1109 ( .A0(n822), .A1(n80), .B0(n869), .B1(n257), .C0(n345), .C1(
        n298), .Y(n540) );
  AOI222XL U1110 ( .A0(n328), .A1(n302), .B0(n304), .B1(n346), .C0(
        ALUinA_com[8]), .C1(n325), .Y(n539) );
  MX2XL U1111 ( .A(n466), .B(n295), .S0(n375), .Y(n1178) );
  NAND4X1 U1112 ( .A(n465), .B(n464), .C(n463), .D(n462), .Y(n466) );
  AOI222XL U1113 ( .A0(n822), .A1(n263), .B0(n869), .B1(n85), .C0(n343), .C1(
        n290), .Y(n465) );
  AOI222XL U1114 ( .A0(n824), .A1(n294), .B0(n296), .B1(n347), .C0(
        ALUinA_com[16]), .C1(n326), .Y(n464) );
  MX2XL U1115 ( .A(n461), .B(n296), .S0(n375), .Y(n1179) );
  NAND4X1 U1116 ( .A(n460), .B(n459), .C(n458), .D(n457), .Y(n461) );
  AOI222XL U1117 ( .A0(n822), .A1(n262), .B0(n869), .B1(n264), .C0(n343), .C1(
        n291), .Y(n460) );
  AOI222XL U1118 ( .A0(n824), .A1(n295), .B0(n297), .B1(n347), .C0(
        ALUinA_com[15]), .C1(n326), .Y(n459) );
  MX2XL U1119 ( .A(n481), .B(n300), .S0(n374), .Y(n1183) );
  NAND4X1 U1120 ( .A(n480), .B(n479), .C(n478), .D(n477), .Y(n481) );
  AOI222XL U1121 ( .A0(n822), .A1(n86), .B0(n869), .B1(n94), .C0(n343), .C1(
        n295), .Y(n480) );
  AOI222XL U1122 ( .A0(n824), .A1(n299), .B0(n301), .B1(n347), .C0(
        ALUinA_com[11]), .C1(n326), .Y(n479) );
  MX2XL U1123 ( .A(n476), .B(n301), .S0(n375), .Y(n1184) );
  NAND4X1 U1124 ( .A(n475), .B(n474), .C(n473), .D(n472), .Y(n476) );
  AOI222XL U1125 ( .A0(n822), .A1(n257), .B0(n869), .B1(n78), .C0(n343), .C1(
        n296), .Y(n475) );
  AOI222XL U1126 ( .A0(n824), .A1(n300), .B0(n302), .B1(n347), .C0(
        ALUinA_com[10]), .C1(n326), .Y(n474) );
  MX2XL U1127 ( .A(n471), .B(n302), .S0(n374), .Y(n1185) );
  NAND4X1 U1128 ( .A(n470), .B(n469), .C(n468), .D(n467), .Y(n471) );
  AOI222XL U1129 ( .A0(n822), .A1(n256), .B0(n869), .B1(n86), .C0(n343), .C1(
        n297), .Y(n470) );
  AOI222XL U1130 ( .A0(n824), .A1(n301), .B0(n303), .B1(n347), .C0(
        ALUinA_com[9]), .C1(n326), .Y(n469) );
  MX2XL U1131 ( .A(n496), .B(n305), .S0(n883), .Y(n1188) );
  NAND4X1 U1132 ( .A(n495), .B(n494), .C(n493), .D(n492), .Y(n496) );
  AOI222XL U1133 ( .A0(n822), .A1(n253), .B0(n869), .B1(n80), .C0(n345), .C1(
        n300), .Y(n495) );
  AOI222XL U1134 ( .A0(n824), .A1(n304), .B0(n306), .B1(n347), .C0(
        ALUinA_com[6]), .C1(n326), .Y(n494) );
  MX2XL U1135 ( .A(n801), .B(n284), .S0(n374), .Y(n1167) );
  NAND4X1 U1136 ( .A(n800), .B(n799), .C(n798), .D(n797), .Y(n801) );
  AOI222XL U1137 ( .A0(n822), .A1(n274), .B0(n869), .B1(n145), .C0(
        tempresult[0]), .C1(n345), .Y(n800) );
  AOI222XL U1138 ( .A0(n328), .A1(n283), .B0(n285), .B1(n347), .C0(
        ALUinA_com[27]), .C1(n325), .Y(n799) );
  NAND4X1 U1139 ( .A(n425), .B(n424), .C(n423), .D(n422), .Y(n426) );
  AOI222XL U1140 ( .A0(n822), .A1(n271), .B0(n869), .B1(n273), .C0(n343), .C1(
        n282), .Y(n425) );
  NAND4X1 U1141 ( .A(n805), .B(n804), .C(n803), .D(n802), .Y(n806) );
  AOI222XL U1142 ( .A0(n822), .A1(n81), .B0(n869), .B1(n271), .C0(n343), .C1(
        n284), .Y(n805) );
  AOI222XL U1143 ( .A0(n824), .A1(n288), .B0(n290), .B1(n346), .C0(
        ALUinA_com[22]), .C1(n325), .Y(n804) );
  NAND4X1 U1144 ( .A(n810), .B(n809), .C(n808), .D(n807), .Y(n811) );
  AOI222XL U1145 ( .A0(n822), .A1(n264), .B0(n869), .B1(n266), .C0(n343), .C1(
        n289), .Y(n810) );
  AOI222XL U1146 ( .A0(n824), .A1(n293), .B0(n295), .B1(n346), .C0(
        ALUinA_com[17]), .C1(n325), .Y(n809) );
  MX2XL U1147 ( .A(n816), .B(n299), .S0(n374), .Y(n1182) );
  NAND4X1 U1148 ( .A(n815), .B(n814), .C(n813), .D(n812), .Y(n816) );
  AOI222XL U1149 ( .A0(n822), .A1(n78), .B0(n869), .B1(n261), .C0(n343), .C1(
        n294), .Y(n815) );
  AOI222XL U1150 ( .A0(n824), .A1(n298), .B0(n300), .B1(n346), .C0(
        ALUinA_com[12]), .C1(n325), .Y(n814) );
  MX2XL U1151 ( .A(n821), .B(n304), .S0(n374), .Y(n1187) );
  NAND4X1 U1152 ( .A(n820), .B(n819), .C(n818), .D(n817), .Y(n821) );
  AOI222XL U1153 ( .A0(n822), .A1(n254), .B0(n869), .B1(n256), .C0(n343), .C1(
        n299), .Y(n820) );
  AOI222XL U1154 ( .A0(n824), .A1(n303), .B0(n305), .B1(n346), .C0(
        ALUinA_com[7]), .C1(n325), .Y(n819) );
  CLKINVX1 U1155 ( .A(n840), .Y(n843) );
  AO21XL U1156 ( .A0(n905), .A1(n206), .B0(n894), .Y(n875) );
  AO21X1 U1157 ( .A0(stateplus1[5]), .A1(n898), .B0(n863), .Y(state_next[5])
         );
  OAI221XL U1158 ( .A0(n862), .A1(n25), .B0(n1558), .B1(n861), .C0(n909), .Y(
        n863) );
  NOR4XL U1159 ( .A(n858), .B(n857), .C(n905), .D(n343), .Y(n861) );
  AOI222XL U1160 ( .A0(n897), .A1(n854), .B0(n894), .B1(n890), .C0(n892), .C1(
        n891), .Y(n862) );
  CLKINVX1 U1161 ( .A(n283), .Y(n1504) );
  CLKINVX1 U1162 ( .A(n285), .Y(n1482) );
  INVXL U1163 ( .A(n755), .Y(n415) );
  NAND3BX1 U1164 ( .AN(n908), .B(n420), .C(n1013), .Y(n558) );
  NAND2XL U1165 ( .A(n760), .B(n759), .Y(n794) );
  MX2XL U1166 ( .A(n973), .B(n991), .S0(n248), .Y(n759) );
  AOI2BB1XL U1167 ( .A0N(n203), .A1N(n844), .B0(n886), .Y(n848) );
  NAND2XL U1168 ( .A(n906), .B(n1129), .Y(n856) );
  AOI2BB1XL U1169 ( .A0N(n846), .A1N(n203), .B0(n845), .Y(n847) );
  CLKINVX1 U1170 ( .A(tempresult[0]), .Y(n563) );
  CLKINVX1 U1171 ( .A(n844), .Y(n853) );
  CLKINVX1 U1172 ( .A(n555), .Y(n1573) );
  NAND2BXL U1173 ( .AN(\halfresult[32] ), .B(n206), .Y(n555) );
  NAND2X1 U1174 ( .A(n760), .B(n758), .Y(n793) );
  MX2XL U1175 ( .A(n991), .B(n973), .S0(n248), .Y(n758) );
  CLKINVX1 U1176 ( .A(n281), .Y(n548) );
  OAI222XL U1177 ( .A0(n1505), .A1(n1251), .B0(n1507), .B1(n1256), .C0(n1503), 
        .C1(n1155), .Y(n1259) );
  CLKINVX1 U1178 ( .A(n304), .Y(n1251) );
  OAI222XL U1179 ( .A0(n1505), .A1(n1406), .B0(n1507), .B1(n1412), .C0(n1503), 
        .C1(n1141), .Y(n1415) );
  CLKINVX1 U1180 ( .A(n290), .Y(n1406) );
  AOI222X1 U1181 ( .A0(subaluinA[17]), .A1(n241), .B0(n158), .B1(n242), .C0(
        n294), .C1(n389), .Y(n1361) );
  AOI222X1 U1182 ( .A0(n67), .A1(n241), .B0(n160), .B1(n242), .C0(n300), .C1(
        n390), .Y(n1299) );
  AOI222X1 U1183 ( .A0(subaluinA[6]), .A1(n241), .B0(n184), .B1(n242), .C0(
        n305), .C1(n390), .Y(n1241) );
  AOI222X1 U1184 ( .A0(subaluinA[22]), .A1(n241), .B0(n15), .B1(n242), .C0(
        n289), .C1(n389), .Y(n1429) );
  AOI222X1 U1185 ( .A0(subaluinA[20]), .A1(n241), .B0(n185), .B1(n242), .C0(
        n291), .C1(n389), .Y(n1396) );
  AOI32XL U1186 ( .A0(n243), .A1(n262), .A2(n242), .B0(n298), .B1(n390), .Y(
        n1323) );
  AO22X1 U1187 ( .A0(reg_lo[0]), .A1(n191), .B0(n985), .B1(n943), .Y(n946) );
  OAI222XL U1188 ( .A0(n1505), .A1(n1013), .B0(n1507), .B1(n1018), .C0(n1503), 
        .C1(n1159), .Y(n1021) );
  NAND2X1 U1189 ( .A(n379), .B(n1438), .Y(n1441) );
  NAND2XL U1190 ( .A(n165), .B(n240), .Y(n1231) );
  OA22XL U1191 ( .A0(n1506), .A1(n1028), .B0(n1029), .B1(n381), .Y(n1135) );
  NAND2XL U1192 ( .A(n175), .B(n240), .Y(n1291) );
  NAND2X1 U1193 ( .A(n380), .B(n1289), .Y(n1292) );
  NAND2X1 U1194 ( .A(n380), .B(n1308), .Y(n1311) );
  BUFX20 U1195 ( .A(ALUinB[31]), .Y(n248) );
  BUFX20 U1196 ( .A(ALUinB[26]), .Y(n246) );
  NAND3BXL U1197 ( .AN(n976), .B(funct_regD[0]), .C(n178), .Y(n1535) );
  OAI221XL U1198 ( .A0(n1436), .A1(n321), .B0(n376), .B1(n34), .C0(n768), .Y(
        n1090) );
  NAND2X1 U1199 ( .A(ALUinB_com[23]), .B(n320), .Y(n768) );
  OAI221XL U1200 ( .A0(n214), .A1(n322), .B0(n377), .B1(n54), .C0(n780), .Y(
        n1078) );
  NAND2X1 U1201 ( .A(ALUinB_com[11]), .B(n791), .Y(n780) );
  OAI221XL U1202 ( .A0(n235), .A1(n322), .B0(n377), .B1(n35), .C0(n774), .Y(
        n1084) );
  OAI221XL U1203 ( .A0(n1347), .A1(n322), .B0(n377), .B1(n36), .C0(n775), .Y(
        n1083) );
  OAI221XL U1204 ( .A0(n132), .A1(n321), .B0(n376), .B1(n37), .C0(n772), .Y(
        n1086) );
  OAI221XL U1205 ( .A0(n1425), .A1(n321), .B0(n376), .B1(n38), .C0(n769), .Y(
        n1089) );
  OAI221XL U1206 ( .A0(n1521), .A1(n321), .B0(n376), .B1(n39), .C0(n762), .Y(
        n1096) );
  OAI221XL U1207 ( .A0(n1407), .A1(n321), .B0(n376), .B1(n40), .C0(n770), .Y(
        n1088) );
  OAI221XL U1208 ( .A0(n1532), .A1(n321), .B0(n376), .B1(n41), .C0(n761), .Y(
        n1097) );
  OAI221XL U1209 ( .A0(n1448), .A1(n321), .B0(n376), .B1(n32), .C0(n767), .Y(
        n1091) );
  OAI221XL U1210 ( .A0(n1306), .A1(n322), .B0(n377), .B1(n42), .C0(n779), .Y(
        n1079) );
  OAI221XL U1211 ( .A0(n114), .A1(n322), .B0(n377), .B1(n43), .C0(n776), .Y(
        n1082) );
  OAI221XL U1212 ( .A0(n1287), .A1(n322), .B0(n377), .B1(n44), .C0(n781), .Y(
        n1077) );
  NAND2XL U1213 ( .A(ALUOp_regD[2]), .B(n190), .Y(n980) );
  OAI221XL U1214 ( .A0(n1464), .A1(n321), .B0(n376), .B1(n45), .C0(n766), .Y(
        n1092) );
  OAI221XL U1215 ( .A0(n1315), .A1(n322), .B0(n377), .B1(n46), .C0(n778), .Y(
        n1080) );
  OAI221XL U1216 ( .A0(n1491), .A1(n321), .B0(n376), .B1(n55), .C0(n764), .Y(
        n1094) );
  NAND2XL U1217 ( .A(ALUinB_com[27]), .B(n320), .Y(n764) );
  OAI221XL U1218 ( .A0(n1392), .A1(n321), .B0(n376), .B1(n47), .C0(n771), .Y(
        n1087) );
  OAI221XL U1219 ( .A0(n1477), .A1(n321), .B0(n376), .B1(n53), .C0(n765), .Y(
        n1093) );
  OAI221XL U1220 ( .A0(n1508), .A1(n321), .B0(n376), .B1(n56), .C0(n763), .Y(
        n1095) );
  OAI221XL U1221 ( .A0(n1328), .A1(n322), .B0(n377), .B1(n57), .C0(n777), .Y(
        n1081) );
  OAI2BB2XL U1222 ( .B0(n757), .B1(n756), .A0N(n1066), .A1N(n865), .Y(n1098)
         );
  AOI32XL U1223 ( .A0(ALUinB_com[31]), .A1(n248), .A2(n991), .B0(n973), .B1(
        n754), .Y(n757) );
  CLKINVX1 U1224 ( .A(ALUinB_com[31]), .Y(n753) );
  MXI2X1 U1225 ( .A(n937), .B(n936), .S0(funct_regD[5]), .Y(n969) );
  NAND4BXL U1226 ( .AN(n935), .B(funct_regD[3]), .C(n976), .D(n933), .Y(n937)
         );
  NAND2XL U1227 ( .A(funct_regD[0]), .B(n934), .Y(n935) );
  NAND2XL U1228 ( .A(ALUOp_regD[0]), .B(n959), .Y(n960) );
  MX2XL U1229 ( .A(ALUOp_regD[0]), .B(n959), .S0(n958), .Y(n961) );
  INVXL U1230 ( .A(n908), .Y(n421) );
  NAND3BX1 U1231 ( .AN(n752), .B(n751), .C(n750), .Y(n1225) );
  OA22XL U1232 ( .A0(n1131), .A1(n748), .B0(n315), .B1(n747), .Y(n751) );
  AOI2BB2XL U1233 ( .B0(hi_com[31]), .B1(n319), .A0N(n738), .A1N(n95), .Y(n750) );
  OAI222XL U1234 ( .A0(n746), .A1(n745), .B0(n871), .B1(n744), .C0(n1131), 
        .C1(n743), .Y(n752) );
  AOI222XL U1235 ( .A0(lo_com[3]), .A1(n371), .B0(n304), .B1(n361), .C0(n305), 
        .C1(n331), .Y(n542) );
  AOI222XL U1236 ( .A0(lo_com[28]), .A1(n371), .B0(tempresult[0]), .B1(n361), 
        .C0(reg_lo[31]), .C1(n331), .Y(n517) );
  AOI222X1 U1237 ( .A0(lo_com[13]), .A1(n371), .B0(n294), .B1(n361), .C0(n295), 
        .C1(n331), .Y(n532) );
  AOI222X1 U1238 ( .A0(lo_com[7]), .A1(n371), .B0(n300), .B1(n361), .C0(n301), 
        .C1(n331), .Y(n817) );
  AOI222XL U1239 ( .A0(lo_com[2]), .A1(n371), .B0(n305), .B1(n361), .C0(n306), 
        .C1(n331), .Y(n826) );
  AOI222XL U1240 ( .A0(lo_com[29]), .A1(n372), .B0(tempresult[1]), .B1(n362), 
        .C0(tempresult[0]), .C1(n332), .Y(n512) );
  AOI222X1 U1241 ( .A0(lo_com[9]), .A1(n372), .B0(n298), .B1(n362), .C0(n299), 
        .C1(n332), .Y(n467) );
  AOI222X1 U1242 ( .A0(lo_com[6]), .A1(n372), .B0(n301), .B1(n362), .C0(n302), 
        .C1(n332), .Y(n492) );
  AOI222XL U1243 ( .A0(lo_com[5]), .A1(n372), .B0(n302), .B1(n362), .C0(n303), 
        .C1(n332), .Y(n487) );
  AOI222XL U1244 ( .A0(n306), .A1(n361), .B0(reg_lo[3]), .B1(n355), .C0(n351), 
        .C1(reg_lo[1]), .Y(n880) );
  AOI222XL U1245 ( .A0(n352), .A1(n282), .B0(ALUinA_com[27]), .B1(n329), .C0(
        reg_lo[31]), .C1(n355), .Y(n513) );
  AOI222XL U1246 ( .A0(n351), .A1(reg_lo[3]), .B0(n330), .B1(ALUinA_com[1]), 
        .C0(n306), .C1(n355), .Y(n543) );
  AOI222XL U1247 ( .A0(n352), .A1(reg_lo[4]), .B0(n330), .B1(ALUinA_com[2]), 
        .C0(n305), .C1(n356), .Y(n483) );
  AOI222XL U1248 ( .A0(n351), .A1(reg_lo[2]), .B0(ALUinA_com[0]), .B1(n330), 
        .C0(reg_lo[4]), .C1(n356), .Y(n827) );
  AOI222XL U1249 ( .A0(subaluinA[0]), .A1(n351), .B0(tempresult[1]), .B1(n824), 
        .C0(tempresult[2]), .C1(n355), .Y(n560) );
  OAI221XL U1250 ( .A0(n498), .A1(n558), .B0(n359), .B1(n1002), .C0(n497), .Y(
        n503) );
  CLKINVX1 U1251 ( .A(n306), .Y(n498) );
  AOI2BB2XL U1252 ( .B0(lo_com[0]), .B1(n373), .A0N(n368), .A1N(n877), .Y(n497) );
  OAI221XL U1253 ( .A0(n1275), .A1(n322), .B0(n377), .B1(n48), .C0(n782), .Y(
        n1076) );
  OAI221XL U1254 ( .A0(n217), .A1(n322), .B0(n377), .B1(n49), .C0(n783), .Y(
        n1075) );
  NAND2XL U1255 ( .A(ALUinB_com[8]), .B(n791), .Y(n783) );
  AOI2BB2XL U1256 ( .B0(lo_com[1]), .B1(n373), .A0N(n339), .A1N(n877), .Y(n879) );
  AND2XL U1257 ( .A(n1046), .B(n324), .Y(subaluinB[11]) );
  AND2XL U1258 ( .A(n1044), .B(n324), .Y(subaluinB[9]) );
  AND2XL U1259 ( .A(n1051), .B(n324), .Y(subaluinB[16]) );
  AND2XL U1260 ( .A(n1045), .B(n324), .Y(subaluinB[10]) );
  AND2XL U1261 ( .A(n1048), .B(n324), .Y(subaluinB[13]) );
  AND2XL U1262 ( .A(n1052), .B(n324), .Y(subaluinB[17]) );
  AND2XL U1263 ( .A(n1060), .B(n323), .Y(subaluinB[25]) );
  AND2XL U1264 ( .A(n1047), .B(n324), .Y(subaluinB[12]) );
  AND2XL U1265 ( .A(n1054), .B(n324), .Y(subaluinB[19]) );
  AND2XL U1266 ( .A(n1040), .B(n324), .Y(subaluinB[5]) );
  AND2XL U1267 ( .A(n1039), .B(n324), .Y(subaluinB[4]) );
  AND2XL U1268 ( .A(n1037), .B(n324), .Y(subaluinB[2]) );
  AND2XL U1269 ( .A(n1036), .B(n324), .Y(subaluinB[1]) );
  AND2XL U1270 ( .A(n1038), .B(n324), .Y(subaluinB[3]) );
  OAI2BB2XL U1271 ( .B0(n374), .B1(n506), .A0N(reg_lo[0]), .A1N(n505), .Y(
        n1191) );
  NAND2XL U1272 ( .A(n743), .B(n504), .Y(n505) );
  NOR4X1 U1273 ( .A(n503), .B(n502), .C(n501), .D(n500), .Y(n506) );
  AOI2BB1XL U1274 ( .A0N(n869), .A1N(n325), .B0(n918), .Y(n500) );
  NAND4BXL U1275 ( .AN(n947), .B(funct_regD[3]), .C(n991), .D(n967), .Y(n948)
         );
  NAND4X1 U1276 ( .A(n742), .B(n741), .C(n740), .D(n739), .Y(n1224) );
  OA22XL U1277 ( .A0(n747), .A1(n313), .B0(n314), .B1(n736), .Y(n741) );
  AOI222XL U1278 ( .A0(n735), .A1(subaluinA[30]), .B0(n734), .B1(subaluinA[29]), .C0(hi_com[30]), .C1(n319), .Y(n742) );
  AOI222XL U1279 ( .A0(ALUinA_com[30]), .A1(n329), .B0(n822), .B1(n278), .C0(
        tempresult[31]), .C1(n824), .Y(n740) );
  NAND4X1 U1280 ( .A(n733), .B(n732), .C(n731), .D(n730), .Y(n1223) );
  OA22XL U1281 ( .A0(n314), .A1(n728), .B0(n871), .B1(n747), .Y(n731) );
  AOI2BB2XL U1282 ( .B0(hi_com[29]), .B1(n319), .A0N(n313), .A1N(n736), .Y(
        n732) );
  OA22X1 U1283 ( .A0(n1133), .A1(n310), .B0(n1134), .B1(n95), .Y(n733) );
  AO22X1 U1284 ( .A0(n897), .A1(state[2]), .B0(n892), .B1(n853), .Y(n840) );
  NAND3XL U1285 ( .A(n867), .B(n866), .C(n865), .Y(state_next[0]) );
  MXI2XL U1286 ( .A(n892), .B(n864), .S0(\stateplus2[0] ), .Y(n866) );
  NAND2X1 U1287 ( .A(n898), .B(stateplus1[0]), .Y(n867) );
  OA22XL U1288 ( .A0(n359), .A1(n744), .B0(n738), .B1(n743), .Y(n739) );
  MX2XL U1289 ( .A(n554), .B(reg_lo[31]), .S0(n374), .Y(n1163) );
  OR4X1 U1290 ( .A(n553), .B(n552), .C(n551), .D(n550), .Y(n554) );
  OAI222XL U1291 ( .A0(n1522), .A1(n549), .B0(n558), .B1(n587), .C0(n349), 
        .C1(n548), .Y(n552) );
  OAI222XL U1292 ( .A0(n871), .A1(n563), .B0(n873), .B1(n745), .C0(n746), .C1(
        n547), .Y(n553) );
  MX2XL U1293 ( .A(n486), .B(reg_lo[4]), .S0(n883), .Y(n1190) );
  NAND4X1 U1294 ( .A(n485), .B(n484), .C(n483), .D(n482), .Y(n486) );
  AOI222XL U1295 ( .A0(n822), .A1(n251), .B0(n869), .B1(n88), .C0(n343), .C1(
        n302), .Y(n485) );
  AOI222XL U1296 ( .A0(n824), .A1(n306), .B0(reg_lo[3]), .B1(n347), .C0(
        ALUinA_com[4]), .C1(n326), .Y(n484) );
  MX2XL U1297 ( .A(n546), .B(reg_lo[3]), .S0(n374), .Y(n1222) );
  NAND4X1 U1298 ( .A(n545), .B(n544), .C(n543), .D(n542), .Y(n546) );
  AOI222XL U1299 ( .A0(n822), .A1(n250), .B0(n869), .B1(n89), .C0(n345), .C1(
        n303), .Y(n545) );
  AOI222XL U1300 ( .A0(n824), .A1(reg_lo[4]), .B0(reg_lo[2]), .B1(n346), .C0(
        ALUinA_com[3]), .C1(n325), .Y(n544) );
  MX2XL U1301 ( .A(n436), .B(n285), .S0(n375), .Y(n1168) );
  NAND4X1 U1302 ( .A(n435), .B(n434), .C(n433), .D(n432), .Y(n436) );
  AOI222XL U1303 ( .A0(n822), .A1(n273), .B0(n869), .B1(n275), .C0(n343), .C1(
        reg_lo[31]), .Y(n435) );
  AOI222XL U1304 ( .A0(lo_com[26]), .A1(n373), .B0(n281), .B1(n362), .C0(n282), 
        .C1(n333), .Y(n432) );
  MX2XL U1305 ( .A(n884), .B(reg_lo[1]), .S0(n883), .Y(n1192) );
  NAND4X1 U1306 ( .A(n882), .B(n881), .C(n880), .D(n879), .Y(n884) );
  AOI222XL U1307 ( .A0(reg_lo[0]), .A1(n346), .B0(n869), .B1(n250), .C0(n343), 
        .C1(n305), .Y(n882) );
  OA22XL U1308 ( .A0(n873), .A1(n872), .B0(n1002), .B1(n871), .Y(n881) );
  MX2XL U1309 ( .A(n830), .B(reg_lo[2]), .S0(n374), .Y(n1193) );
  NAND4X1 U1310 ( .A(n829), .B(n828), .C(n827), .D(n826), .Y(n830) );
  AOI222XL U1311 ( .A0(n822), .A1(n249), .B0(n869), .B1(n251), .C0(n343), .C1(
        n304), .Y(n829) );
  AOI222XL U1312 ( .A0(n824), .A1(reg_lo[3]), .B0(reg_lo[1]), .B1(n346), .C0(
        ALUinA_com[2]), .C1(n326), .Y(n828) );
  MX2XL U1313 ( .A(n511), .B(n281), .S0(n883), .Y(n1164) );
  NAND4X1 U1314 ( .A(n510), .B(n509), .C(n508), .D(n507), .Y(n511) );
  AOI222XL U1315 ( .A0(n822), .A1(n92), .B0(n869), .B1(n278), .C0(
        tempresult[3]), .C1(n345), .Y(n510) );
  AOI222XL U1316 ( .A0(n824), .A1(reg_lo[31]), .B0(n282), .B1(n347), .C0(
        ALUinA_com[30]), .C1(n326), .Y(n509) );
  MX2XL U1317 ( .A(n491), .B(n306), .S0(n883), .Y(n1189) );
  NAND4X1 U1318 ( .A(n490), .B(n489), .C(n488), .D(n487), .Y(n491) );
  AOI222XL U1319 ( .A0(n822), .A1(n89), .B0(n869), .B1(n82), .C0(n345), .C1(
        n301), .Y(n490) );
  AOI222XL U1320 ( .A0(n824), .A1(n305), .B0(reg_lo[4]), .B1(n347), .C0(
        ALUinA_com[5]), .C1(n326), .Y(n489) );
  AO22X1 U1321 ( .A0(lo_com[31]), .A1(n373), .B0(tempresult[2]), .B1(n333), 
        .Y(n551) );
  OAI2BB1X1 U1322 ( .A0N(stateplus1[4]), .A1N(n898), .B0(n851), .Y(
        state_next[4]) );
  MX2XL U1323 ( .A(n850), .B(n849), .S0(state[4]), .Y(n851) );
  AOI211XL U1324 ( .A0(n894), .A1(n852), .B0(n848), .C0(n847), .Y(n849) );
  OA22XL U1325 ( .A0(n843), .A1(n203), .B0(n852), .B1(n842), .Y(n850) );
  OAI2BB1X1 U1326 ( .A0N(stateplus1[1]), .A1N(n898), .B0(n889), .Y(
        state_next[1]) );
  MX2XL U1327 ( .A(n888), .B(n887), .S0(\stateplus4[1] ), .Y(n889) );
  AOI2BB1XL U1328 ( .A0N(n26), .A1N(n886), .B0(n897), .Y(n887) );
  INVX1 U1329 ( .A(n885), .Y(n888) );
  OAI2BB1X1 U1330 ( .A0N(stateplus1[3]), .A1N(n898), .B0(n839), .Y(
        state_next[3]) );
  MX2XL U1331 ( .A(n838), .B(n837), .S0(state[3]), .Y(n839) );
  AOI222XL U1332 ( .A0(n894), .A1(n19), .B0(n864), .B1(n846), .C0(n892), .C1(
        n844), .Y(n837) );
  AOI2BB1XL U1333 ( .A0N(n841), .A1N(n842), .B0(n840), .Y(n838) );
  AO21X1 U1334 ( .A0(stateplus1[2]), .A1(n898), .B0(n835), .Y(state_next[2])
         );
  MX2XL U1335 ( .A(n834), .B(n833), .S0(state[2]), .Y(n835) );
  OAI221XL U1336 ( .A0(n832), .A1(n886), .B0(n19), .B1(n842), .C0(n845), .Y(
        n834) );
  AND2XL U1337 ( .A(n885), .B(n19), .Y(n833) );
  OAI221XL U1338 ( .A0(n103), .A1(n322), .B0(n377), .B1(n50), .C0(n784), .Y(
        n1074) );
  OAI221XL U1339 ( .A0(n123), .A1(n321), .B0(n378), .B1(n22), .C0(n792), .Y(
        n1068) );
  NAND2X1 U1340 ( .A(ALUinB_com[1]), .B(n320), .Y(n792) );
  OAI221XL U1341 ( .A0(n127), .A1(n322), .B0(n378), .B1(n23), .C0(n790), .Y(
        n1069) );
  NAND2XL U1342 ( .A(ALUinB_com[2]), .B(n320), .Y(n790) );
  OAI221XL U1343 ( .A0(n405), .A1(n793), .B0(n378), .B1(n24), .C0(n789), .Y(
        n1070) );
  NAND2XL U1344 ( .A(ALUinB_com[3]), .B(n320), .Y(n789) );
  OAI221XL U1345 ( .A0(n101), .A1(n793), .B0(n378), .B1(n788), .C0(n787), .Y(
        n1071) );
  NAND2XL U1346 ( .A(ALUinB_com[4]), .B(n320), .Y(n787) );
  OAI221XL U1347 ( .A0(n117), .A1(n322), .B0(n378), .B1(n51), .C0(n786), .Y(
        n1072) );
  NAND2XL U1348 ( .A(ALUinB_com[5]), .B(n320), .Y(n786) );
  OAI221XL U1349 ( .A0(n135), .A1(n322), .B0(n378), .B1(n52), .C0(n785), .Y(
        n1073) );
  NAND2XL U1350 ( .A(ALUinB_com[6]), .B(n320), .Y(n785) );
  OR2X1 U1351 ( .A(n841), .B(n203), .Y(n852) );
  NAND3XL U1352 ( .A(state[4]), .B(state[3]), .C(n853), .Y(n891) );
  OR2X1 U1353 ( .A(n852), .B(n204), .Y(n890) );
  AND2XL U1354 ( .A(n1056), .B(n323), .Y(subaluinB[21]) );
  AND2XL U1355 ( .A(n1055), .B(n323), .Y(subaluinB[20]) );
  AND2XL U1356 ( .A(n1066), .B(n323), .Y(subaluinB[31]) );
  AND2XL U1357 ( .A(n1058), .B(n323), .Y(subaluinB[23]) );
  AND2XL U1358 ( .A(n1050), .B(n324), .Y(subaluinB[15]) );
  AND2XL U1359 ( .A(n1065), .B(n323), .Y(subaluinB[30]) );
  AND2XL U1360 ( .A(n1062), .B(n323), .Y(subaluinB[27]) );
  AND2XL U1361 ( .A(n1053), .B(n324), .Y(subaluinB[18]) );
  AND2XL U1362 ( .A(n1064), .B(n323), .Y(subaluinB[29]) );
  AND2XL U1363 ( .A(n1042), .B(n324), .Y(subaluinB[7]) );
  NAND2XL U1364 ( .A(\stateplus4[1] ), .B(state[2]), .Y(n841) );
  INVXL U1365 ( .A(reg_lo[31]), .Y(n556) );
  INVXL U1366 ( .A(reg_lo[4]), .Y(n877) );
  NOR2BX1 U1367 ( .AN(n373), .B(n206), .Y(n205) );
  AO22XL U1368 ( .A0(n400), .A1(n795), .B0(n1035), .B1(n865), .Y(n1067) );
  NAND2XL U1369 ( .A(n794), .B(n793), .Y(n795) );
  CLKINVX1 U1370 ( .A(n1138), .Y(n706) );
  CLKINVX1 U1371 ( .A(n1139), .Y(n700) );
  CLKINVX1 U1372 ( .A(n1140), .Y(n694) );
  CLKINVX1 U1373 ( .A(n1141), .Y(n688) );
  CLKINVX1 U1374 ( .A(n1142), .Y(n682) );
  CLKINVX1 U1375 ( .A(n1143), .Y(n676) );
  CLKINVX1 U1376 ( .A(n1144), .Y(n670) );
  CLKINVX1 U1377 ( .A(n1145), .Y(n664) );
  CLKINVX1 U1378 ( .A(n1146), .Y(n658) );
  CLKINVX1 U1379 ( .A(n1148), .Y(n646) );
  CLKINVX1 U1380 ( .A(n1149), .Y(n640) );
  CLKINVX1 U1381 ( .A(n1150), .Y(n634) );
  CLKINVX1 U1382 ( .A(n1152), .Y(n622) );
  CLKINVX1 U1383 ( .A(n1153), .Y(n616) );
  CLKINVX1 U1384 ( .A(n1154), .Y(n610) );
  CLKINVX1 U1385 ( .A(n1155), .Y(n604) );
  CLKINVX1 U1386 ( .A(n1156), .Y(n598) );
  CLKINVX1 U1387 ( .A(n1157), .Y(n592) );
  CLKINVX1 U1388 ( .A(n1158), .Y(n586) );
  CLKINVX1 U1389 ( .A(n1159), .Y(n580) );
  CLKINVX1 U1390 ( .A(n1160), .Y(n574) );
  CLKINVX1 U1391 ( .A(n1161), .Y(n568) );
  CLKINVX1 U1392 ( .A(n1134), .Y(n722) );
  INVXL U1393 ( .A(n209), .Y(n1306) );
  INVXL U1394 ( .A(n125), .Y(n1287) );
  INVXL U1395 ( .A(ALUinB[9]), .Y(n1275) );
  NAND2X1 U1396 ( .A(ALUinB[21]), .B(n83), .Y(n1412) );
  NAND4BX4 U1397 ( .AN(n966), .B(n965), .C(n964), .D(n963), .Y(ALUout[0]) );
  INVX8 U1398 ( .A(n1419), .Y(n1565) );
  INVX12 U1399 ( .A(n1416), .Y(n1564) );
  INVX8 U1400 ( .A(n1506), .Y(n1550) );
  INVX12 U1401 ( .A(n1566), .Y(n1354) );
  CLKBUFX20 U1402 ( .A(ALUOp_regD[4]), .Y(n280) );
  NAND2X2 U1403 ( .A(n26), .B(n19), .Y(n836) );
  NAND3BX2 U1404 ( .AN(funct_regD[2]), .B(funct_regD[4]), .C(n967), .Y(n414)
         );
  CLKINVX3 U1405 ( .A(n756), .Y(n760) );
  NAND2X2 U1406 ( .A(funct_regD[1]), .B(n975), .Y(n938) );
  NAND3BX2 U1407 ( .AN(n846), .B(state[4]), .C(state[3]), .Y(n854) );
  CLKINVX3 U1408 ( .A(n854), .Y(n896) );
  NAND2X2 U1409 ( .A(n896), .B(n25), .Y(n410) );
  CLKINVX3 U1410 ( .A(n836), .Y(n832) );
  NAND3BX2 U1411 ( .AN(n410), .B(n196), .C(n832), .Y(n908) );
  CLKINVX3 U1412 ( .A(reg_lo[2]), .Y(n1002) );
  CLKINVX3 U1413 ( .A(reg_lo[3]), .Y(n1013) );
  NAND2X2 U1414 ( .A(n418), .B(n908), .Y(n904) );
  NAND2X2 U1415 ( .A(n905), .B(state[6]), .Y(n499) );
  OAI31X2 U1416 ( .A0(n415), .A1(n414), .A2(n939), .B0(n198), .Y(n743) );
  NAND3BX2 U1417 ( .AN(reg_lo[1]), .B(n902), .C(n416), .Y(n842) );
  CLKINVX3 U1418 ( .A(n417), .Y(n878) );
  CLKINVX3 U1419 ( .A(n499), .Y(n860) );
  NAND2X2 U1420 ( .A(tempresult[31]), .B(n348), .Y(n749) );
  NAND2X2 U1421 ( .A(n760), .B(n755), .Y(n865) );
  NAND4X2 U1422 ( .A(n916), .B(n915), .C(n914), .D(n913), .Y(stall_muldiv) );
  CLKINVX3 U1423 ( .A(ALUOp_regD[5]), .Y(n920) );
  CLKINVX3 U1424 ( .A(ALUOp_regD[3]), .Y(n923) );
  NAND2X2 U1425 ( .A(n190), .B(n962), .Y(n982) );
  CLKINVX3 U1426 ( .A(n280), .Y(n1562) );
  AOI211X2 U1427 ( .A0(n928), .A1(n927), .B0(n983), .C0(n951), .Y(n966) );
  NAND4X2 U1428 ( .A(ALUOp_regD[2]), .B(n958), .C(n954), .D(n197), .Y(n1506)
         );
  NAND4X2 U1429 ( .A(n962), .B(n396), .C(n961), .D(n960), .Y(n1419) );
  NAND2X2 U1430 ( .A(N953), .B(n238), .Y(n963) );
  CLKINVX3 U1431 ( .A(n968), .Y(n992) );
  NAND2X2 U1432 ( .A(funct_regD[1]), .B(n992), .Y(n1416) );
  NAND2X2 U1433 ( .A(n984), .B(n969), .Y(n1566) );
  CLKINVX3 U1434 ( .A(n970), .Y(n971) );
  NAND2X2 U1435 ( .A(n191), .B(n984), .Y(n1505) );
  NAND2X2 U1436 ( .A(n178), .B(n991), .Y(n1507) );
  AOI211X2 U1437 ( .A0(N986), .A1(n239), .B0(n990), .C0(n989), .Y(n994) );
  NAND2X2 U1438 ( .A(N1050), .B(n170), .Y(n993) );
  AOI2BB1X2 U1439 ( .A0N(n392), .A1N(n998), .B0(n387), .Y(n999) );
  NAND4X2 U1440 ( .A(n1006), .B(n1005), .C(n1004), .D(n1003), .Y(n1007) );
  AOI221X2 U1441 ( .A0(N987), .A1(n239), .B0(N955), .B1(n1354), .C0(n1007), 
        .Y(n1009) );
  NAND2X2 U1442 ( .A(N1051), .B(n170), .Y(n1008) );
  OAI211X2 U1443 ( .A0(n1419), .A1(n1010), .B0(n1009), .C0(n1008), .Y(n1011)
         );
  NAND2X2 U1444 ( .A(N1084), .B(n1564), .Y(n1027) );
  CLKINVX3 U1445 ( .A(n1014), .Y(n1019) );
  OAI221X2 U1446 ( .A0(n1019), .A1(n1560), .B0(n1506), .B1(n1018), .C0(n1017), 
        .Y(n1020) );
  AOI211X2 U1447 ( .A0(N956), .A1(n1354), .B0(n1021), .C0(n1020), .Y(n1025) );
  NAND2X2 U1448 ( .A(N988), .B(n239), .Y(n1024) );
  NAND2X2 U1449 ( .A(N1052), .B(n170), .Y(n1022) );
  NAND4X2 U1450 ( .A(n1025), .B(n1024), .C(n1023), .D(n1022), .Y(n1026) );
  OA22X4 U1451 ( .A0(n1032), .A1(n1560), .B0(n1032), .B1(n1031), .Y(n1034) );
  NAND4X2 U1452 ( .A(n1135), .B(n1132), .C(n1034), .D(n1033), .Y(n1136) );
  AOI221X2 U1453 ( .A0(N957), .A1(n238), .B0(N989), .B1(n239), .C0(n1136), .Y(
        n1227) );
  NAND3BX2 U1454 ( .AN(n280), .B(N1053), .C(n170), .Y(n1151) );
  NAND2X2 U1455 ( .A(n1564), .B(n395), .Y(n1137) );
  NAND2X2 U1456 ( .A(N1085), .B(n1443), .Y(n1147) );
  NAND4X2 U1457 ( .A(n1233), .B(n1232), .C(n1231), .D(n1230), .Y(n1234) );
  AOI221X2 U1458 ( .A0(N958), .A1(n238), .B0(N958), .B1(n1354), .C0(n1234), 
        .Y(n1236) );
  NAND2X2 U1459 ( .A(N1086), .B(n1564), .Y(n1235) );
  NAND2X2 U1460 ( .A(N1087), .B(n1564), .Y(n1250) );
  CLKMX2X4 U1461 ( .A(n1239), .B(n382), .S0(n1238), .Y(n1244) );
  NAND2X2 U1462 ( .A(N991), .B(n239), .Y(n1247) );
  CLKINVX3 U1463 ( .A(N959), .Y(n1245) );
  AO22X4 U1464 ( .A0(N1056), .A1(n170), .B0(N992), .B1(n239), .Y(n1261) );
  OA21X4 U1465 ( .A0(n238), .A1(n1354), .B0(N960), .Y(n1260) );
  AOI2BB1X2 U1466 ( .A0N(n392), .A1N(n157), .B0(n387), .Y(n1264) );
  AOI2BB1X2 U1467 ( .A0N(n392), .A1N(n174), .B0(n387), .Y(n1276) );
  AND4X4 U1468 ( .A(n1281), .B(n1280), .C(n1279), .D(n1278), .Y(n1286) );
  OAI221X2 U1469 ( .A0(n280), .A1(n1286), .B0(n1285), .B1(n1284), .C0(n1283), 
        .Y(ALUout[9]) );
  AOI2BB1X2 U1470 ( .A0N(n392), .A1N(n175), .B0(n387), .Y(n1288) );
  NAND4X2 U1471 ( .A(n1293), .B(n1292), .C(n1291), .D(n1290), .Y(n1294) );
  NAND3BX2 U1472 ( .AN(n280), .B(n239), .C(N996), .Y(n1305) );
  NAND4X2 U1473 ( .A(n1312), .B(n1311), .C(n1310), .D(n1309), .Y(n1313) );
  NAND2BX2 U1474 ( .AN(n1317), .B(n1450), .Y(n1318) );
  NAND3BX2 U1475 ( .AN(n280), .B(n239), .C(N998), .Y(n1327) );
  CLKMX2X4 U1476 ( .A(n1330), .B(n382), .S0(n1329), .Y(n1335) );
  CLKMX2X4 U1477 ( .A(n1339), .B(n382), .S0(n1338), .Y(n1344) );
  AOI2BB1X2 U1478 ( .A0N(n392), .A1N(n156), .B0(n388), .Y(n1348) );
  NAND3BX2 U1479 ( .AN(n280), .B(n1564), .C(N1097), .Y(n1356) );
  NAND2X2 U1480 ( .A(n1354), .B(n395), .Y(n1417) );
  CLKMX2X4 U1481 ( .A(n1359), .B(n382), .S0(n1358), .Y(n1364) );
  NAND3BX2 U1482 ( .AN(n280), .B(N1066), .C(n170), .Y(n1366) );
  CLKMX2X4 U1483 ( .A(n1394), .B(n381), .S0(n1393), .Y(n1399) );
  NAND2X2 U1484 ( .A(N1101), .B(n1564), .Y(n1400) );
  NAND3BX2 U1485 ( .AN(n1566), .B(N973), .C(n395), .Y(n1404) );
  AOI32X2 U1486 ( .A0(N1069), .A1(n394), .A2(n170), .B0(N973), .B1(n238), .Y(
        n1403) );
  AOI2BB1X2 U1487 ( .A0N(n391), .A1N(n1409), .B0(n388), .Y(n1410) );
  AOI2BB1X2 U1488 ( .A0N(n1415), .A1N(n1414), .B0(n280), .Y(n1424) );
  NAND3BX2 U1489 ( .AN(n1416), .B(N1102), .C(n395), .Y(n1423) );
  AOI2BB1X2 U1490 ( .A0N(n391), .A1N(n15), .B0(n388), .Y(n1427) );
  AOI2BB1X2 U1491 ( .A0N(n391), .A1N(n180), .B0(n388), .Y(n1437) );
  AOI222X2 U1492 ( .A0(subaluinA[23]), .A1(n241), .B0(n180), .B1(n242), .C0(
        n288), .C1(n389), .Y(n1439) );
  NAND4X2 U1493 ( .A(n1442), .B(n1441), .C(n1440), .D(n1439), .Y(n1444) );
  AOI211X2 U1494 ( .A0(n379), .A1(n1455), .B0(n1454), .C0(n1453), .Y(n1456) );
  AOI221X2 U1495 ( .A0(N1073), .A1(n152), .B0(n1459), .B1(n394), .C0(n1458), 
        .Y(n1461) );
  AOI2BB1X2 U1496 ( .A0N(n392), .A1N(n1465), .B0(n388), .Y(n1468) );
  CLKMX2X4 U1497 ( .A(n1468), .B(n381), .S0(n1467), .Y(n1471) );
  AOI222X2 U1498 ( .A0(n63), .A1(n241), .B0(n1465), .B1(n242), .C0(n286), .C1(
        n389), .Y(n1469) );
  NAND4X2 U1499 ( .A(n1472), .B(n1471), .C(n1470), .D(n1469), .Y(n1473) );
  OAI221X2 U1500 ( .A0(N1106), .A1(n1473), .B0(n1564), .B1(n1473), .C0(n395), 
        .Y(n1474) );
  NAND2X4 U1501 ( .A(N1075), .B(n152), .Y(n1490) );
  AOI2BB1X2 U1502 ( .A0N(n391), .A1N(n1476), .B0(n388), .Y(n1479) );
  OAI221X2 U1503 ( .A0(N1107), .A1(n1487), .B0(n1564), .B1(n1487), .C0(n395), 
        .Y(n1489) );
  CLKMX2X4 U1504 ( .A(n1494), .B(n381), .S0(n1493), .Y(n1495) );
  OAI221X2 U1505 ( .A0(N1108), .A1(n1499), .B0(n1564), .B1(n1499), .C0(n395), 
        .Y(n1502) );
  AOI2BB1X2 U1506 ( .A0N(n391), .A1N(n1511), .B0(n388), .Y(n1512) );
  OAI221X2 U1507 ( .A0(N1109), .A1(n1517), .B0(n1564), .B1(n1517), .C0(n395), 
        .Y(n1519) );
  NAND2X4 U1508 ( .A(N1078), .B(n152), .Y(n1531) );
  AOI222X2 U1509 ( .A0(n186), .A1(n1534), .B0(n282), .B1(n389), .C0(
        subaluinA[29]), .C1(n241), .Y(n1526) );
  OAI211X2 U1510 ( .A0(n1539), .A1(n1560), .B0(n1538), .C0(n1537), .Y(n1540)
         );
  OAI221X2 U1511 ( .A0(N1111), .A1(n1540), .B0(n1564), .B1(n1540), .C0(n395), 
        .Y(n1545) );
  AOI22X4 U1512 ( .A0(N983), .A1(n1542), .B0(N1015), .B1(n1541), .Y(n1543) );
  OAI221X2 U1513 ( .A0(n1561), .A1(n1560), .B0(n391), .B1(n1558), .C0(n1557), 
        .Y(n1563) );
endmodule


module MIPS_Pipeline_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n38;

  CLKAND2X8 U1 ( .A(A[14]), .B(n24), .Y(n26) );
  AND2X2 U2 ( .A(A[11]), .B(n28), .Y(n27) );
  CLKXOR2X2 U3 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  INVX1 U4 ( .A(A[2]), .Y(SUM[2]) );
  CLKAND2X8 U5 ( .A(A[4]), .B(n9), .Y(n14) );
  XOR2X1 U6 ( .A(A[8]), .B(n16), .Y(SUM[8]) );
  CLKAND2X12 U7 ( .A(A[16]), .B(n23), .Y(n25) );
  CLKAND2X12 U8 ( .A(A[15]), .B(n26), .Y(n23) );
  CLKAND2X12 U9 ( .A(A[24]), .B(n10), .Y(n11) );
  CLKAND2X12 U10 ( .A(A[23]), .B(n13), .Y(n10) );
  CLKAND2X12 U11 ( .A(A[22]), .B(n18), .Y(n13) );
  CLKAND2X12 U12 ( .A(A[5]), .B(n14), .Y(n34) );
  CLKAND2X8 U13 ( .A(A[17]), .B(n25), .Y(n22) );
  NAND2X2 U14 ( .A(A[30]), .B(n15), .Y(n38) );
  CLKAND2X12 U15 ( .A(A[29]), .B(n32), .Y(n15) );
  CLKAND2X6 U16 ( .A(A[21]), .B(n20), .Y(n18) );
  CLKAND2X12 U17 ( .A(A[20]), .B(n19), .Y(n20) );
  CLKAND2X8 U18 ( .A(A[3]), .B(A[2]), .Y(n9) );
  CLKAND2X4 U19 ( .A(A[18]), .B(n22), .Y(n21) );
  XNOR2X2 U20 ( .A(A[31]), .B(n38), .Y(SUM[31]) );
  AND2X6 U21 ( .A(A[28]), .B(n17), .Y(n32) );
  AND2X8 U22 ( .A(A[9]), .B(n33), .Y(n31) );
  AND2X4 U23 ( .A(A[19]), .B(n21), .Y(n19) );
  AND2X8 U24 ( .A(A[26]), .B(n29), .Y(n12) );
  NAND2X2 U25 ( .A(A[28]), .B(n2), .Y(n3) );
  NAND2X1 U26 ( .A(n1), .B(n17), .Y(n4) );
  NAND2X4 U27 ( .A(n3), .B(n4), .Y(SUM[28]) );
  CLKINVX1 U28 ( .A(A[28]), .Y(n1) );
  CLKINVX1 U29 ( .A(n17), .Y(n2) );
  AND2X4 U30 ( .A(A[27]), .B(n12), .Y(n17) );
  NAND2X4 U31 ( .A(A[29]), .B(n6), .Y(n7) );
  NAND2X4 U32 ( .A(n5), .B(n32), .Y(n8) );
  NAND2X6 U33 ( .A(n7), .B(n8), .Y(SUM[29]) );
  CLKINVX1 U34 ( .A(A[29]), .Y(n5) );
  INVX2 U35 ( .A(n32), .Y(n6) );
  AND2X8 U36 ( .A(A[8]), .B(n16), .Y(n33) );
  AND2X8 U37 ( .A(A[7]), .B(n35), .Y(n16) );
  XOR2X4 U38 ( .A(A[30]), .B(n15), .Y(SUM[30]) );
  XOR2XL U39 ( .A(A[4]), .B(n9), .Y(SUM[4]) );
  AND2X4 U40 ( .A(A[6]), .B(n34), .Y(n35) );
  CLKXOR2X1 U41 ( .A(A[5]), .B(n14), .Y(SUM[5]) );
  CLKAND2X2 U42 ( .A(A[13]), .B(n30), .Y(n24) );
  AND2X2 U43 ( .A(A[10]), .B(n31), .Y(n28) );
  AND2X4 U44 ( .A(A[25]), .B(n11), .Y(n29) );
  XOR2X1 U45 ( .A(A[26]), .B(n29), .Y(SUM[26]) );
  XOR2X1 U46 ( .A(A[24]), .B(n10), .Y(SUM[24]) );
  XOR2X1 U47 ( .A(A[27]), .B(n12), .Y(SUM[27]) );
  XOR2X1 U48 ( .A(A[25]), .B(n11), .Y(SUM[25]) );
  AND2X2 U49 ( .A(A[12]), .B(n27), .Y(n30) );
  XOR2X1 U50 ( .A(A[22]), .B(n18), .Y(SUM[22]) );
  XOR2X1 U51 ( .A(A[20]), .B(n19), .Y(SUM[20]) );
  XOR2X1 U52 ( .A(A[18]), .B(n22), .Y(SUM[18]) );
  XOR2X1 U53 ( .A(A[23]), .B(n13), .Y(SUM[23]) );
  XOR2X1 U54 ( .A(A[21]), .B(n20), .Y(SUM[21]) );
  XOR2X1 U55 ( .A(A[19]), .B(n21), .Y(SUM[19]) );
  XOR2X1 U56 ( .A(A[17]), .B(n25), .Y(SUM[17]) );
  XOR2X1 U57 ( .A(A[15]), .B(n26), .Y(SUM[15]) );
  XOR2X1 U58 ( .A(A[16]), .B(n23), .Y(SUM[16]) );
  XOR2X1 U59 ( .A(A[10]), .B(n31), .Y(SUM[10]) );
  XOR2X1 U60 ( .A(A[11]), .B(n28), .Y(SUM[11]) );
  XOR2X1 U61 ( .A(A[13]), .B(n30), .Y(SUM[13]) );
  CLKXOR2X1 U62 ( .A(A[7]), .B(n35), .Y(SUM[7]) );
  XOR2X1 U63 ( .A(A[14]), .B(n24), .Y(SUM[14]) );
  CLKXOR2X1 U64 ( .A(A[9]), .B(n33), .Y(SUM[9]) );
  XOR2X1 U65 ( .A(A[12]), .B(n27), .Y(SUM[12]) );
  CLKXOR2X1 U66 ( .A(A[6]), .B(n34), .Y(SUM[6]) );
  CLKBUFX3 U67 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U68 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, flush, stallcache, stall_lw_use, JumpReg_m, MemRead_m,
         MemWrite_m, ALUsrc, RegWrite_m, Branch_DEC_m, MemRead_regD,
         MemWrite_regD, ALUsrc_regD, RegWrite_regD, JumpReg_regD, Branch_regD,
         RegWrite_regE, RegWrite_regM, Branch_DEC, MemRead, MemWrite, RegWrite,
         JumpReg, ExtOp, branchpred_his, pred_cond, stall_muldiv, predict,
         Jump_IF, Branch_IF, n16, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n149, n150, n161, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n201,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231;
  wire   [31:0] PCplus4;
  wire   [15:0] branchOffset_D;
  wire   [5:0] opcode;
  wire   [4:0] Rs;
  wire   [4:0] Rt;
  wire   [4:0] Rd;
  wire   [4:0] shamt;
  wire   [5:0] funct;
  wire   [15:0] immediate;
  wire   [31:0] PCplus4_regI;
  wire   [1:0] MemtoReg;
  wire   [5:0] ALUOp;
  wire   [5:0] funct_m;
  wire   [31:0] A_f;
  wire   [31:0] B_f;
  wire   [31:0] ExtOut;
  wire   [4:0] wsel;
  wire   [1:0] MemtoReg_regD;
  wire   [5:0] ALUOp_regD;
  wire   [5:0] funct_regD;
  wire   [31:0] A_regD;
  wire   [31:0] B_regD;
  wire   [31:0] ExtOut_regD;
  wire   [4:0] Rs_regD;
  wire   [4:0] Rt_regD;
  wire   [4:0] wsel_regD;
  wire   [31:0] PCplus4_regD;
  wire   [15:0] branchOffset_regD;
  wire   [31:0] tempALUinB;
  wire   [31:0] ALUout;
  wire   [1:0] MemtoReg_regE;
  wire   [4:0] wsel_regE;
  wire   [1:0] ALUout_regE;
  wire   [1:0] MemtoReg_regM;
  wire   [31:0] ALUout_regM;
  wire   [4:0] wsel_regM;
  wire   [31:0] dataOut_regM;
  wire   [1:0] RegDst;
  wire   [31:0] WriteData;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [1:0] FU_Asel;
  wire   [31:0] ALUinA;
  wire   [1:0] FU_Bsel;
  wire   [1:0] PCcur;
  wire   [2:0] PCsrc;
  wire   [31:0] PCnext;
  wire   [31:0] ALUinB;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;

  IF_DEC_regFile i_IF_DEC_regFile ( .clk(clk), .rst_n(ICACHE_ren), .flush(
        flush), .stallcache(n197), .stall_lw_use(stall_lw_use), 
        .instruction_next({n82, ICACHE_rdata[30:0]}), .PCplus4({PCplus4[31], 
        n132, n134, PCplus4[28], n133, PCplus4[26:5], n44, PCplus4[3:0]}), 
        .branchOffset(branchOffset_D), .opcode(opcode), .Rs(Rs), .Rt(Rt), .Rd(
        Rd), .shamt(shamt), .funct(funct), .immediate(immediate), 
        .PCplus4_regI(PCplus4_regI) );
  DEC_EX_regFile i_DEC_EX_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(n197), .MemtoReg(MemtoReg), .ALUOp(ALUOp), .JumpReg(
        JumpReg_m), .MemRead(MemRead_m), .MemWrite(MemWrite_m), .ALUsrc(ALUsrc), .RegWrite(RegWrite_m), .Branch(Branch_DEC_m), .PCplus4_regI(PCplus4_regI), 
        .funct(funct_m), .branchOffset_D(branchOffset_D), .A(A_f), .B(B_f), 
        .ExtOut(ExtOut), .Rs({n196, n195, n194, n193, n192}), .Rt({n191, n190, 
        n189, n188, n187}), .wsel(wsel), .MemtoReg_regD(MemtoReg_regD), 
        .ALUOp_regD(ALUOp_regD), .MemRead_regD(MemRead_regD), .MemWrite_regD(
        MemWrite_regD), .ALUsrc_regD(ALUsrc_regD), .RegWrite_regD(
        RegWrite_regD), .funct_regD(funct_regD), .A_regD(A_regD), .B_regD(
        B_regD), .ExtOut_regD(ExtOut_regD), .Rs_regD(Rs_regD), .Rt_regD(
        Rt_regD), .wsel_regD(wsel_regD), .JumpReg_regD(JumpReg_regD), 
        .Branch_regD(Branch_regD), .PCplus4_regD(PCplus4_regD), 
        .branchOffset_regD(branchOffset_regD) );
  EX_MEM_regFile i_EX_MEM_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(n197), .MemtoReg_regD(MemtoReg_regD), .MemRead_regD(
        MemRead_regD), .MemWrite_regD(MemWrite_regD), .RegWrite_regD(
        RegWrite_regD), .B_regD({tempALUinB[31:29], n131, n128, 
        tempALUinB[26:24], n130, tempALUinB[22:21], n97, tempALUinB[19:3], n41, 
        tempALUinB[1:0]}), .wsel_regD(wsel_regD), .ALUout({ALUout[31], n125, 
        ALUout[29:25], n109, ALUout[23:20], n90, ALUout[18:17], n121, 
        ALUout[15:14], n112, ALUout[12], n78, ALUout[10:7], n88, ALUout[5], 
        n63, ALUout[3], n126, ALUout[1], n89}), .MemtoReg_regE(MemtoReg_regE), 
        .MemRead_regE(DCACHE_ren), .MemWrite_regE(DCACHE_wen), .RegWrite_regE(
        RegWrite_regE), .B_regE(DCACHE_wdata), .wsel_regE(wsel_regE), 
        .ALUout_regE({DCACHE_addr[29], n232, n233, DCACHE_addr[26], n234, 
        DCACHE_addr[24:22], n235, n236, DCACHE_addr[19], n237, n238, n239, 
        n240, n241, n242, n243, n244, n245, DCACHE_addr[9], n246, n247, n248, 
        n249, n250, n251, n252, n253, n254, ALUout_regE}) );
  MEM_WB_regFile i_MEM_WB_regFile ( .clk(clk), .rst_n(ICACHE_ren), 
        .stallcache(n197), .MemtoReg_regE(MemtoReg_regE), .RegWrite_regE(
        RegWrite_regE), .ALUout_regE({DCACHE_addr, ALUout_regE}), .wsel_regE(
        wsel_regE), .dataOut({DCACHE_rdata[31:6], n43, DCACHE_rdata[4:0]}), 
        .MemtoReg_regM(MemtoReg_regM), .RegWrite_regM(RegWrite_regM), 
        .ALUout_regM(ALUout_regM), .wsel_regM(wsel_regM), .dataOut_regM(
        dataOut_regM) );
  maincontrol i_maincontrol ( .opcode(opcode), .funct(funct), .RegDst(RegDst), 
        .MemtoReg(MemtoReg), .ALUOp(ALUOp), .Branch(Branch_DEC), .MemRead(
        MemRead), .MemWrite(MemWrite), .ALUsrc(ALUsrc), .RegWrite(RegWrite), 
        .JumpReg(JumpReg), .ExtOp(ExtOp) );
  registerFile i_registrefFile ( .clk(clk), .rst_n(ICACHE_ren), .rsel1({n196, 
        n195, n194, n193, n192}), .rsel2({n191, n190, n189, n188, n187}), 
        .wsel({n127, n119, n116, n161, n123}), .wen(RegWrite_regM), .wdata({
        WriteData[31:21], n135, WriteData[19], n137, WriteData[17:2], n124, 
        n73}), .rdata1(A), .rdata2(B) );
  extender i_extender ( .shamt_i(shamt), .immed_i(immediate), .ExtOp_i(ExtOp), 
        .ExtOut_o(ExtOut) );
  MUX_5_3to1 MUX_wsel ( .data0_i({n191, n190, n189, n188, n187}), .data1_i(Rd), 
        .data2_i({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .select_i(RegDst), .data_o(
        wsel) );
  MUX_32_3to1_0 MUX_WriteData ( .data0_i(dataOut_regM), .data1_i({
        ALUout_regM[31:4], n58, ALUout_regM[2:0]}), .data2_i({
        ALUout_regM[31:4], n58, ALUout_regM[2:0]}), .select_i(MemtoReg_regM), 
        .data_o(WriteData) );
  MUX_32_3to1_2 MUX_ALUinA ( .data0_i(A_regD), .data1_i({WriteData[31:21], 
        n135, WriteData[19], n137, WriteData[17:2], n124, WriteData[0]}), 
        .data2_i({DCACHE_addr, ALUout_regE}), .select_i(FU_Asel), .data_o(
        ALUinA) );
  MUX_32_3to1_1 MUX_ALUinB ( .data0_i(B_regD), .data1_i({WriteData[31:21], 
        n135, WriteData[19], n137, WriteData[17:2], n124, WriteData[0]}), 
        .data2_i({DCACHE_addr, ALUout_regE}), .select_i(FU_Bsel), .data_o(
        tempALUinB) );
  forwarding i_forwarding ( .Rs_regD(Rs_regD), .Rt_regD(Rt_regD), 
        .RegWrite_regE(RegWrite_regE), .wsel_regE(wsel_regE), .RegWrite_regM(
        RegWrite_regM), .wsel_regM(wsel_regM), .FU_Asel(FU_Asel), .FU_Bsel(
        FU_Bsel) );
  hazard_detection i_hazard_detection ( .Branch_EX(Branch_regD), .equal(n143), 
        .branchpred_his(branchpred_his), .JumpReg_regD(JumpReg_regD), 
        .MemRead_regD(MemRead_regD), .Rt_regD({n92, Rt_regD[3:2], n101, n45}), 
        .Rs({n196, n195, n194, n193, n192}), .Rt({n191, n190, n189, n188, n187}), .ICACHE_stall(ICACHE_stall), .DCACHE_stall(DCACHE_stall), .stall_lw_use(
        stall_lw_use), .stallcache(stallcache), .flush(flush), .pred_cond(
        pred_cond), .stall_muldiv(stall_muldiv) );
  branch_prediction i_branch_prediction ( .clk(clk), .rst_n(ICACHE_ren), 
        .branch(Branch_regD), .equal(n231), .predict(predict), 
        .branchpred_his(branchpred_his) );
  precontrolDec i_precontrolDec ( .instruction_next(ICACHE_rdata), .Jump_IF(
        Jump_IF), .Branch_IF(Branch_IF) );
  nextPCcalculator i_nextPCcalculator ( .PCcur({ICACHE_addr, PCcur}), 
        .PCplus4({PCplus4[31], n132, n134, PCplus4[28], n133, PCplus4[26:5], 
        n44, PCplus4[3:0]}), .PCplus4_regD(PCplus4_regD), .targetAddr(
        ICACHE_rdata[25:0]), .branchOffset_I(ICACHE_rdata[15:0]), 
        .branchOffset_regD(branchOffset_regD), .JumpRegAddr({ALUinA[31:29], 
        n111, ALUinA[27], n118, ALUinA[25:24], n70, n77, ALUinA[21], n49, 
        ALUinA[19], n60, ALUinA[17:13], n39, n86, ALUinA[10], n57, n114, n47, 
        n72, n65, n62, n80, n68, ALUinA[1:0]}), .PCsrc(PCsrc), .PCnext(PCnext)
         );
  PCsrcLogic i_PCsrcLogic ( .pred_cond(pred_cond), .Branch_EX(Branch_regD), 
        .Branch_IF(Branch_IF), .equal(n231), .Jump(Jump_IF), .JumpReg(
        JumpReg_regD), .predict(predict), .stallcache(n197), .stall_lw_use(
        stall_lw_use), .PCsrc(PCsrc) );
  ALU i_ALU ( .clk(clk), .rst_n(ICACHE_ren), .ALUOp_regD(ALUOp_regD), 
        .funct_regD(funct_regD), .ALUinA(ALUinA), .ALUinB({ALUinB[31], n75, 
        ALUinB[29:22], n149, ALUinB[20:10], n150, ALUinB[8:7], n37, 
        ALUinB[5:2], n230, ALUinB[0]}), .ALUout(ALUout), .stall_muldiv(
        stall_muldiv) );
  MIPS_Pipeline_DW01_add_0 add_417 ( .A({ICACHE_addr, PCcur}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(PCplus4) );
  DFFRX4 \PCreg_reg[2]  ( .D(PCnext[2]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[0]) );
  DFFRX4 \PCreg_reg[3]  ( .D(PCnext[3]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[1]) );
  DFFRX4 \PCreg_reg[4]  ( .D(PCnext[4]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[2]) );
  DFFRX4 \PCreg_reg[29]  ( .D(PCnext[29]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[27]) );
  DFFRX4 \PCreg_reg[28]  ( .D(PCnext[28]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[26]) );
  DFFRX4 \PCreg_reg[22]  ( .D(PCnext[22]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[20]) );
  DFFRX4 \PCreg_reg[26]  ( .D(PCnext[26]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[24]) );
  DFFRX4 \PCreg_reg[25]  ( .D(PCnext[25]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[23]) );
  DFFRX4 \PCreg_reg[5]  ( .D(PCnext[5]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[3]) );
  DFFRX4 \PCreg_reg[6]  ( .D(PCnext[6]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[4]) );
  DFFRX4 \PCreg_reg[20]  ( .D(PCnext[20]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[18]) );
  DFFRX4 \PCreg_reg[24]  ( .D(PCnext[24]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[22]) );
  DFFRX4 \PCreg_reg[7]  ( .D(PCnext[7]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[5]) );
  DFFRX4 \PCreg_reg[9]  ( .D(PCnext[9]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[7]) );
  DFFRX2 \PCreg_reg[12]  ( .D(PCnext[12]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[10]) );
  DFFRX4 \PCreg_reg[8]  ( .D(PCnext[8]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[6]) );
  DFFRX2 \PCreg_reg[15]  ( .D(PCnext[15]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[13]) );
  DFFRX4 \PCreg_reg[19]  ( .D(PCnext[19]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[17]) );
  DFFRX2 \PCreg_reg[14]  ( .D(PCnext[14]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[12]) );
  DFFRX4 \PCreg_reg[30]  ( .D(PCnext[30]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[28]) );
  DFFRX4 \PCreg_reg[27]  ( .D(PCnext[27]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[25]) );
  DFFRX4 \PCreg_reg[31]  ( .D(PCnext[31]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[29]) );
  DFFRX4 \PCreg_reg[18]  ( .D(PCnext[18]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[16]) );
  DFFRX2 \PCreg_reg[11]  ( .D(PCnext[11]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[9]) );
  DFFRX2 \PCreg_reg[13]  ( .D(PCnext[13]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[11]) );
  DFFRX4 \PCreg_reg[0]  ( .D(PCnext[0]), .CK(clk), .RN(n203), .Q(PCcur[0]) );
  DFFRHQX2 \PCreg_reg[17]  ( .D(PCnext[17]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[15]) );
  DFFRHQX2 \PCreg_reg[16]  ( .D(PCnext[16]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[14]) );
  DFFRX2 \PCreg_reg[23]  ( .D(PCnext[23]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[21]) );
  DFFRX2 \PCreg_reg[21]  ( .D(PCnext[21]), .CK(clk), .RN(n203), .Q(
        ICACHE_addr[19]) );
  DFFRX4 \PCreg_reg[1]  ( .D(PCnext[1]), .CK(clk), .RN(ICACHE_ren), .Q(
        PCcur[1]) );
  DFFRX4 \PCreg_reg[10]  ( .D(PCnext[10]), .CK(clk), .RN(ICACHE_ren), .Q(
        ICACHE_addr[8]) );
  NOR3X6 U37 ( .A(ALUout[23]), .B(ALUout[3]), .C(ALUout[4]), .Y(n221) );
  INVX6 U38 ( .A(ALUout[16]), .Y(n120) );
  BUFX16 U39 ( .A(tempALUinB[27]), .Y(n128) );
  CLKMX2X6 U40 ( .A(tempALUinB[7]), .B(ExtOut_regD[7]), .S0(n36), .Y(ALUinB[7]) );
  CLKINVX20 U41 ( .A(n182), .Y(n36) );
  NAND2X6 U42 ( .A(tempALUinB[0]), .B(n182), .Y(n98) );
  CLKMX2X6 U43 ( .A(ExtOut_regD[6]), .B(tempALUinB[6]), .S0(ALUsrc_regD), .Y(
        n37) );
  INVXL U44 ( .A(ALUinA[12]), .Y(n38) );
  INVX1 U45 ( .A(n38), .Y(n39) );
  INVXL U46 ( .A(tempALUinB[2]), .Y(n40) );
  CLKINVX1 U47 ( .A(n40), .Y(n41) );
  NOR3X6 U48 ( .A(ALUout[20]), .B(ALUout[16]), .C(ALUout[24]), .Y(n218) );
  NAND3X8 U49 ( .A(n211), .B(n213), .C(n212), .Y(n214) );
  NOR2X8 U50 ( .A(ALUout[7]), .B(ALUout[22]), .Y(n211) );
  NOR2X8 U51 ( .A(n226), .B(n225), .Y(n227) );
  NOR2X8 U52 ( .A(ALUout[30]), .B(ALUout[9]), .Y(n219) );
  CLKINVX8 U53 ( .A(ALUout[0]), .Y(n206) );
  NAND2X8 U54 ( .A(n206), .B(n207), .Y(n216) );
  NOR4X8 U55 ( .A(n217), .B(n216), .C(n215), .D(n214), .Y(n228) );
  CLKINVX3 U56 ( .A(ExtOut_regD[5]), .Y(n50) );
  INVX16 U57 ( .A(n185), .Y(n183) );
  BUFX16 U58 ( .A(n252), .Y(DCACHE_addr[2]) );
  BUFX16 U59 ( .A(n251), .Y(DCACHE_addr[3]) );
  CLKINVX6 U60 ( .A(tempALUinB[23]), .Y(n129) );
  BUFX16 U61 ( .A(n186), .Y(n184) );
  INVX12 U62 ( .A(n93), .Y(n150) );
  INVX1 U63 ( .A(ExtOut_regD[9]), .Y(n94) );
  BUFX6 U64 ( .A(Rt[0]), .Y(n187) );
  CLKBUFX2 U65 ( .A(ALUout[30]), .Y(n125) );
  BUFX20 U66 ( .A(n201), .Y(ICACHE_ren) );
  BUFX2 U67 ( .A(n179), .Y(n178) );
  BUFX2 U68 ( .A(n179), .Y(n177) );
  INVX1 U69 ( .A(n170), .Y(n179) );
  BUFX2 U70 ( .A(n180), .Y(n175) );
  BUFX2 U71 ( .A(n180), .Y(n176) );
  CLKINVX3 U72 ( .A(n181), .Y(n173) );
  CLKINVX3 U73 ( .A(n181), .Y(n174) );
  INVX6 U74 ( .A(ALUsrc_regD), .Y(n186) );
  BUFX12 U75 ( .A(n186), .Y(n185) );
  CLKINVX12 U76 ( .A(n182), .Y(n55) );
  INVX1 U77 ( .A(n170), .Y(n180) );
  INVX8 U78 ( .A(n55), .Y(n95) );
  INVX1 U79 ( .A(n170), .Y(n181) );
  CLKBUFX3 U80 ( .A(PCplus4[4]), .Y(n44) );
  NOR2BX4 U81 ( .AN(n229), .B(stall_lw_use), .Y(n42) );
  INVX8 U82 ( .A(n66), .Y(n229) );
  AND2X1 U83 ( .A(Branch_DEC), .B(n42), .Y(Branch_DEC_m) );
  AND2X1 U84 ( .A(JumpReg), .B(n42), .Y(JumpReg_m) );
  AND2X1 U85 ( .A(MemRead), .B(n42), .Y(MemRead_m) );
  BUFX6 U86 ( .A(DCACHE_rdata[5]), .Y(n43) );
  CLKBUFX2 U87 ( .A(Rt_regD[0]), .Y(n45) );
  CLKMX2X6 U88 ( .A(ExtOut_regD[13]), .B(tempALUinB[13]), .S0(n182), .Y(
        ALUinB[13]) );
  NAND2X4 U89 ( .A(tempALUinB[8]), .B(n183), .Y(n52) );
  INVXL U90 ( .A(ALUinA[7]), .Y(n46) );
  CLKINVX1 U91 ( .A(n46), .Y(n47) );
  INVXL U92 ( .A(ALUinA[20]), .Y(n48) );
  INVX1 U93 ( .A(n48), .Y(n49) );
  OAI2BB2X4 U94 ( .B0(n50), .B1(n95), .A0N(tempALUinB[5]), .A1N(n95), .Y(
        ALUinB[5]) );
  NAND2X2 U95 ( .A(ExtOut_regD[8]), .B(n55), .Y(n51) );
  NAND2X8 U96 ( .A(n51), .B(n52), .Y(ALUinB[8]) );
  CLKAND2X3 U97 ( .A(n227), .B(n228), .Y(n231) );
  AND2X8 U98 ( .A(n227), .B(n228), .Y(n143) );
  NAND2X2 U99 ( .A(ExtOut_regD[15]), .B(n185), .Y(n53) );
  NAND2X6 U100 ( .A(tempALUinB[15]), .B(n183), .Y(n54) );
  NAND2X8 U101 ( .A(n53), .B(n54), .Y(ALUinB[15]) );
  MXI2X8 U102 ( .A(tempALUinB[21]), .B(ExtOut_regD[21]), .S0(n55), .Y(n145) );
  INVX4 U103 ( .A(n115), .Y(n116) );
  INVX4 U104 ( .A(ExtOut_regD[29]), .Y(n74) );
  BUFX8 U105 ( .A(n107), .Y(n119) );
  CLKMX2X4 U106 ( .A(ExtOut_regD[3]), .B(tempALUinB[3]), .S0(ALUsrc_regD), .Y(
        ALUinB[3]) );
  INVXL U107 ( .A(ALUinA[9]), .Y(n56) );
  CLKINVX1 U108 ( .A(n56), .Y(n57) );
  BUFX16 U109 ( .A(ALUout_regM[3]), .Y(n58) );
  INVXL U110 ( .A(ALUinA[18]), .Y(n59) );
  INVX1 U111 ( .A(n59), .Y(n60) );
  INVXL U112 ( .A(ALUinA[4]), .Y(n61) );
  INVX1 U113 ( .A(n61), .Y(n62) );
  CLKBUFX2 U114 ( .A(ALUout[4]), .Y(n63) );
  INVXL U115 ( .A(ALUinA[5]), .Y(n64) );
  CLKINVX1 U116 ( .A(n64), .Y(n65) );
  CLKBUFX2 U117 ( .A(flush), .Y(n66) );
  INVXL U118 ( .A(ALUinA[2]), .Y(n67) );
  CLKINVX1 U119 ( .A(n67), .Y(n68) );
  INVXL U120 ( .A(ALUinA[23]), .Y(n69) );
  INVX1 U121 ( .A(n69), .Y(n70) );
  CLKBUFX2 U122 ( .A(wsel_regM[1]), .Y(n161) );
  INVXL U123 ( .A(ALUinA[6]), .Y(n71) );
  CLKINVX1 U124 ( .A(n71), .Y(n72) );
  CLKBUFX2 U125 ( .A(wsel_regM[4]), .Y(n127) );
  CLKBUFX2 U126 ( .A(WriteData[0]), .Y(n73) );
  OAI2BB2X4 U127 ( .B0(n74), .B1(n95), .A0N(tempALUinB[29]), .A1N(n182), .Y(
        ALUinB[29]) );
  BUFX20 U128 ( .A(ALUinB[30]), .Y(n75) );
  INVXL U129 ( .A(ALUinA[22]), .Y(n76) );
  INVX1 U130 ( .A(n76), .Y(n77) );
  INVXL U131 ( .A(n209), .Y(n78) );
  INVXL U132 ( .A(ALUinA[3]), .Y(n79) );
  CLKINVX1 U133 ( .A(n79), .Y(n80) );
  INVXL U134 ( .A(ICACHE_rdata[31]), .Y(n81) );
  CLKINVX3 U135 ( .A(n81), .Y(n82) );
  INVXL U136 ( .A(ALUinA[11]), .Y(n85) );
  INVX1 U137 ( .A(n85), .Y(n86) );
  INVXL U138 ( .A(ALUout[24]), .Y(n108) );
  INVXL U139 ( .A(ALUout[6]), .Y(n87) );
  CLKINVX3 U140 ( .A(n87), .Y(n88) );
  INVXL U141 ( .A(n206), .Y(n89) );
  BUFX8 U142 ( .A(ALUout[19]), .Y(n90) );
  INVXL U143 ( .A(Rt_regD[4]), .Y(n91) );
  INVX1 U144 ( .A(n91), .Y(n92) );
  AOI2BB2X4 U145 ( .B0(tempALUinB[9]), .B1(n183), .A0N(n94), .A1N(n95), .Y(n93) );
  CLKBUFX20 U146 ( .A(n232), .Y(DCACHE_addr[28]) );
  INVXL U147 ( .A(tempALUinB[20]), .Y(n96) );
  CLKINVX1 U148 ( .A(n96), .Y(n97) );
  NAND3X6 U149 ( .A(n224), .B(n223), .C(n222), .Y(n225) );
  NAND2X8 U150 ( .A(ExtOut_regD[0]), .B(n185), .Y(n99) );
  NAND2X8 U151 ( .A(n98), .B(n99), .Y(ALUinB[0]) );
  CLKINVX20 U152 ( .A(n184), .Y(n182) );
  INVXL U153 ( .A(Rt_regD[1]), .Y(n100) );
  INVX3 U154 ( .A(n100), .Y(n101) );
  BUFX12 U155 ( .A(WriteData[20]), .Y(n135) );
  NAND2X2 U156 ( .A(ExtOut_regD[17]), .B(n185), .Y(n102) );
  NAND2X6 U157 ( .A(tempALUinB[17]), .B(n183), .Y(n103) );
  NAND2X8 U158 ( .A(n102), .B(n103), .Y(ALUinB[17]) );
  NOR2X8 U159 ( .A(ALUout[8]), .B(ALUout[18]), .Y(n208) );
  NAND2XL U160 ( .A(ExtOut_regD[19]), .B(n185), .Y(n104) );
  NAND2X8 U161 ( .A(tempALUinB[19]), .B(n183), .Y(n105) );
  NAND2X8 U162 ( .A(n104), .B(n105), .Y(ALUinB[19]) );
  INVXL U163 ( .A(wsel_regM[3]), .Y(n106) );
  INVX1 U164 ( .A(n106), .Y(n107) );
  INVX6 U165 ( .A(ALUout[2]), .Y(n212) );
  NAND2X6 U166 ( .A(tempALUinB[18]), .B(n182), .Y(n142) );
  CLKMX2X6 U167 ( .A(ExtOut_regD[20]), .B(tempALUinB[20]), .S0(n182), .Y(
        ALUinB[20]) );
  INVX1 U168 ( .A(ALUinA[26]), .Y(n117) );
  CLKINVX2 U169 ( .A(n108), .Y(n109) );
  INVXL U170 ( .A(ALUinA[28]), .Y(n110) );
  INVX1 U171 ( .A(n110), .Y(n111) );
  CLKBUFX2 U172 ( .A(ALUout[13]), .Y(n112) );
  INVXL U173 ( .A(ALUinA[8]), .Y(n113) );
  CLKINVX1 U174 ( .A(n113), .Y(n114) );
  INVXL U175 ( .A(wsel_regM[2]), .Y(n115) );
  INVX1 U176 ( .A(n117), .Y(n118) );
  INVX20 U177 ( .A(n145), .Y(n149) );
  CLKINVX8 U178 ( .A(ALUout[11]), .Y(n209) );
  CLKMX2X6 U179 ( .A(ExtOut_regD[28]), .B(n131), .S0(n182), .Y(ALUinB[28]) );
  INVX1 U180 ( .A(n120), .Y(n121) );
  INVXL U181 ( .A(wsel_regM[0]), .Y(n122) );
  INVX4 U182 ( .A(n122), .Y(n123) );
  BUFX16 U183 ( .A(WriteData[1]), .Y(n124) );
  NOR2BX4 U184 ( .AN(n229), .B(stall_lw_use), .Y(n144) );
  NOR2X8 U185 ( .A(ALUout[6]), .B(ALUout[1]), .Y(n213) );
  NOR4X8 U186 ( .A(n90), .B(ALUout[27]), .C(ALUout[29]), .D(ALUout[28]), .Y(
        n220) );
  NOR2X8 U187 ( .A(ALUout[31]), .B(ALUout[26]), .Y(n207) );
  NOR2X8 U188 ( .A(ALUout[13]), .B(ALUout[25]), .Y(n210) );
  INVXL U189 ( .A(n212), .Y(n126) );
  NAND4X6 U190 ( .A(n218), .B(n221), .C(n220), .D(n219), .Y(n226) );
  OR2X8 U191 ( .A(ALUout[21]), .B(ALUout[17]), .Y(n217) );
  NAND3X8 U192 ( .A(n208), .B(n210), .C(n209), .Y(n215) );
  NOR2X4 U193 ( .A(ALUout[15]), .B(ALUout[14]), .Y(n224) );
  NAND2X8 U194 ( .A(n130), .B(n183), .Y(n139) );
  NOR2X4 U195 ( .A(ALUout[12]), .B(ALUout[10]), .Y(n223) );
  BUFX20 U196 ( .A(stallcache), .Y(n197) );
  CLKBUFX20 U197 ( .A(n241), .Y(DCACHE_addr[14]) );
  CLKBUFX20 U198 ( .A(n248), .Y(DCACHE_addr[6]) );
  INVX8 U199 ( .A(ALUout[5]), .Y(n222) );
  BUFX16 U200 ( .A(PCplus4[29]), .Y(n134) );
  BUFX8 U201 ( .A(tempALUinB[28]), .Y(n131) );
  CLKMX2X4 U202 ( .A(ExtOut_regD[31]), .B(tempALUinB[31]), .S0(n182), .Y(
        ALUinB[31]) );
  CLKBUFX20 U203 ( .A(n246), .Y(DCACHE_addr[8]) );
  INVX8 U204 ( .A(n129), .Y(n130) );
  BUFX8 U205 ( .A(PCplus4[30]), .Y(n132) );
  BUFX6 U206 ( .A(PCplus4[27]), .Y(n133) );
  CLKINVX4 U207 ( .A(WriteData[18]), .Y(n136) );
  INVX6 U208 ( .A(n136), .Y(n137) );
  AO22X4 U209 ( .A0(ExtOut_regD[27]), .A1(n184), .B0(n128), .B1(n182), .Y(
        ALUinB[27]) );
  NAND2XL U210 ( .A(ExtOut_regD[23]), .B(n184), .Y(n138) );
  NAND2X8 U211 ( .A(n138), .B(n139), .Y(ALUinB[23]) );
  AND2X1 U212 ( .A(RegWrite), .B(n144), .Y(RegWrite_m) );
  AND2X1 U213 ( .A(MemWrite), .B(n144), .Y(MemWrite_m) );
  CLKBUFX4 U214 ( .A(n201), .Y(n203) );
  BUFX6 U215 ( .A(n16), .Y(n170) );
  INVXL U216 ( .A(n182), .Y(n146) );
  INVX3 U217 ( .A(n204), .Y(n205) );
  NAND2XL U218 ( .A(ExtOut_regD[1]), .B(n184), .Y(n204) );
  BUFX16 U219 ( .A(n250), .Y(DCACHE_addr[4]) );
  BUFX6 U220 ( .A(Rt[3]), .Y(n190) );
  BUFX6 U221 ( .A(Rt[2]), .Y(n189) );
  BUFX6 U222 ( .A(Rt[4]), .Y(n191) );
  BUFX6 U223 ( .A(Rs[3]), .Y(n195) );
  BUFX6 U224 ( .A(Rs[2]), .Y(n194) );
  BUFX16 U225 ( .A(Rt[1]), .Y(n188) );
  BUFX12 U226 ( .A(Rs[0]), .Y(n192) );
  BUFX12 U227 ( .A(Rs[1]), .Y(n193) );
  NAND2X2 U228 ( .A(ExtOut_regD[18]), .B(n140), .Y(n141) );
  NAND2X8 U229 ( .A(n141), .B(n142), .Y(ALUinB[18]) );
  INVXL U230 ( .A(n182), .Y(n140) );
  INVX3 U231 ( .A(n175), .Y(n171) );
  INVX3 U232 ( .A(n175), .Y(n172) );
  CLKBUFX3 U233 ( .A(rst_n), .Y(n201) );
  NOR2BX2 U234 ( .AN(MemtoReg[1]), .B(MemtoReg[0]), .Y(n16) );
  AOI2BB2X4 U235 ( .B0(n146), .B1(n204), .A0N(tempALUinB[1]), .A1N(n205), .Y(
        n230) );
  AND2XL U236 ( .A(funct[0]), .B(n229), .Y(funct_m[0]) );
  AND2XL U237 ( .A(funct[1]), .B(n229), .Y(funct_m[1]) );
  AND2XL U238 ( .A(funct[2]), .B(n229), .Y(funct_m[2]) );
  AND2XL U239 ( .A(funct[3]), .B(n229), .Y(funct_m[3]) );
  AND2XL U240 ( .A(funct[4]), .B(n229), .Y(funct_m[4]) );
  AND2XL U241 ( .A(funct[5]), .B(n229), .Y(funct_m[5]) );
  AO22X1 U242 ( .A0(B[0]), .A1(n176), .B0(PCplus4_regI[0]), .B1(n173), .Y(
        B_f[0]) );
  AO22X1 U243 ( .A0(B[1]), .A1(n177), .B0(PCplus4_regI[1]), .B1(n174), .Y(
        B_f[1]) );
  AO22X1 U244 ( .A0(B[2]), .A1(n178), .B0(PCplus4_regI[2]), .B1(n174), .Y(
        B_f[2]) );
  AO22X1 U245 ( .A0(B[3]), .A1(n176), .B0(PCplus4_regI[3]), .B1(n174), .Y(
        B_f[3]) );
  AO22X1 U246 ( .A0(B[4]), .A1(n176), .B0(PCplus4_regI[4]), .B1(n174), .Y(
        B_f[4]) );
  AO22X1 U247 ( .A0(B[5]), .A1(n176), .B0(PCplus4_regI[5]), .B1(n173), .Y(
        B_f[5]) );
  AO22X1 U248 ( .A0(B[6]), .A1(n176), .B0(PCplus4_regI[6]), .B1(n173), .Y(
        B_f[6]) );
  AO22X1 U249 ( .A0(B[7]), .A1(n179), .B0(PCplus4_regI[7]), .B1(n173), .Y(
        B_f[7]) );
  AO22X1 U250 ( .A0(B[8]), .A1(n178), .B0(PCplus4_regI[8]), .B1(n173), .Y(
        B_f[8]) );
  AO22X1 U251 ( .A0(B[9]), .A1(n177), .B0(PCplus4_regI[9]), .B1(n174), .Y(
        B_f[9]) );
  AO22X1 U252 ( .A0(B[10]), .A1(n178), .B0(PCplus4_regI[10]), .B1(n173), .Y(
        B_f[10]) );
  AO22X1 U253 ( .A0(B[11]), .A1(n177), .B0(PCplus4_regI[11]), .B1(n173), .Y(
        B_f[11]) );
  AO22X1 U254 ( .A0(B[12]), .A1(n175), .B0(PCplus4_regI[12]), .B1(n173), .Y(
        B_f[12]) );
  AO22X1 U255 ( .A0(B[13]), .A1(n176), .B0(PCplus4_regI[13]), .B1(n173), .Y(
        B_f[13]) );
  AO22X1 U256 ( .A0(B[14]), .A1(n176), .B0(PCplus4_regI[14]), .B1(n173), .Y(
        B_f[14]) );
  AO22X1 U257 ( .A0(B[15]), .A1(n176), .B0(PCplus4_regI[15]), .B1(n173), .Y(
        B_f[15]) );
  AO22X1 U258 ( .A0(B[16]), .A1(n176), .B0(PCplus4_regI[16]), .B1(n173), .Y(
        B_f[16]) );
  AO22X1 U259 ( .A0(B[17]), .A1(n176), .B0(PCplus4_regI[17]), .B1(n173), .Y(
        B_f[17]) );
  AO22X1 U260 ( .A0(B[18]), .A1(n176), .B0(PCplus4_regI[18]), .B1(n174), .Y(
        B_f[18]) );
  AO22X1 U261 ( .A0(B[19]), .A1(n176), .B0(PCplus4_regI[19]), .B1(n174), .Y(
        B_f[19]) );
  AO22X1 U262 ( .A0(B[20]), .A1(n177), .B0(PCplus4_regI[20]), .B1(n174), .Y(
        B_f[20]) );
  AO22X1 U263 ( .A0(B[21]), .A1(n177), .B0(PCplus4_regI[21]), .B1(n174), .Y(
        B_f[21]) );
  AO22X1 U264 ( .A0(B[22]), .A1(n177), .B0(PCplus4_regI[22]), .B1(n174), .Y(
        B_f[22]) );
  AO22X1 U265 ( .A0(B[23]), .A1(n177), .B0(PCplus4_regI[23]), .B1(n174), .Y(
        B_f[23]) );
  AO22X1 U266 ( .A0(B[24]), .A1(n177), .B0(PCplus4_regI[24]), .B1(n174), .Y(
        B_f[24]) );
  AO22X1 U267 ( .A0(B[25]), .A1(n178), .B0(PCplus4_regI[25]), .B1(n174), .Y(
        B_f[25]) );
  AO22X1 U268 ( .A0(B[26]), .A1(n178), .B0(PCplus4_regI[26]), .B1(n174), .Y(
        B_f[26]) );
  AO22X1 U269 ( .A0(B[27]), .A1(n178), .B0(PCplus4_regI[27]), .B1(n174), .Y(
        B_f[27]) );
  AO22X1 U270 ( .A0(B[28]), .A1(n178), .B0(PCplus4_regI[28]), .B1(n174), .Y(
        B_f[28]) );
  AO22X1 U271 ( .A0(B[29]), .A1(n178), .B0(PCplus4_regI[29]), .B1(n174), .Y(
        B_f[29]) );
  AO22X1 U272 ( .A0(B[30]), .A1(n176), .B0(PCplus4_regI[30]), .B1(n174), .Y(
        B_f[30]) );
  AO22X1 U273 ( .A0(B[31]), .A1(n176), .B0(PCplus4_regI[31]), .B1(n174), .Y(
        B_f[31]) );
  NOR2BX1 U274 ( .AN(A[0]), .B(n171), .Y(A_f[0]) );
  NOR2BX1 U275 ( .AN(A[1]), .B(n171), .Y(A_f[1]) );
  NOR2BX1 U276 ( .AN(A[2]), .B(n172), .Y(A_f[2]) );
  NOR2BX1 U277 ( .AN(A[3]), .B(n172), .Y(A_f[3]) );
  NOR2BX1 U278 ( .AN(A[4]), .B(n173), .Y(A_f[4]) );
  NOR2BX1 U279 ( .AN(A[5]), .B(n173), .Y(A_f[5]) );
  NOR2BX1 U280 ( .AN(A[6]), .B(n173), .Y(A_f[6]) );
  NOR2BX1 U281 ( .AN(A[7]), .B(n173), .Y(A_f[7]) );
  NOR2BX1 U282 ( .AN(A[8]), .B(n173), .Y(A_f[8]) );
  NOR2BX1 U283 ( .AN(A[9]), .B(n173), .Y(A_f[9]) );
  NOR2BX1 U284 ( .AN(A[10]), .B(n171), .Y(A_f[10]) );
  NOR2BX1 U285 ( .AN(A[11]), .B(n171), .Y(A_f[11]) );
  NOR2BX1 U286 ( .AN(A[12]), .B(n171), .Y(A_f[12]) );
  NOR2BX1 U287 ( .AN(A[13]), .B(n171), .Y(A_f[13]) );
  NOR2BX1 U288 ( .AN(A[14]), .B(n171), .Y(A_f[14]) );
  NOR2BX1 U289 ( .AN(A[15]), .B(n171), .Y(A_f[15]) );
  NOR2BX1 U290 ( .AN(A[16]), .B(n171), .Y(A_f[16]) );
  NOR2BX1 U291 ( .AN(A[17]), .B(n171), .Y(A_f[17]) );
  NOR2BX1 U292 ( .AN(A[18]), .B(n171), .Y(A_f[18]) );
  NOR2BX1 U293 ( .AN(A[19]), .B(n171), .Y(A_f[19]) );
  NOR2BX1 U294 ( .AN(A[20]), .B(n171), .Y(A_f[20]) );
  NOR2BX1 U295 ( .AN(A[21]), .B(n172), .Y(A_f[21]) );
  NOR2BX1 U296 ( .AN(A[22]), .B(n172), .Y(A_f[22]) );
  NOR2BX1 U297 ( .AN(A[23]), .B(n172), .Y(A_f[23]) );
  NOR2BX1 U298 ( .AN(A[24]), .B(n172), .Y(A_f[24]) );
  NOR2BX1 U299 ( .AN(A[25]), .B(n172), .Y(A_f[25]) );
  NOR2BX1 U300 ( .AN(A[26]), .B(n172), .Y(A_f[26]) );
  NOR2BX1 U301 ( .AN(A[27]), .B(n172), .Y(A_f[27]) );
  NOR2BX1 U302 ( .AN(A[28]), .B(n172), .Y(A_f[28]) );
  NOR2BX1 U303 ( .AN(A[29]), .B(n172), .Y(A_f[29]) );
  NOR2BX1 U304 ( .AN(A[30]), .B(n172), .Y(A_f[30]) );
  NOR2BX1 U305 ( .AN(A[31]), .B(n172), .Y(A_f[31]) );
  BUFX8 U306 ( .A(Rs[4]), .Y(n196) );
  BUFX20 U307 ( .A(n244), .Y(DCACHE_addr[11]) );
  BUFX20 U308 ( .A(n234), .Y(DCACHE_addr[25]) );
  BUFX20 U309 ( .A(n235), .Y(DCACHE_addr[21]) );
  BUFX20 U310 ( .A(n239), .Y(DCACHE_addr[16]) );
  BUFX20 U311 ( .A(n237), .Y(DCACHE_addr[18]) );
  BUFX20 U312 ( .A(n240), .Y(DCACHE_addr[15]) );
  BUFX20 U313 ( .A(n236), .Y(DCACHE_addr[20]) );
  BUFX20 U314 ( .A(n238), .Y(DCACHE_addr[17]) );
  BUFX20 U315 ( .A(n249), .Y(DCACHE_addr[5]) );
  BUFX20 U316 ( .A(n233), .Y(DCACHE_addr[27]) );
  BUFX20 U317 ( .A(n242), .Y(DCACHE_addr[13]) );
  BUFX20 U318 ( .A(n245), .Y(DCACHE_addr[10]) );
  BUFX20 U319 ( .A(n243), .Y(DCACHE_addr[12]) );
  BUFX20 U320 ( .A(n254), .Y(DCACHE_addr[0]) );
  BUFX20 U321 ( .A(n253), .Y(DCACHE_addr[1]) );
  BUFX20 U322 ( .A(n247), .Y(DCACHE_addr[7]) );
  AO22X4 U323 ( .A0(ExtOut_regD[2]), .A1(n55), .B0(tempALUinB[2]), .B1(n183), 
        .Y(ALUinB[2]) );
  AO22X4 U324 ( .A0(ExtOut_regD[4]), .A1(n55), .B0(tempALUinB[4]), .B1(n183), 
        .Y(ALUinB[4]) );
  AO22X4 U325 ( .A0(ExtOut_regD[10]), .A1(n185), .B0(tempALUinB[10]), .B1(n183), .Y(ALUinB[10]) );
  AO22X4 U326 ( .A0(ExtOut_regD[11]), .A1(n185), .B0(tempALUinB[11]), .B1(n183), .Y(ALUinB[11]) );
  AO22X4 U327 ( .A0(ExtOut_regD[12]), .A1(n185), .B0(tempALUinB[12]), .B1(n183), .Y(ALUinB[12]) );
  AO22X4 U328 ( .A0(ExtOut_regD[14]), .A1(n185), .B0(tempALUinB[14]), .B1(n183), .Y(ALUinB[14]) );
  AO22X4 U329 ( .A0(ExtOut_regD[16]), .A1(n185), .B0(tempALUinB[16]), .B1(n183), .Y(ALUinB[16]) );
  AO22X4 U330 ( .A0(ExtOut_regD[22]), .A1(n185), .B0(tempALUinB[22]), .B1(n183), .Y(ALUinB[22]) );
  CLKMX2X4 U331 ( .A(ExtOut_regD[24]), .B(tempALUinB[24]), .S0(n182), .Y(
        ALUinB[24]) );
  CLKMX2X4 U332 ( .A(ExtOut_regD[25]), .B(tempALUinB[25]), .S0(n182), .Y(
        ALUinB[25]) );
  AO22X4 U333 ( .A0(ExtOut_regD[26]), .A1(n184), .B0(tempALUinB[26]), .B1(n183), .Y(ALUinB[26]) );
  AO22X4 U334 ( .A0(ExtOut_regD[30]), .A1(n185), .B0(tempALUinB[30]), .B1(n183), .Y(ALUinB[30]) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         \blocktag[7][21] , \blocktag[7][20] , \blocktag[7][18] ,
         \blocktag[7][17] , \blocktag[7][16] , \blocktag[7][15] ,
         \blocktag[7][13] , \blocktag[7][11] , \blocktag[7][9] ,
         \blocktag[7][8] , \blocktag[7][7] , \blocktag[7][6] ,
         \blocktag[7][5] , \blocktag[7][2] , \blocktag[7][1] ,
         \blocktag[7][0] , \blocktag[6][21] , \blocktag[6][20] ,
         \blocktag[6][18] , \blocktag[6][17] , \blocktag[6][16] ,
         \blocktag[6][15] , \blocktag[6][13] , \blocktag[6][11] ,
         \blocktag[6][9] , \blocktag[6][8] , \blocktag[6][7] ,
         \blocktag[6][6] , \blocktag[6][5] , \blocktag[6][2] ,
         \blocktag[6][1] , \blocktag[6][0] , \blocktag[5][21] ,
         \blocktag[5][20] , \blocktag[5][18] , \blocktag[5][17] ,
         \blocktag[5][16] , \blocktag[5][15] , \blocktag[5][13] ,
         \blocktag[5][11] , \blocktag[5][9] , \blocktag[5][8] ,
         \blocktag[5][7] , \blocktag[5][6] , \blocktag[5][5] ,
         \blocktag[5][2] , \blocktag[5][1] , \blocktag[5][0] ,
         \blocktag[4][21] , \blocktag[4][20] , \blocktag[4][18] ,
         \blocktag[4][17] , \blocktag[4][16] , \blocktag[4][15] ,
         \blocktag[4][13] , \blocktag[4][11] , \blocktag[4][9] ,
         \blocktag[4][8] , \blocktag[4][7] , \blocktag[4][6] ,
         \blocktag[4][5] , \blocktag[4][2] , \blocktag[4][1] ,
         \blocktag[4][0] , \blocktag[3][21] , \blocktag[3][20] ,
         \blocktag[3][18] , \blocktag[3][17] , \blocktag[3][16] ,
         \blocktag[3][15] , \blocktag[3][13] , \blocktag[3][11] ,
         \blocktag[3][9] , \blocktag[3][8] , \blocktag[3][7] ,
         \blocktag[3][6] , \blocktag[3][5] , \blocktag[3][2] ,
         \blocktag[3][1] , \blocktag[3][0] , \blocktag[2][21] ,
         \blocktag[2][20] , \blocktag[2][18] , \blocktag[2][17] ,
         \blocktag[2][16] , \blocktag[2][15] , \blocktag[2][13] ,
         \blocktag[2][11] , \blocktag[2][9] , \blocktag[2][8] ,
         \blocktag[2][7] , \blocktag[2][6] , \blocktag[2][5] ,
         \blocktag[2][2] , \blocktag[2][1] , \blocktag[2][0] ,
         \blocktag[1][21] , \blocktag[1][20] , \blocktag[1][18] ,
         \blocktag[1][17] , \blocktag[1][16] , \blocktag[1][15] ,
         \blocktag[1][13] , \blocktag[1][11] , \blocktag[1][9] ,
         \blocktag[1][8] , \blocktag[1][7] , \blocktag[1][6] ,
         \blocktag[1][5] , \blocktag[1][2] , \blocktag[1][1] ,
         \blocktag[1][0] , \blocktag[0][21] , \blocktag[0][20] ,
         \blocktag[0][18] , \blocktag[0][17] , \blocktag[0][16] ,
         \blocktag[0][15] , \blocktag[0][13] , \blocktag[0][11] ,
         \blocktag[0][9] , \blocktag[0][8] , \blocktag[0][7] ,
         \blocktag[0][6] , \blocktag[0][5] , \blocktag[0][2] ,
         \blocktag[0][1] , \blocktag[0][0] , valid, dirty, \block[7][127] ,
         \block[7][126] , \block[7][125] , \block[7][124] , \block[7][123] ,
         \block[7][122] , \block[7][121] , \block[7][120] , \block[7][119] ,
         \block[7][118] , \block[7][117] , \block[7][116] , \block[7][115] ,
         \block[7][114] , \block[7][113] , \block[7][112] , \block[7][111] ,
         \block[7][110] , \block[7][109] , \block[7][108] , \block[7][107] ,
         \block[7][106] , \block[7][105] , \block[7][104] , \block[7][103] ,
         \block[7][102] , \block[7][101] , \block[7][100] , \block[7][99] ,
         \block[7][98] , \block[7][97] , \block[7][96] , \block[7][95] ,
         \block[7][94] , \block[7][93] , \block[7][92] , \block[7][91] ,
         \block[7][90] , \block[7][89] , \block[7][88] , \block[7][87] ,
         \block[7][86] , \block[7][85] , \block[7][84] , \block[7][83] ,
         \block[7][82] , \block[7][81] , \block[7][80] , \block[7][79] ,
         \block[7][78] , \block[7][77] , \block[7][76] , \block[7][75] ,
         \block[7][74] , \block[7][73] , \block[7][72] , \block[7][71] ,
         \block[7][70] , \block[7][69] , \block[7][68] , \block[7][67] ,
         \block[7][66] , \block[7][65] , \block[7][64] , \block[7][63] ,
         \block[7][62] , \block[7][61] , \block[7][60] , \block[7][59] ,
         \block[7][58] , \block[7][57] , \block[7][56] , \block[7][55] ,
         \block[7][54] , \block[7][53] , \block[7][52] , \block[7][51] ,
         \block[7][50] , \block[7][49] , \block[7][48] , \block[7][47] ,
         \block[7][46] , \block[7][45] , \block[7][44] , \block[7][43] ,
         \block[7][42] , \block[7][41] , \block[7][40] , \block[7][39] ,
         \block[7][38] , \block[7][37] , \block[7][36] , \block[7][35] ,
         \block[7][34] , \block[7][33] , \block[7][32] , \block[7][31] ,
         \block[7][30] , \block[7][29] , \block[7][28] , \block[7][27] ,
         \block[7][26] , \block[7][25] , \block[7][24] , \block[7][23] ,
         \block[7][22] , \block[7][21] , \block[7][20] , \block[7][19] ,
         \block[7][18] , \block[7][17] , \block[7][16] , \block[7][15] ,
         \block[7][14] , \block[7][13] , \block[7][12] , \block[7][11] ,
         \block[7][10] , \block[7][9] , \block[7][8] , \block[7][7] ,
         \block[7][6] , \block[7][5] , \block[7][4] , \block[7][3] ,
         \block[7][2] , \block[7][1] , \block[7][0] , \block[6][127] ,
         \block[6][126] , \block[6][125] , \block[6][124] , \block[6][123] ,
         \block[6][122] , \block[6][121] , \block[6][120] , \block[6][119] ,
         \block[6][118] , \block[6][117] , \block[6][116] , \block[6][115] ,
         \block[6][114] , \block[6][113] , \block[6][112] , \block[6][111] ,
         \block[6][110] , \block[6][109] , \block[6][108] , \block[6][107] ,
         \block[6][106] , \block[6][105] , \block[6][104] , \block[6][103] ,
         \block[6][102] , \block[6][101] , \block[6][100] , \block[6][99] ,
         \block[6][98] , \block[6][97] , \block[6][96] , \block[6][95] ,
         \block[6][94] , \block[6][93] , \block[6][92] , \block[6][91] ,
         \block[6][90] , \block[6][89] , \block[6][88] , \block[6][87] ,
         \block[6][86] , \block[6][85] , \block[6][84] , \block[6][83] ,
         \block[6][82] , \block[6][81] , \block[6][80] , \block[6][79] ,
         \block[6][78] , \block[6][77] , \block[6][76] , \block[6][75] ,
         \block[6][74] , \block[6][73] , \block[6][72] , \block[6][71] ,
         \block[6][70] , \block[6][69] , \block[6][68] , \block[6][67] ,
         \block[6][66] , \block[6][65] , \block[6][64] , \block[6][63] ,
         \block[6][62] , \block[6][61] , \block[6][60] , \block[6][59] ,
         \block[6][58] , \block[6][57] , \block[6][56] , \block[6][55] ,
         \block[6][54] , \block[6][53] , \block[6][52] , \block[6][51] ,
         \block[6][50] , \block[6][49] , \block[6][48] , \block[6][47] ,
         \block[6][46] , \block[6][45] , \block[6][44] , \block[6][43] ,
         \block[6][42] , \block[6][41] , \block[6][40] , \block[6][39] ,
         \block[6][38] , \block[6][37] , \block[6][36] , \block[6][35] ,
         \block[6][34] , \block[6][33] , \block[6][32] , \block[6][31] ,
         \block[6][30] , \block[6][29] , \block[6][28] , \block[6][27] ,
         \block[6][26] , \block[6][25] , \block[6][24] , \block[6][23] ,
         \block[6][22] , \block[6][21] , \block[6][20] , \block[6][19] ,
         \block[6][18] , \block[6][17] , \block[6][16] , \block[6][15] ,
         \block[6][14] , \block[6][13] , \block[6][12] , \block[6][11] ,
         \block[6][10] , \block[6][9] , \block[6][8] , \block[6][7] ,
         \block[6][6] , \block[6][5] , \block[6][4] , \block[6][3] ,
         \block[6][2] , \block[6][1] , \block[6][0] , \block[5][127] ,
         \block[5][126] , \block[5][125] , \block[5][124] , \block[5][123] ,
         \block[5][122] , \block[5][121] , \block[5][120] , \block[5][119] ,
         \block[5][118] , \block[5][117] , \block[5][116] , \block[5][115] ,
         \block[5][114] , \block[5][113] , \block[5][112] , \block[5][111] ,
         \block[5][110] , \block[5][109] , \block[5][108] , \block[5][107] ,
         \block[5][106] , \block[5][105] , \block[5][104] , \block[5][103] ,
         \block[5][102] , \block[5][101] , \block[5][100] , \block[5][99] ,
         \block[5][98] , \block[5][97] , \block[5][96] , \block[5][95] ,
         \block[5][94] , \block[5][93] , \block[5][92] , \block[5][91] ,
         \block[5][90] , \block[5][89] , \block[5][88] , \block[5][87] ,
         \block[5][86] , \block[5][85] , \block[5][84] , \block[5][83] ,
         \block[5][82] , \block[5][81] , \block[5][80] , \block[5][79] ,
         \block[5][78] , \block[5][77] , \block[5][76] , \block[5][75] ,
         \block[5][74] , \block[5][73] , \block[5][72] , \block[5][71] ,
         \block[5][70] , \block[5][69] , \block[5][68] , \block[5][67] ,
         \block[5][66] , \block[5][65] , \block[5][64] , \block[5][63] ,
         \block[5][62] , \block[5][61] , \block[5][60] , \block[5][59] ,
         \block[5][58] , \block[5][57] , \block[5][56] , \block[5][55] ,
         \block[5][54] , \block[5][53] , \block[5][52] , \block[5][51] ,
         \block[5][50] , \block[5][49] , \block[5][48] , \block[5][47] ,
         \block[5][46] , \block[5][45] , \block[5][44] , \block[5][43] ,
         \block[5][42] , \block[5][41] , \block[5][40] , \block[5][39] ,
         \block[5][38] , \block[5][37] , \block[5][36] , \block[5][35] ,
         \block[5][34] , \block[5][33] , \block[5][32] , \block[5][31] ,
         \block[5][30] , \block[5][29] , \block[5][28] , \block[5][27] ,
         \block[5][26] , \block[5][25] , \block[5][24] , \block[5][23] ,
         \block[5][22] , \block[5][21] , \block[5][20] , \block[5][19] ,
         \block[5][18] , \block[5][17] , \block[5][16] , \block[5][15] ,
         \block[5][14] , \block[5][13] , \block[5][12] , \block[5][11] ,
         \block[5][10] , \block[5][9] , \block[5][8] , \block[5][7] ,
         \block[5][6] , \block[5][5] , \block[5][4] , \block[5][3] ,
         \block[5][2] , \block[5][1] , \block[5][0] , \block[4][127] ,
         \block[4][126] , \block[4][125] , \block[4][124] , \block[4][123] ,
         \block[4][122] , \block[4][121] , \block[4][120] , \block[4][119] ,
         \block[4][118] , \block[4][117] , \block[4][116] , \block[4][115] ,
         \block[4][114] , \block[4][113] , \block[4][112] , \block[4][111] ,
         \block[4][110] , \block[4][109] , \block[4][108] , \block[4][107] ,
         \block[4][106] , \block[4][105] , \block[4][104] , \block[4][103] ,
         \block[4][102] , \block[4][101] , \block[4][100] , \block[4][99] ,
         \block[4][98] , \block[4][97] , \block[4][96] , \block[4][95] ,
         \block[4][94] , \block[4][93] , \block[4][92] , \block[4][91] ,
         \block[4][90] , \block[4][89] , \block[4][88] , \block[4][87] ,
         \block[4][86] , \block[4][85] , \block[4][84] , \block[4][83] ,
         \block[4][82] , \block[4][81] , \block[4][80] , \block[4][79] ,
         \block[4][78] , \block[4][77] , \block[4][76] , \block[4][75] ,
         \block[4][74] , \block[4][73] , \block[4][72] , \block[4][71] ,
         \block[4][70] , \block[4][69] , \block[4][68] , \block[4][67] ,
         \block[4][66] , \block[4][65] , \block[4][64] , \block[4][63] ,
         \block[4][62] , \block[4][61] , \block[4][60] , \block[4][59] ,
         \block[4][58] , \block[4][57] , \block[4][56] , \block[4][55] ,
         \block[4][54] , \block[4][53] , \block[4][52] , \block[4][51] ,
         \block[4][50] , \block[4][49] , \block[4][48] , \block[4][47] ,
         \block[4][46] , \block[4][45] , \block[4][44] , \block[4][43] ,
         \block[4][42] , \block[4][41] , \block[4][40] , \block[4][39] ,
         \block[4][38] , \block[4][37] , \block[4][36] , \block[4][35] ,
         \block[4][34] , \block[4][33] , \block[4][32] , \block[4][31] ,
         \block[4][30] , \block[4][29] , \block[4][28] , \block[4][27] ,
         \block[4][26] , \block[4][25] , \block[4][24] , \block[4][23] ,
         \block[4][22] , \block[4][21] , \block[4][20] , \block[4][19] ,
         \block[4][18] , \block[4][17] , \block[4][16] , \block[4][15] ,
         \block[4][14] , \block[4][13] , \block[4][12] , \block[4][11] ,
         \block[4][10] , \block[4][9] , \block[4][8] , \block[4][7] ,
         \block[4][6] , \block[4][5] , \block[4][4] , \block[4][3] ,
         \block[4][2] , \block[4][1] , \block[4][0] , \block[3][127] ,
         \block[3][126] , \block[3][125] , \block[3][124] , \block[3][123] ,
         \block[3][122] , \block[3][121] , \block[3][120] , \block[3][119] ,
         \block[3][118] , \block[3][117] , \block[3][116] , \block[3][115] ,
         \block[3][114] , \block[3][113] , \block[3][112] , \block[3][111] ,
         \block[3][110] , \block[3][109] , \block[3][108] , \block[3][107] ,
         \block[3][106] , \block[3][105] , \block[3][104] , \block[3][103] ,
         \block[3][102] , \block[3][101] , \block[3][100] , \block[3][99] ,
         \block[3][98] , \block[3][97] , \block[3][96] , \block[3][95] ,
         \block[3][94] , \block[3][93] , \block[3][92] , \block[3][91] ,
         \block[3][90] , \block[3][89] , \block[3][88] , \block[3][87] ,
         \block[3][86] , \block[3][85] , \block[3][84] , \block[3][83] ,
         \block[3][82] , \block[3][81] , \block[3][80] , \block[3][79] ,
         \block[3][78] , \block[3][77] , \block[3][76] , \block[3][75] ,
         \block[3][74] , \block[3][73] , \block[3][72] , \block[3][71] ,
         \block[3][70] , \block[3][69] , \block[3][68] , \block[3][67] ,
         \block[3][66] , \block[3][65] , \block[3][64] , \block[3][63] ,
         \block[3][62] , \block[3][61] , \block[3][60] , \block[3][59] ,
         \block[3][58] , \block[3][57] , \block[3][56] , \block[3][55] ,
         \block[3][54] , \block[3][53] , \block[3][52] , \block[3][51] ,
         \block[3][50] , \block[3][49] , \block[3][48] , \block[3][47] ,
         \block[3][46] , \block[3][45] , \block[3][44] , \block[3][43] ,
         \block[3][42] , \block[3][41] , \block[3][40] , \block[3][39] ,
         \block[3][38] , \block[3][37] , \block[3][36] , \block[3][35] ,
         \block[3][34] , \block[3][33] , \block[3][32] , \block[3][31] ,
         \block[3][30] , \block[3][29] , \block[3][28] , \block[3][27] ,
         \block[3][26] , \block[3][25] , \block[3][24] , \block[3][23] ,
         \block[3][22] , \block[3][21] , \block[3][20] , \block[3][19] ,
         \block[3][18] , \block[3][17] , \block[3][16] , \block[3][15] ,
         \block[3][14] , \block[3][13] , \block[3][12] , \block[3][11] ,
         \block[3][10] , \block[3][9] , \block[3][8] , \block[3][7] ,
         \block[3][6] , \block[3][4] , \block[3][3] , \block[3][2] ,
         \block[3][1] , \block[3][0] , \block[2][127] , \block[2][126] ,
         \block[2][125] , \block[2][124] , \block[2][123] , \block[2][122] ,
         \block[2][121] , \block[2][120] , \block[2][119] , \block[2][118] ,
         \block[2][117] , \block[2][116] , \block[2][115] , \block[2][114] ,
         \block[2][113] , \block[2][112] , \block[2][111] , \block[2][110] ,
         \block[2][109] , \block[2][108] , \block[2][107] , \block[2][106] ,
         \block[2][105] , \block[2][104] , \block[2][103] , \block[2][102] ,
         \block[2][101] , \block[2][100] , \block[2][99] , \block[2][98] ,
         \block[2][97] , \block[2][96] , \block[2][95] , \block[2][94] ,
         \block[2][93] , \block[2][92] , \block[2][91] , \block[2][90] ,
         \block[2][89] , \block[2][88] , \block[2][87] , \block[2][86] ,
         \block[2][85] , \block[2][84] , \block[2][83] , \block[2][82] ,
         \block[2][81] , \block[2][80] , \block[2][79] , \block[2][78] ,
         \block[2][77] , \block[2][76] , \block[2][75] , \block[2][74] ,
         \block[2][73] , \block[2][72] , \block[2][71] , \block[2][70] ,
         \block[2][69] , \block[2][68] , \block[2][67] , \block[2][66] ,
         \block[2][65] , \block[2][64] , \block[2][63] , \block[2][62] ,
         \block[2][61] , \block[2][60] , \block[2][59] , \block[2][58] ,
         \block[2][57] , \block[2][56] , \block[2][55] , \block[2][54] ,
         \block[2][53] , \block[2][52] , \block[2][51] , \block[2][50] ,
         \block[2][49] , \block[2][48] , \block[2][47] , \block[2][46] ,
         \block[2][45] , \block[2][44] , \block[2][43] , \block[2][42] ,
         \block[2][41] , \block[2][40] , \block[2][39] , \block[2][38] ,
         \block[2][37] , \block[2][36] , \block[2][35] , \block[2][34] ,
         \block[2][33] , \block[2][32] , \block[2][31] , \block[2][30] ,
         \block[2][29] , \block[2][28] , \block[2][27] , \block[2][26] ,
         \block[2][25] , \block[2][24] , \block[2][23] , \block[2][22] ,
         \block[2][21] , \block[2][20] , \block[2][19] , \block[2][18] ,
         \block[2][17] , \block[2][16] , \block[2][15] , \block[2][14] ,
         \block[2][13] , \block[2][12] , \block[2][11] , \block[2][10] ,
         \block[2][9] , \block[2][8] , \block[2][7] , \block[2][6] ,
         \block[2][4] , \block[2][3] , \block[2][2] , \block[2][1] ,
         \block[2][0] , \block[1][127] , \block[1][126] , \block[1][125] ,
         \block[1][124] , \block[1][123] , \block[1][122] , \block[1][121] ,
         \block[1][120] , \block[1][119] , \block[1][118] , \block[1][117] ,
         \block[1][116] , \block[1][115] , \block[1][114] , \block[1][113] ,
         \block[1][112] , \block[1][111] , \block[1][110] , \block[1][109] ,
         \block[1][108] , \block[1][107] , \block[1][106] , \block[1][105] ,
         \block[1][104] , \block[1][103] , \block[1][102] , \block[1][101] ,
         \block[1][100] , \block[1][99] , \block[1][98] , \block[1][97] ,
         \block[1][96] , \block[1][95] , \block[1][94] , \block[1][93] ,
         \block[1][92] , \block[1][91] , \block[1][90] , \block[1][89] ,
         \block[1][88] , \block[1][87] , \block[1][86] , \block[1][85] ,
         \block[1][84] , \block[1][83] , \block[1][82] , \block[1][81] ,
         \block[1][80] , \block[1][79] , \block[1][78] , \block[1][77] ,
         \block[1][76] , \block[1][75] , \block[1][74] , \block[1][73] ,
         \block[1][72] , \block[1][71] , \block[1][70] , \block[1][69] ,
         \block[1][68] , \block[1][67] , \block[1][66] , \block[1][65] ,
         \block[1][64] , \block[1][63] , \block[1][62] , \block[1][61] ,
         \block[1][60] , \block[1][59] , \block[1][58] , \block[1][57] ,
         \block[1][56] , \block[1][55] , \block[1][54] , \block[1][53] ,
         \block[1][52] , \block[1][51] , \block[1][50] , \block[1][49] ,
         \block[1][48] , \block[1][47] , \block[1][46] , \block[1][45] ,
         \block[1][44] , \block[1][43] , \block[1][42] , \block[1][41] ,
         \block[1][40] , \block[1][39] , \block[1][38] , \block[1][37] ,
         \block[1][36] , \block[1][35] , \block[1][34] , \block[1][33] ,
         \block[1][32] , \block[1][31] , \block[1][30] , \block[1][29] ,
         \block[1][28] , \block[1][27] , \block[1][26] , \block[1][25] ,
         \block[1][24] , \block[1][23] , \block[1][22] , \block[1][21] ,
         \block[1][20] , \block[1][19] , \block[1][18] , \block[1][17] ,
         \block[1][16] , \block[1][15] , \block[1][14] , \block[1][13] ,
         \block[1][12] , \block[1][11] , \block[1][10] , \block[1][9] ,
         \block[1][8] , \block[1][7] , \block[1][6] , \block[1][4] ,
         \block[1][3] , \block[1][2] , \block[1][1] , \block[1][0] ,
         \block[0][127] , \block[0][126] , \block[0][125] , \block[0][124] ,
         \block[0][123] , \block[0][122] , \block[0][121] , \block[0][120] ,
         \block[0][119] , \block[0][118] , \block[0][117] , \block[0][116] ,
         \block[0][115] , \block[0][114] , \block[0][113] , \block[0][112] ,
         \block[0][111] , \block[0][110] , \block[0][109] , \block[0][108] ,
         \block[0][107] , \block[0][106] , \block[0][105] , \block[0][104] ,
         \block[0][103] , \block[0][102] , \block[0][101] , \block[0][100] ,
         \block[0][99] , \block[0][98] , \block[0][97] , \block[0][96] ,
         \block[0][95] , \block[0][94] , \block[0][93] , \block[0][92] ,
         \block[0][91] , \block[0][90] , \block[0][89] , \block[0][88] ,
         \block[0][87] , \block[0][86] , \block[0][85] , \block[0][84] ,
         \block[0][83] , \block[0][82] , \block[0][81] , \block[0][80] ,
         \block[0][79] , \block[0][78] , \block[0][77] , \block[0][76] ,
         \block[0][75] , \block[0][74] , \block[0][73] , \block[0][72] ,
         \block[0][71] , \block[0][70] , \block[0][69] , \block[0][68] ,
         \block[0][67] , \block[0][66] , \block[0][65] , \block[0][64] ,
         \block[0][63] , \block[0][62] , \block[0][61] , \block[0][60] ,
         \block[0][59] , \block[0][58] , \block[0][57] , \block[0][56] ,
         \block[0][55] , \block[0][54] , \block[0][53] , \block[0][52] ,
         \block[0][51] , \block[0][50] , \block[0][49] , \block[0][48] ,
         \block[0][47] , \block[0][46] , \block[0][45] , \block[0][44] ,
         \block[0][43] , \block[0][42] , \block[0][41] , \block[0][40] ,
         \block[0][39] , \block[0][38] , \block[0][37] , \block[0][36] ,
         \block[0][35] , \block[0][34] , \block[0][33] , \block[0][32] ,
         \block[0][31] , \block[0][30] , \block[0][29] , \block[0][28] ,
         \block[0][27] , \block[0][26] , \block[0][25] , \block[0][24] ,
         \block[0][23] , \block[0][22] , \block[0][21] , \block[0][20] ,
         \block[0][19] , \block[0][18] , \block[0][17] , \block[0][16] ,
         \block[0][15] , \block[0][14] , \block[0][13] , \block[0][12] ,
         \block[0][11] , \block[0][10] , \block[0][9] , \block[0][8] ,
         \block[0][7] , \block[0][6] , \block[0][4] , \block[0][3] ,
         \block[0][2] , \block[0][1] , \block[0][0] , n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n503, n1, n2, n3, n5, n7, n9, n11, n13,
         n15, n17, n19, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39, n41,
         n43, n45, n47, n49, n51, n53, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n502, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n788, n789, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  EDFFXL \block_reg[7][116]  ( .D(block_next[116]), .E(n651), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFXL \block_reg[7][115]  ( .D(block_next[115]), .E(n651), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFXL \block_reg[7][114]  ( .D(block_next[114]), .E(n651), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFXL \block_reg[7][113]  ( .D(block_next[113]), .E(n651), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFXL \block_reg[7][112]  ( .D(block_next[112]), .E(n651), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFXL \block_reg[7][111]  ( .D(block_next[111]), .E(n651), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFXL \block_reg[7][110]  ( .D(block_next[110]), .E(n651), .CK(clk), .Q(
        \block[7][110] ) );
  EDFFXL \block_reg[7][109]  ( .D(block_next[109]), .E(n651), .CK(clk), .Q(
        \block[7][109] ) );
  EDFFXL \block_reg[7][108]  ( .D(block_next[108]), .E(n651), .CK(clk), .Q(
        \block[7][108] ) );
  EDFFXL \block_reg[7][107]  ( .D(block_next[107]), .E(n651), .CK(clk), .Q(
        \block[7][107] ) );
  EDFFXL \block_reg[7][106]  ( .D(block_next[106]), .E(n651), .CK(clk), .Q(
        \block[7][106] ) );
  EDFFXL \block_reg[7][105]  ( .D(block_next[105]), .E(n651), .CK(clk), .Q(
        \block[7][105] ) );
  EDFFXL \block_reg[7][104]  ( .D(block_next[104]), .E(n650), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFXL \block_reg[7][103]  ( .D(block_next[103]), .E(n650), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFXL \block_reg[7][102]  ( .D(block_next[102]), .E(n650), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFXL \block_reg[7][101]  ( .D(block_next[101]), .E(n650), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFXL \block_reg[7][100]  ( .D(block_next[100]), .E(n650), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFXL \block_reg[7][99]  ( .D(block_next[99]), .E(n650), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFXL \block_reg[7][98]  ( .D(block_next[98]), .E(n650), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFXL \block_reg[7][97]  ( .D(block_next[97]), .E(n650), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFXL \block_reg[7][96]  ( .D(block_next[96]), .E(n650), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFXL \block_reg[7][95]  ( .D(block_next[95]), .E(n650), .CK(clk), .Q(
        \block[7][95] ) );
  EDFFXL \block_reg[7][94]  ( .D(block_next[94]), .E(n650), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFXL \block_reg[7][93]  ( .D(block_next[93]), .E(n650), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFXL \block_reg[7][92]  ( .D(block_next[92]), .E(n650), .CK(clk), .Q(
        \block[7][92] ) );
  EDFFXL \block_reg[7][91]  ( .D(block_next[91]), .E(n649), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFXL \block_reg[7][90]  ( .D(block_next[90]), .E(n649), .CK(clk), .Q(
        \block[7][90] ) );
  EDFFXL \block_reg[7][89]  ( .D(block_next[89]), .E(n649), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFXL \block_reg[7][88]  ( .D(block_next[88]), .E(n649), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFXL \block_reg[7][87]  ( .D(block_next[87]), .E(n649), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFXL \block_reg[7][86]  ( .D(block_next[86]), .E(n649), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFXL \block_reg[7][85]  ( .D(block_next[85]), .E(n649), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFXL \block_reg[7][84]  ( .D(block_next[84]), .E(n649), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFXL \block_reg[7][83]  ( .D(block_next[83]), .E(n649), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFXL \block_reg[7][82]  ( .D(block_next[82]), .E(n649), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFXL \block_reg[7][81]  ( .D(block_next[81]), .E(n649), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFXL \block_reg[7][80]  ( .D(block_next[80]), .E(n649), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFXL \block_reg[7][79]  ( .D(block_next[79]), .E(n649), .CK(clk), .Q(
        \block[7][79] ) );
  EDFFXL \block_reg[7][78]  ( .D(block_next[78]), .E(n648), .CK(clk), .Q(
        \block[7][78] ) );
  EDFFXL \block_reg[7][77]  ( .D(block_next[77]), .E(n648), .CK(clk), .Q(
        \block[7][77] ) );
  EDFFXL \block_reg[7][76]  ( .D(block_next[76]), .E(n648), .CK(clk), .Q(
        \block[7][76] ) );
  EDFFXL \block_reg[7][75]  ( .D(block_next[75]), .E(n648), .CK(clk), .Q(
        \block[7][75] ) );
  EDFFXL \block_reg[7][74]  ( .D(block_next[74]), .E(n648), .CK(clk), .Q(
        \block[7][74] ) );
  EDFFXL \block_reg[7][73]  ( .D(block_next[73]), .E(n648), .CK(clk), .Q(
        \block[7][73] ) );
  EDFFXL \block_reg[7][72]  ( .D(block_next[72]), .E(n648), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFXL \block_reg[7][71]  ( .D(block_next[71]), .E(n648), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFXL \block_reg[7][70]  ( .D(block_next[70]), .E(n648), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFXL \block_reg[7][69]  ( .D(block_next[69]), .E(n648), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFXL \block_reg[7][68]  ( .D(block_next[68]), .E(n648), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFXL \block_reg[7][67]  ( .D(block_next[67]), .E(n648), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFXL \block_reg[7][66]  ( .D(block_next[66]), .E(n648), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFXL \block_reg[7][65]  ( .D(block_next[65]), .E(n647), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFXL \block_reg[7][64]  ( .D(block_next[64]), .E(n647), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFX1 \block_reg[7][63]  ( .D(block_next[63]), .E(n647), .CK(clk), .Q(
        \block[7][63] ) );
  EDFFX1 \block_reg[7][53]  ( .D(block_next[53]), .E(n647), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFX1 \block_reg[7][52]  ( .D(block_next[52]), .E(n646), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFX1 \block_reg[7][49]  ( .D(block_next[49]), .E(n646), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFX1 \block_reg[7][41]  ( .D(block_next[41]), .E(n646), .CK(clk), .Q(
        \block[7][41] ) );
  EDFFX1 \block_reg[7][38]  ( .D(block_next[38]), .E(n645), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFX1 \block_reg[7][37]  ( .D(block_next[37]), .E(n645), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFX1 \block_reg[7][36]  ( .D(block_next[36]), .E(n645), .CK(clk), .Q(
        \block[7][36] ) );
  EDFFX1 \block_reg[7][35]  ( .D(block_next[35]), .E(n645), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFX1 \block_reg[7][34]  ( .D(block_next[34]), .E(n645), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFX1 \block_reg[7][32]  ( .D(block_next[32]), .E(n645), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFX1 \block_reg[7][21]  ( .D(block_next[21]), .E(n644), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFX1 \block_reg[7][20]  ( .D(block_next[20]), .E(n644), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFX1 \block_reg[7][19]  ( .D(block_next[19]), .E(n644), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFX1 \block_reg[7][18]  ( .D(block_next[18]), .E(n644), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFX1 \block_reg[7][17]  ( .D(block_next[17]), .E(n644), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFX1 \block_reg[7][16]  ( .D(block_next[16]), .E(n644), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFX1 \block_reg[7][15]  ( .D(block_next[15]), .E(n644), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFX1 \block_reg[7][14]  ( .D(block_next[14]), .E(n644), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFX1 \block_reg[7][13]  ( .D(block_next[13]), .E(n643), .CK(clk), .Q(
        \block[7][13] ) );
  EDFFX1 \block_reg[7][12]  ( .D(block_next[12]), .E(n643), .CK(clk), .Q(
        \block[7][12] ) );
  EDFFX1 \block_reg[7][11]  ( .D(block_next[11]), .E(n643), .CK(clk), .Q(
        \block[7][11] ) );
  EDFFX1 \block_reg[7][10]  ( .D(block_next[10]), .E(n643), .CK(clk), .Q(
        \block[7][10] ) );
  EDFFX1 \block_reg[7][9]  ( .D(block_next[9]), .E(n643), .CK(clk), .Q(
        \block[7][9] ) );
  EDFFX1 \block_reg[7][8]  ( .D(block_next[8]), .E(n643), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFX1 \block_reg[7][7]  ( .D(block_next[7]), .E(n643), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFX1 \block_reg[7][0]  ( .D(block_next[0]), .E(n642), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFXL \block_reg[7][127]  ( .D(block_next[127]), .E(n652), .CK(clk), .Q(
        \block[7][127] ) );
  EDFFXL \block_reg[7][126]  ( .D(block_next[126]), .E(n652), .CK(clk), .Q(
        \block[7][126] ) );
  EDFFXL \block_reg[7][125]  ( .D(block_next[125]), .E(n652), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFXL \block_reg[7][124]  ( .D(block_next[124]), .E(n652), .CK(clk), .Q(
        \block[7][124] ) );
  EDFFXL \block_reg[7][123]  ( .D(block_next[123]), .E(n652), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFXL \block_reg[7][122]  ( .D(block_next[122]), .E(n652), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFXL \block_reg[7][121]  ( .D(block_next[121]), .E(n652), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFXL \block_reg[7][120]  ( .D(block_next[120]), .E(n652), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFXL \block_reg[7][119]  ( .D(block_next[119]), .E(n652), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFXL \block_reg[7][118]  ( .D(block_next[118]), .E(n652), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFXL \block_reg[7][117]  ( .D(block_next[117]), .E(n651), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFXL \block_reg[3][116]  ( .D(block_next[116]), .E(n724), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFXL \block_reg[3][115]  ( .D(block_next[115]), .E(n724), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFXL \block_reg[3][114]  ( .D(block_next[114]), .E(n724), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFXL \block_reg[3][113]  ( .D(block_next[113]), .E(n724), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFXL \block_reg[3][112]  ( .D(block_next[112]), .E(n724), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFXL \block_reg[3][111]  ( .D(block_next[111]), .E(n724), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFXL \block_reg[3][110]  ( .D(block_next[110]), .E(n724), .CK(clk), .Q(
        \block[3][110] ) );
  EDFFXL \block_reg[3][109]  ( .D(block_next[109]), .E(n724), .CK(clk), .Q(
        \block[3][109] ) );
  EDFFXL \block_reg[3][108]  ( .D(block_next[108]), .E(n724), .CK(clk), .Q(
        \block[3][108] ) );
  EDFFXL \block_reg[3][107]  ( .D(block_next[107]), .E(n724), .CK(clk), .Q(
        \block[3][107] ) );
  EDFFXL \block_reg[3][106]  ( .D(block_next[106]), .E(n724), .CK(clk), .Q(
        \block[3][106] ) );
  EDFFXL \block_reg[3][105]  ( .D(block_next[105]), .E(n724), .CK(clk), .Q(
        \block[3][105] ) );
  EDFFXL \block_reg[3][104]  ( .D(block_next[104]), .E(n723), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFXL \block_reg[3][103]  ( .D(block_next[103]), .E(n723), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFXL \block_reg[3][102]  ( .D(block_next[102]), .E(n723), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFXL \block_reg[3][101]  ( .D(block_next[101]), .E(n723), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFXL \block_reg[3][100]  ( .D(block_next[100]), .E(n723), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFXL \block_reg[3][99]  ( .D(block_next[99]), .E(n723), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFXL \block_reg[3][98]  ( .D(block_next[98]), .E(n723), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFXL \block_reg[3][97]  ( .D(block_next[97]), .E(n723), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFXL \block_reg[3][96]  ( .D(block_next[96]), .E(n723), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFXL \block_reg[3][95]  ( .D(block_next[95]), .E(n723), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFXL \block_reg[3][94]  ( .D(block_next[94]), .E(n723), .CK(clk), .Q(
        \block[3][94] ) );
  EDFFXL \block_reg[3][93]  ( .D(block_next[93]), .E(n723), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFXL \block_reg[3][92]  ( .D(block_next[92]), .E(n723), .CK(clk), .Q(
        \block[3][92] ) );
  EDFFXL \block_reg[3][91]  ( .D(block_next[91]), .E(n722), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFXL \block_reg[3][90]  ( .D(block_next[90]), .E(n722), .CK(clk), .Q(
        \block[3][90] ) );
  EDFFXL \block_reg[3][89]  ( .D(block_next[89]), .E(n722), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFXL \block_reg[3][88]  ( .D(block_next[88]), .E(n722), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFXL \block_reg[3][87]  ( .D(block_next[87]), .E(n722), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFXL \block_reg[3][86]  ( .D(block_next[86]), .E(n722), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFXL \block_reg[3][85]  ( .D(block_next[85]), .E(n722), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFXL \block_reg[3][84]  ( .D(block_next[84]), .E(n722), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFXL \block_reg[3][83]  ( .D(block_next[83]), .E(n722), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFXL \block_reg[3][82]  ( .D(block_next[82]), .E(n722), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFXL \block_reg[3][81]  ( .D(block_next[81]), .E(n722), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFXL \block_reg[3][80]  ( .D(block_next[80]), .E(n722), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFXL \block_reg[3][79]  ( .D(block_next[79]), .E(n722), .CK(clk), .Q(
        \block[3][79] ) );
  EDFFXL \block_reg[3][78]  ( .D(block_next[78]), .E(n721), .CK(clk), .Q(
        \block[3][78] ) );
  EDFFXL \block_reg[3][77]  ( .D(block_next[77]), .E(n721), .CK(clk), .Q(
        \block[3][77] ) );
  EDFFXL \block_reg[3][76]  ( .D(block_next[76]), .E(n721), .CK(clk), .Q(
        \block[3][76] ) );
  EDFFXL \block_reg[3][75]  ( .D(block_next[75]), .E(n721), .CK(clk), .Q(
        \block[3][75] ) );
  EDFFXL \block_reg[3][74]  ( .D(block_next[74]), .E(n721), .CK(clk), .Q(
        \block[3][74] ) );
  EDFFXL \block_reg[3][73]  ( .D(block_next[73]), .E(n721), .CK(clk), .Q(
        \block[3][73] ) );
  EDFFXL \block_reg[3][72]  ( .D(block_next[72]), .E(n721), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFXL \block_reg[3][71]  ( .D(block_next[71]), .E(n721), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFXL \block_reg[3][70]  ( .D(block_next[70]), .E(n721), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFXL \block_reg[3][69]  ( .D(block_next[69]), .E(n721), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFXL \block_reg[3][68]  ( .D(block_next[68]), .E(n721), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFXL \block_reg[3][67]  ( .D(block_next[67]), .E(n721), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFXL \block_reg[3][66]  ( .D(block_next[66]), .E(n721), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFXL \block_reg[3][65]  ( .D(block_next[65]), .E(n720), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFXL \block_reg[3][64]  ( .D(block_next[64]), .E(n720), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFX1 \block_reg[3][63]  ( .D(block_next[63]), .E(n720), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFX1 \block_reg[3][53]  ( .D(block_next[53]), .E(n720), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFX1 \block_reg[3][52]  ( .D(block_next[52]), .E(n719), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFX1 \block_reg[3][49]  ( .D(block_next[49]), .E(n719), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFX1 \block_reg[3][41]  ( .D(block_next[41]), .E(n719), .CK(clk), .Q(
        \block[3][41] ) );
  EDFFX1 \block_reg[3][38]  ( .D(block_next[38]), .E(n718), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFX1 \block_reg[3][37]  ( .D(block_next[37]), .E(n718), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFX1 \block_reg[3][36]  ( .D(block_next[36]), .E(n718), .CK(clk), .Q(
        \block[3][36] ) );
  EDFFX1 \block_reg[3][35]  ( .D(block_next[35]), .E(n718), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFX1 \block_reg[3][34]  ( .D(block_next[34]), .E(n718), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFX1 \block_reg[3][32]  ( .D(block_next[32]), .E(n718), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFX1 \block_reg[3][21]  ( .D(block_next[21]), .E(n717), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFX1 \block_reg[3][20]  ( .D(block_next[20]), .E(n717), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFX1 \block_reg[3][19]  ( .D(block_next[19]), .E(n717), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFX1 \block_reg[3][18]  ( .D(block_next[18]), .E(n717), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFX1 \block_reg[3][17]  ( .D(block_next[17]), .E(n717), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFX1 \block_reg[3][16]  ( .D(block_next[16]), .E(n717), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFX1 \block_reg[3][15]  ( .D(block_next[15]), .E(n717), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFX1 \block_reg[3][14]  ( .D(block_next[14]), .E(n717), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFX1 \block_reg[3][13]  ( .D(block_next[13]), .E(n716), .CK(clk), .Q(
        \block[3][13] ) );
  EDFFX1 \block_reg[3][12]  ( .D(block_next[12]), .E(n716), .CK(clk), .Q(
        \block[3][12] ) );
  EDFFX1 \block_reg[3][11]  ( .D(block_next[11]), .E(n716), .CK(clk), .Q(
        \block[3][11] ) );
  EDFFX1 \block_reg[3][10]  ( .D(block_next[10]), .E(n716), .CK(clk), .Q(
        \block[3][10] ) );
  EDFFX1 \block_reg[3][9]  ( .D(block_next[9]), .E(n716), .CK(clk), .Q(
        \block[3][9] ) );
  EDFFX1 \block_reg[3][8]  ( .D(block_next[8]), .E(n716), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFX1 \block_reg[3][7]  ( .D(block_next[7]), .E(n716), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFX1 \block_reg[3][0]  ( .D(block_next[0]), .E(n715), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFXL \block_reg[3][127]  ( .D(block_next[127]), .E(n725), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFXL \block_reg[3][126]  ( .D(block_next[126]), .E(n725), .CK(clk), .Q(
        \block[3][126] ) );
  EDFFXL \block_reg[3][125]  ( .D(block_next[125]), .E(n725), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFXL \block_reg[3][124]  ( .D(block_next[124]), .E(n725), .CK(clk), .Q(
        \block[3][124] ) );
  EDFFXL \block_reg[3][123]  ( .D(block_next[123]), .E(n725), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFXL \block_reg[3][122]  ( .D(block_next[122]), .E(n725), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFXL \block_reg[3][121]  ( .D(block_next[121]), .E(n725), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFXL \block_reg[3][120]  ( .D(block_next[120]), .E(n725), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFXL \block_reg[3][119]  ( .D(block_next[119]), .E(n725), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFXL \block_reg[3][118]  ( .D(block_next[118]), .E(n725), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFXL \block_reg[3][117]  ( .D(block_next[117]), .E(n724), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFXL \block_reg[5][116]  ( .D(block_next[116]), .E(n689), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFXL \block_reg[5][115]  ( .D(block_next[115]), .E(n689), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFXL \block_reg[5][114]  ( .D(block_next[114]), .E(n689), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFXL \block_reg[5][113]  ( .D(block_next[113]), .E(n689), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFXL \block_reg[5][112]  ( .D(block_next[112]), .E(n689), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFXL \block_reg[5][111]  ( .D(block_next[111]), .E(n689), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFXL \block_reg[5][110]  ( .D(block_next[110]), .E(n689), .CK(clk), .Q(
        \block[5][110] ) );
  EDFFXL \block_reg[5][109]  ( .D(block_next[109]), .E(n689), .CK(clk), .Q(
        \block[5][109] ) );
  EDFFXL \block_reg[5][108]  ( .D(block_next[108]), .E(n689), .CK(clk), .Q(
        \block[5][108] ) );
  EDFFXL \block_reg[5][107]  ( .D(block_next[107]), .E(n689), .CK(clk), .Q(
        \block[5][107] ) );
  EDFFXL \block_reg[5][106]  ( .D(block_next[106]), .E(n689), .CK(clk), .Q(
        \block[5][106] ) );
  EDFFXL \block_reg[5][105]  ( .D(block_next[105]), .E(n689), .CK(clk), .Q(
        \block[5][105] ) );
  EDFFXL \block_reg[5][104]  ( .D(block_next[104]), .E(n688), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFXL \block_reg[5][103]  ( .D(block_next[103]), .E(n688), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFXL \block_reg[5][102]  ( .D(block_next[102]), .E(n688), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFXL \block_reg[5][101]  ( .D(block_next[101]), .E(n688), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFXL \block_reg[5][100]  ( .D(block_next[100]), .E(n688), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFXL \block_reg[5][99]  ( .D(block_next[99]), .E(n688), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFXL \block_reg[5][98]  ( .D(block_next[98]), .E(n688), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFXL \block_reg[5][97]  ( .D(block_next[97]), .E(n688), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFXL \block_reg[5][96]  ( .D(block_next[96]), .E(n688), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFXL \block_reg[5][95]  ( .D(block_next[95]), .E(n688), .CK(clk), .Q(
        \block[5][95] ) );
  EDFFXL \block_reg[5][94]  ( .D(block_next[94]), .E(n688), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFXL \block_reg[5][93]  ( .D(block_next[93]), .E(n688), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFXL \block_reg[5][92]  ( .D(block_next[92]), .E(n688), .CK(clk), .Q(
        \block[5][92] ) );
  EDFFXL \block_reg[5][91]  ( .D(block_next[91]), .E(n687), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFXL \block_reg[5][90]  ( .D(block_next[90]), .E(n687), .CK(clk), .Q(
        \block[5][90] ) );
  EDFFXL \block_reg[5][89]  ( .D(block_next[89]), .E(n687), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFXL \block_reg[5][88]  ( .D(block_next[88]), .E(n687), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFXL \block_reg[5][87]  ( .D(block_next[87]), .E(n687), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFXL \block_reg[5][86]  ( .D(block_next[86]), .E(n687), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFXL \block_reg[5][85]  ( .D(block_next[85]), .E(n687), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFXL \block_reg[5][84]  ( .D(block_next[84]), .E(n687), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFXL \block_reg[5][83]  ( .D(block_next[83]), .E(n687), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFXL \block_reg[5][82]  ( .D(block_next[82]), .E(n687), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFXL \block_reg[5][81]  ( .D(block_next[81]), .E(n687), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFXL \block_reg[5][80]  ( .D(block_next[80]), .E(n687), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFXL \block_reg[5][79]  ( .D(block_next[79]), .E(n687), .CK(clk), .Q(
        \block[5][79] ) );
  EDFFXL \block_reg[5][78]  ( .D(block_next[78]), .E(n686), .CK(clk), .Q(
        \block[5][78] ) );
  EDFFXL \block_reg[5][77]  ( .D(block_next[77]), .E(n686), .CK(clk), .Q(
        \block[5][77] ) );
  EDFFXL \block_reg[5][76]  ( .D(block_next[76]), .E(n686), .CK(clk), .Q(
        \block[5][76] ) );
  EDFFXL \block_reg[5][75]  ( .D(block_next[75]), .E(n686), .CK(clk), .Q(
        \block[5][75] ) );
  EDFFXL \block_reg[5][74]  ( .D(block_next[74]), .E(n686), .CK(clk), .Q(
        \block[5][74] ) );
  EDFFXL \block_reg[5][73]  ( .D(block_next[73]), .E(n686), .CK(clk), .Q(
        \block[5][73] ) );
  EDFFXL \block_reg[5][72]  ( .D(block_next[72]), .E(n686), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFXL \block_reg[5][71]  ( .D(block_next[71]), .E(n686), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFXL \block_reg[5][70]  ( .D(block_next[70]), .E(n686), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFXL \block_reg[5][69]  ( .D(block_next[69]), .E(n686), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFXL \block_reg[5][68]  ( .D(block_next[68]), .E(n686), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFXL \block_reg[5][67]  ( .D(block_next[67]), .E(n686), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFXL \block_reg[5][66]  ( .D(block_next[66]), .E(n686), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFXL \block_reg[5][65]  ( .D(block_next[65]), .E(n685), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFXL \block_reg[5][64]  ( .D(block_next[64]), .E(n685), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFX1 \block_reg[5][63]  ( .D(block_next[63]), .E(n685), .CK(clk), .Q(
        \block[5][63] ) );
  EDFFX1 \block_reg[5][53]  ( .D(block_next[53]), .E(n685), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFX1 \block_reg[5][52]  ( .D(block_next[52]), .E(n684), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFX1 \block_reg[5][49]  ( .D(block_next[49]), .E(n684), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFX1 \block_reg[5][41]  ( .D(block_next[41]), .E(n684), .CK(clk), .Q(
        \block[5][41] ) );
  EDFFX1 \block_reg[5][38]  ( .D(block_next[38]), .E(n683), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFX1 \block_reg[5][37]  ( .D(block_next[37]), .E(n683), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFX1 \block_reg[5][36]  ( .D(block_next[36]), .E(n683), .CK(clk), .Q(
        \block[5][36] ) );
  EDFFX1 \block_reg[5][35]  ( .D(block_next[35]), .E(n683), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFX1 \block_reg[5][32]  ( .D(block_next[32]), .E(n683), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFX1 \block_reg[5][21]  ( .D(block_next[21]), .E(n682), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFX1 \block_reg[5][20]  ( .D(block_next[20]), .E(n682), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFX1 \block_reg[5][19]  ( .D(block_next[19]), .E(n682), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFX1 \block_reg[5][18]  ( .D(block_next[18]), .E(n682), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFX1 \block_reg[5][17]  ( .D(block_next[17]), .E(n682), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFX1 \block_reg[5][16]  ( .D(block_next[16]), .E(n682), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFX1 \block_reg[5][15]  ( .D(block_next[15]), .E(n682), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFX1 \block_reg[5][14]  ( .D(block_next[14]), .E(n682), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFX1 \block_reg[5][13]  ( .D(block_next[13]), .E(n681), .CK(clk), .Q(
        \block[5][13] ) );
  EDFFX1 \block_reg[5][12]  ( .D(block_next[12]), .E(n681), .CK(clk), .Q(
        \block[5][12] ) );
  EDFFX1 \block_reg[5][11]  ( .D(block_next[11]), .E(n681), .CK(clk), .Q(
        \block[5][11] ) );
  EDFFX1 \block_reg[5][10]  ( .D(block_next[10]), .E(n681), .CK(clk), .Q(
        \block[5][10] ) );
  EDFFX1 \block_reg[5][9]  ( .D(block_next[9]), .E(n681), .CK(clk), .Q(
        \block[5][9] ) );
  EDFFX1 \block_reg[5][8]  ( .D(block_next[8]), .E(n681), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFX1 \block_reg[5][7]  ( .D(block_next[7]), .E(n681), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFX1 \block_reg[5][0]  ( .D(block_next[0]), .E(n680), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFXL \block_reg[5][127]  ( .D(block_next[127]), .E(n690), .CK(clk), .Q(
        \block[5][127] ) );
  EDFFXL \block_reg[5][126]  ( .D(block_next[126]), .E(n690), .CK(clk), .Q(
        \block[5][126] ) );
  EDFFXL \block_reg[5][125]  ( .D(block_next[125]), .E(n690), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFXL \block_reg[5][124]  ( .D(block_next[124]), .E(n690), .CK(clk), .Q(
        \block[5][124] ) );
  EDFFXL \block_reg[5][123]  ( .D(block_next[123]), .E(n690), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFXL \block_reg[5][122]  ( .D(block_next[122]), .E(n690), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFXL \block_reg[5][121]  ( .D(block_next[121]), .E(n690), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFXL \block_reg[5][120]  ( .D(block_next[120]), .E(n690), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFXL \block_reg[5][119]  ( .D(block_next[119]), .E(n690), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFXL \block_reg[5][118]  ( .D(block_next[118]), .E(n690), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFXL \block_reg[5][117]  ( .D(block_next[117]), .E(n689), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFXL \block_reg[1][116]  ( .D(block_next[116]), .E(n758), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFXL \block_reg[1][115]  ( .D(block_next[115]), .E(n758), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFXL \block_reg[1][114]  ( .D(block_next[114]), .E(n758), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFXL \block_reg[1][113]  ( .D(block_next[113]), .E(n758), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFXL \block_reg[1][112]  ( .D(block_next[112]), .E(n758), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFXL \block_reg[1][111]  ( .D(block_next[111]), .E(n758), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFXL \block_reg[1][110]  ( .D(block_next[110]), .E(n758), .CK(clk), .Q(
        \block[1][110] ) );
  EDFFXL \block_reg[1][109]  ( .D(block_next[109]), .E(n758), .CK(clk), .Q(
        \block[1][109] ) );
  EDFFXL \block_reg[1][108]  ( .D(block_next[108]), .E(n758), .CK(clk), .Q(
        \block[1][108] ) );
  EDFFXL \block_reg[1][107]  ( .D(block_next[107]), .E(n758), .CK(clk), .Q(
        \block[1][107] ) );
  EDFFXL \block_reg[1][106]  ( .D(block_next[106]), .E(n758), .CK(clk), .Q(
        \block[1][106] ) );
  EDFFXL \block_reg[1][105]  ( .D(block_next[105]), .E(n758), .CK(clk), .Q(
        \block[1][105] ) );
  EDFFXL \block_reg[1][104]  ( .D(block_next[104]), .E(n757), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFXL \block_reg[1][103]  ( .D(block_next[103]), .E(n757), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFXL \block_reg[1][102]  ( .D(block_next[102]), .E(n757), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFXL \block_reg[1][101]  ( .D(block_next[101]), .E(n757), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFXL \block_reg[1][100]  ( .D(block_next[100]), .E(n757), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFXL \block_reg[1][99]  ( .D(block_next[99]), .E(n757), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFXL \block_reg[1][98]  ( .D(block_next[98]), .E(n757), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFXL \block_reg[1][97]  ( .D(block_next[97]), .E(n757), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFXL \block_reg[1][96]  ( .D(block_next[96]), .E(n757), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFXL \block_reg[1][95]  ( .D(block_next[95]), .E(n757), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFXL \block_reg[1][94]  ( .D(block_next[94]), .E(n757), .CK(clk), .Q(
        \block[1][94] ) );
  EDFFXL \block_reg[1][93]  ( .D(block_next[93]), .E(n757), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFXL \block_reg[1][92]  ( .D(block_next[92]), .E(n757), .CK(clk), .Q(
        \block[1][92] ) );
  EDFFXL \block_reg[1][91]  ( .D(block_next[91]), .E(n756), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFXL \block_reg[1][90]  ( .D(block_next[90]), .E(n756), .CK(clk), .Q(
        \block[1][90] ) );
  EDFFXL \block_reg[1][89]  ( .D(block_next[89]), .E(n756), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFXL \block_reg[1][88]  ( .D(block_next[88]), .E(n756), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFXL \block_reg[1][87]  ( .D(block_next[87]), .E(n756), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFXL \block_reg[1][86]  ( .D(block_next[86]), .E(n756), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFXL \block_reg[1][85]  ( .D(block_next[85]), .E(n756), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFXL \block_reg[1][84]  ( .D(block_next[84]), .E(n756), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFXL \block_reg[1][83]  ( .D(block_next[83]), .E(n756), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFXL \block_reg[1][82]  ( .D(block_next[82]), .E(n756), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFXL \block_reg[1][81]  ( .D(block_next[81]), .E(n756), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFXL \block_reg[1][80]  ( .D(block_next[80]), .E(n756), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFXL \block_reg[1][79]  ( .D(block_next[79]), .E(n756), .CK(clk), .Q(
        \block[1][79] ) );
  EDFFXL \block_reg[1][78]  ( .D(block_next[78]), .E(n755), .CK(clk), .Q(
        \block[1][78] ) );
  EDFFXL \block_reg[1][77]  ( .D(block_next[77]), .E(n755), .CK(clk), .Q(
        \block[1][77] ) );
  EDFFXL \block_reg[1][76]  ( .D(block_next[76]), .E(n755), .CK(clk), .Q(
        \block[1][76] ) );
  EDFFXL \block_reg[1][75]  ( .D(block_next[75]), .E(n755), .CK(clk), .Q(
        \block[1][75] ) );
  EDFFXL \block_reg[1][74]  ( .D(block_next[74]), .E(n755), .CK(clk), .Q(
        \block[1][74] ) );
  EDFFXL \block_reg[1][73]  ( .D(block_next[73]), .E(n755), .CK(clk), .Q(
        \block[1][73] ) );
  EDFFXL \block_reg[1][72]  ( .D(block_next[72]), .E(n755), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFXL \block_reg[1][71]  ( .D(block_next[71]), .E(n755), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFXL \block_reg[1][70]  ( .D(block_next[70]), .E(n755), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFXL \block_reg[1][69]  ( .D(block_next[69]), .E(n755), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFXL \block_reg[1][68]  ( .D(block_next[68]), .E(n755), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFXL \block_reg[1][67]  ( .D(block_next[67]), .E(n755), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFXL \block_reg[1][66]  ( .D(block_next[66]), .E(n755), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFXL \block_reg[1][65]  ( .D(block_next[65]), .E(n754), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFXL \block_reg[1][64]  ( .D(block_next[64]), .E(n754), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFX1 \block_reg[1][63]  ( .D(block_next[63]), .E(n754), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFX1 \block_reg[1][53]  ( .D(block_next[53]), .E(n754), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFX1 \block_reg[1][52]  ( .D(block_next[52]), .E(n753), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFX1 \block_reg[1][49]  ( .D(block_next[49]), .E(n753), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFX1 \block_reg[1][41]  ( .D(block_next[41]), .E(n753), .CK(clk), .Q(
        \block[1][41] ) );
  EDFFX1 \block_reg[1][38]  ( .D(block_next[38]), .E(n752), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFX1 \block_reg[1][37]  ( .D(block_next[37]), .E(n752), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFX1 \block_reg[1][36]  ( .D(block_next[36]), .E(n752), .CK(clk), .Q(
        \block[1][36] ) );
  EDFFX1 \block_reg[1][35]  ( .D(block_next[35]), .E(n752), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFX1 \block_reg[1][32]  ( .D(block_next[32]), .E(n752), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFX1 \block_reg[1][21]  ( .D(block_next[21]), .E(n751), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFX1 \block_reg[1][20]  ( .D(block_next[20]), .E(n751), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFX1 \block_reg[1][19]  ( .D(block_next[19]), .E(n751), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFX1 \block_reg[1][18]  ( .D(block_next[18]), .E(n751), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFX1 \block_reg[1][17]  ( .D(block_next[17]), .E(n751), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFX1 \block_reg[1][16]  ( .D(block_next[16]), .E(n751), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFX1 \block_reg[1][15]  ( .D(block_next[15]), .E(n751), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFX1 \block_reg[1][14]  ( .D(block_next[14]), .E(n751), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFX1 \block_reg[1][13]  ( .D(block_next[13]), .E(n750), .CK(clk), .Q(
        \block[1][13] ) );
  EDFFX1 \block_reg[1][12]  ( .D(block_next[12]), .E(n750), .CK(clk), .Q(
        \block[1][12] ) );
  EDFFX1 \block_reg[1][11]  ( .D(block_next[11]), .E(n750), .CK(clk), .Q(
        \block[1][11] ) );
  EDFFX1 \block_reg[1][10]  ( .D(block_next[10]), .E(n750), .CK(clk), .Q(
        \block[1][10] ) );
  EDFFX1 \block_reg[1][9]  ( .D(block_next[9]), .E(n750), .CK(clk), .Q(
        \block[1][9] ) );
  EDFFX1 \block_reg[1][8]  ( .D(block_next[8]), .E(n750), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFX1 \block_reg[1][7]  ( .D(block_next[7]), .E(n750), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFX1 \block_reg[1][0]  ( .D(block_next[0]), .E(n749), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFXL \block_reg[1][127]  ( .D(block_next[127]), .E(n759), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFXL \block_reg[1][126]  ( .D(block_next[126]), .E(n759), .CK(clk), .Q(
        \block[1][126] ) );
  EDFFXL \block_reg[1][125]  ( .D(block_next[125]), .E(n759), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFXL \block_reg[1][124]  ( .D(block_next[124]), .E(n759), .CK(clk), .Q(
        \block[1][124] ) );
  EDFFXL \block_reg[1][123]  ( .D(block_next[123]), .E(n759), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFXL \block_reg[1][122]  ( .D(block_next[122]), .E(n759), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFXL \block_reg[1][121]  ( .D(block_next[121]), .E(n759), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFXL \block_reg[1][120]  ( .D(block_next[120]), .E(n759), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFXL \block_reg[1][119]  ( .D(block_next[119]), .E(n759), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFXL \block_reg[1][118]  ( .D(block_next[118]), .E(n759), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFXL \block_reg[1][117]  ( .D(block_next[117]), .E(n758), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFXL \block_reg[4][116]  ( .D(block_next[116]), .E(n706), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFXL \block_reg[4][115]  ( .D(block_next[115]), .E(n706), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFXL \block_reg[4][114]  ( .D(block_next[114]), .E(n706), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFXL \block_reg[4][113]  ( .D(block_next[113]), .E(n706), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFXL \block_reg[4][112]  ( .D(block_next[112]), .E(n706), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFXL \block_reg[4][111]  ( .D(block_next[111]), .E(n706), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFXL \block_reg[4][110]  ( .D(block_next[110]), .E(n706), .CK(clk), .Q(
        \block[4][110] ) );
  EDFFXL \block_reg[4][109]  ( .D(block_next[109]), .E(n706), .CK(clk), .Q(
        \block[4][109] ) );
  EDFFXL \block_reg[4][108]  ( .D(block_next[108]), .E(n706), .CK(clk), .Q(
        \block[4][108] ) );
  EDFFXL \block_reg[4][107]  ( .D(block_next[107]), .E(n706), .CK(clk), .Q(
        \block[4][107] ) );
  EDFFXL \block_reg[4][106]  ( .D(block_next[106]), .E(n706), .CK(clk), .Q(
        \block[4][106] ) );
  EDFFXL \block_reg[4][105]  ( .D(block_next[105]), .E(n706), .CK(clk), .Q(
        \block[4][105] ) );
  EDFFXL \block_reg[4][104]  ( .D(block_next[104]), .E(n705), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFXL \block_reg[4][103]  ( .D(block_next[103]), .E(n705), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFXL \block_reg[4][102]  ( .D(block_next[102]), .E(n705), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFXL \block_reg[4][101]  ( .D(block_next[101]), .E(n705), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFXL \block_reg[4][100]  ( .D(block_next[100]), .E(n705), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFXL \block_reg[4][99]  ( .D(block_next[99]), .E(n705), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFXL \block_reg[4][98]  ( .D(block_next[98]), .E(n705), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFXL \block_reg[4][97]  ( .D(block_next[97]), .E(n705), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFXL \block_reg[4][96]  ( .D(block_next[96]), .E(n705), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFXL \block_reg[4][95]  ( .D(block_next[95]), .E(n705), .CK(clk), .Q(
        \block[4][95] ) );
  EDFFXL \block_reg[4][94]  ( .D(block_next[94]), .E(n705), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFXL \block_reg[4][93]  ( .D(block_next[93]), .E(n705), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFXL \block_reg[4][92]  ( .D(block_next[92]), .E(n705), .CK(clk), .Q(
        \block[4][92] ) );
  EDFFXL \block_reg[4][91]  ( .D(block_next[91]), .E(n704), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFXL \block_reg[4][90]  ( .D(block_next[90]), .E(n704), .CK(clk), .Q(
        \block[4][90] ) );
  EDFFXL \block_reg[4][89]  ( .D(block_next[89]), .E(n704), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFXL \block_reg[4][88]  ( .D(block_next[88]), .E(n704), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFXL \block_reg[4][87]  ( .D(block_next[87]), .E(n704), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFXL \block_reg[4][86]  ( .D(block_next[86]), .E(n704), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFXL \block_reg[4][85]  ( .D(block_next[85]), .E(n704), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFXL \block_reg[4][84]  ( .D(block_next[84]), .E(n704), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFXL \block_reg[4][83]  ( .D(block_next[83]), .E(n704), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFXL \block_reg[4][82]  ( .D(block_next[82]), .E(n704), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFXL \block_reg[4][81]  ( .D(block_next[81]), .E(n704), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFXL \block_reg[4][80]  ( .D(block_next[80]), .E(n704), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFXL \block_reg[4][79]  ( .D(block_next[79]), .E(n704), .CK(clk), .Q(
        \block[4][79] ) );
  EDFFXL \block_reg[4][78]  ( .D(block_next[78]), .E(n703), .CK(clk), .Q(
        \block[4][78] ) );
  EDFFXL \block_reg[4][77]  ( .D(block_next[77]), .E(n703), .CK(clk), .Q(
        \block[4][77] ) );
  EDFFXL \block_reg[4][76]  ( .D(block_next[76]), .E(n703), .CK(clk), .Q(
        \block[4][76] ) );
  EDFFXL \block_reg[4][75]  ( .D(block_next[75]), .E(n703), .CK(clk), .Q(
        \block[4][75] ) );
  EDFFXL \block_reg[4][74]  ( .D(block_next[74]), .E(n703), .CK(clk), .Q(
        \block[4][74] ) );
  EDFFXL \block_reg[4][73]  ( .D(block_next[73]), .E(n703), .CK(clk), .Q(
        \block[4][73] ) );
  EDFFXL \block_reg[4][72]  ( .D(block_next[72]), .E(n703), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFXL \block_reg[4][71]  ( .D(block_next[71]), .E(n703), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFXL \block_reg[4][70]  ( .D(block_next[70]), .E(n703), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFXL \block_reg[4][69]  ( .D(block_next[69]), .E(n703), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFXL \block_reg[4][68]  ( .D(block_next[68]), .E(n703), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFXL \block_reg[4][67]  ( .D(block_next[67]), .E(n703), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFXL \block_reg[4][66]  ( .D(block_next[66]), .E(n703), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFXL \block_reg[4][65]  ( .D(block_next[65]), .E(n702), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFXL \block_reg[4][64]  ( .D(block_next[64]), .E(n702), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFX1 \block_reg[4][63]  ( .D(block_next[63]), .E(n702), .CK(clk), .Q(
        \block[4][63] ) );
  EDFFX1 \block_reg[4][53]  ( .D(block_next[53]), .E(n702), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFX1 \block_reg[4][52]  ( .D(block_next[52]), .E(n701), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFX1 \block_reg[4][49]  ( .D(block_next[49]), .E(n701), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFX1 \block_reg[4][41]  ( .D(block_next[41]), .E(n701), .CK(clk), .Q(
        \block[4][41] ) );
  EDFFX1 \block_reg[4][38]  ( .D(block_next[38]), .E(n700), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFX1 \block_reg[4][37]  ( .D(block_next[37]), .E(n700), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFX1 \block_reg[4][36]  ( .D(block_next[36]), .E(n700), .CK(clk), .Q(
        \block[4][36] ) );
  EDFFX1 \block_reg[4][35]  ( .D(block_next[35]), .E(n700), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFX1 \block_reg[4][32]  ( .D(block_next[32]), .E(n700), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFX1 \block_reg[4][21]  ( .D(block_next[21]), .E(n699), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFX1 \block_reg[4][20]  ( .D(block_next[20]), .E(n699), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFX1 \block_reg[4][19]  ( .D(block_next[19]), .E(n699), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFX1 \block_reg[4][18]  ( .D(block_next[18]), .E(n699), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFX1 \block_reg[4][17]  ( .D(block_next[17]), .E(n699), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFX1 \block_reg[4][16]  ( .D(block_next[16]), .E(n699), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFX1 \block_reg[4][15]  ( .D(block_next[15]), .E(n699), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFX1 \block_reg[4][14]  ( .D(block_next[14]), .E(n699), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFX1 \block_reg[4][13]  ( .D(block_next[13]), .E(n698), .CK(clk), .Q(
        \block[4][13] ) );
  EDFFX1 \block_reg[4][12]  ( .D(block_next[12]), .E(n698), .CK(clk), .Q(
        \block[4][12] ) );
  EDFFX1 \block_reg[4][11]  ( .D(block_next[11]), .E(n698), .CK(clk), .Q(
        \block[4][11] ) );
  EDFFX1 \block_reg[4][10]  ( .D(block_next[10]), .E(n698), .CK(clk), .Q(
        \block[4][10] ) );
  EDFFX1 \block_reg[4][9]  ( .D(block_next[9]), .E(n698), .CK(clk), .Q(
        \block[4][9] ) );
  EDFFX1 \block_reg[4][8]  ( .D(block_next[8]), .E(n698), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFX1 \block_reg[4][7]  ( .D(block_next[7]), .E(n698), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFX1 \block_reg[4][0]  ( .D(block_next[0]), .E(n697), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFXL \block_reg[4][127]  ( .D(block_next[127]), .E(n707), .CK(clk), .Q(
        \block[4][127] ) );
  EDFFXL \block_reg[4][126]  ( .D(block_next[126]), .E(n707), .CK(clk), .Q(
        \block[4][126] ) );
  EDFFXL \block_reg[4][125]  ( .D(block_next[125]), .E(n707), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFXL \block_reg[4][124]  ( .D(block_next[124]), .E(n707), .CK(clk), .Q(
        \block[4][124] ) );
  EDFFXL \block_reg[4][123]  ( .D(block_next[123]), .E(n707), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFXL \block_reg[4][122]  ( .D(block_next[122]), .E(n707), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFXL \block_reg[4][121]  ( .D(block_next[121]), .E(n707), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFXL \block_reg[4][120]  ( .D(block_next[120]), .E(n707), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFXL \block_reg[4][119]  ( .D(block_next[119]), .E(n707), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFXL \block_reg[4][118]  ( .D(block_next[118]), .E(n707), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFXL \block_reg[4][117]  ( .D(block_next[117]), .E(n706), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFXL \block_reg[0][116]  ( .D(block_next[116]), .E(n777), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFXL \block_reg[0][115]  ( .D(block_next[115]), .E(n777), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFXL \block_reg[0][114]  ( .D(block_next[114]), .E(n777), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFXL \block_reg[0][113]  ( .D(block_next[113]), .E(n777), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFXL \block_reg[0][112]  ( .D(block_next[112]), .E(n777), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFXL \block_reg[0][111]  ( .D(block_next[111]), .E(n777), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFXL \block_reg[0][110]  ( .D(block_next[110]), .E(n777), .CK(clk), .Q(
        \block[0][110] ) );
  EDFFXL \block_reg[0][109]  ( .D(block_next[109]), .E(n777), .CK(clk), .Q(
        \block[0][109] ) );
  EDFFXL \block_reg[0][108]  ( .D(block_next[108]), .E(n777), .CK(clk), .Q(
        \block[0][108] ) );
  EDFFXL \block_reg[0][107]  ( .D(block_next[107]), .E(n777), .CK(clk), .Q(
        \block[0][107] ) );
  EDFFXL \block_reg[0][106]  ( .D(block_next[106]), .E(n777), .CK(clk), .Q(
        \block[0][106] ) );
  EDFFXL \block_reg[0][105]  ( .D(block_next[105]), .E(n777), .CK(clk), .Q(
        \block[0][105] ) );
  EDFFXL \block_reg[0][104]  ( .D(block_next[104]), .E(n776), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFXL \block_reg[0][103]  ( .D(block_next[103]), .E(n776), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFXL \block_reg[0][102]  ( .D(block_next[102]), .E(n776), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFXL \block_reg[0][101]  ( .D(block_next[101]), .E(n776), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFXL \block_reg[0][100]  ( .D(block_next[100]), .E(n776), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFXL \block_reg[0][99]  ( .D(block_next[99]), .E(n776), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFXL \block_reg[0][98]  ( .D(block_next[98]), .E(n776), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFXL \block_reg[0][97]  ( .D(block_next[97]), .E(n776), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFXL \block_reg[0][96]  ( .D(block_next[96]), .E(n776), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFXL \block_reg[0][95]  ( .D(block_next[95]), .E(n776), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFXL \block_reg[0][94]  ( .D(block_next[94]), .E(n776), .CK(clk), .Q(
        \block[0][94] ) );
  EDFFXL \block_reg[0][93]  ( .D(block_next[93]), .E(n776), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFXL \block_reg[0][92]  ( .D(block_next[92]), .E(n776), .CK(clk), .Q(
        \block[0][92] ) );
  EDFFXL \block_reg[0][91]  ( .D(block_next[91]), .E(n775), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFXL \block_reg[0][90]  ( .D(block_next[90]), .E(n775), .CK(clk), .Q(
        \block[0][90] ) );
  EDFFXL \block_reg[0][89]  ( .D(block_next[89]), .E(n775), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFXL \block_reg[0][88]  ( .D(block_next[88]), .E(n775), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFXL \block_reg[0][87]  ( .D(block_next[87]), .E(n775), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFXL \block_reg[0][86]  ( .D(block_next[86]), .E(n775), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFXL \block_reg[0][85]  ( .D(block_next[85]), .E(n775), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFXL \block_reg[0][84]  ( .D(block_next[84]), .E(n775), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFXL \block_reg[0][83]  ( .D(block_next[83]), .E(n775), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFXL \block_reg[0][82]  ( .D(block_next[82]), .E(n775), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFXL \block_reg[0][81]  ( .D(block_next[81]), .E(n775), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFXL \block_reg[0][80]  ( .D(block_next[80]), .E(n775), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFXL \block_reg[0][79]  ( .D(block_next[79]), .E(n775), .CK(clk), .Q(
        \block[0][79] ) );
  EDFFXL \block_reg[0][78]  ( .D(block_next[78]), .E(n774), .CK(clk), .Q(
        \block[0][78] ) );
  EDFFXL \block_reg[0][77]  ( .D(block_next[77]), .E(n774), .CK(clk), .Q(
        \block[0][77] ) );
  EDFFXL \block_reg[0][76]  ( .D(block_next[76]), .E(n774), .CK(clk), .Q(
        \block[0][76] ) );
  EDFFXL \block_reg[0][75]  ( .D(block_next[75]), .E(n774), .CK(clk), .Q(
        \block[0][75] ) );
  EDFFXL \block_reg[0][74]  ( .D(block_next[74]), .E(n774), .CK(clk), .Q(
        \block[0][74] ) );
  EDFFXL \block_reg[0][73]  ( .D(block_next[73]), .E(n774), .CK(clk), .Q(
        \block[0][73] ) );
  EDFFXL \block_reg[0][72]  ( .D(block_next[72]), .E(n774), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFXL \block_reg[0][71]  ( .D(block_next[71]), .E(n774), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFXL \block_reg[0][70]  ( .D(block_next[70]), .E(n774), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFXL \block_reg[0][69]  ( .D(block_next[69]), .E(n774), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFXL \block_reg[0][68]  ( .D(block_next[68]), .E(n774), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFXL \block_reg[0][67]  ( .D(block_next[67]), .E(n774), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFXL \block_reg[0][66]  ( .D(block_next[66]), .E(n774), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFXL \block_reg[0][65]  ( .D(block_next[65]), .E(n773), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFXL \block_reg[0][64]  ( .D(block_next[64]), .E(n773), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFX1 \block_reg[0][63]  ( .D(block_next[63]), .E(n773), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFX1 \block_reg[0][53]  ( .D(block_next[53]), .E(n773), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFX1 \block_reg[0][52]  ( .D(block_next[52]), .E(n772), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFX1 \block_reg[0][49]  ( .D(block_next[49]), .E(n772), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFX1 \block_reg[0][41]  ( .D(block_next[41]), .E(n772), .CK(clk), .Q(
        \block[0][41] ) );
  EDFFX1 \block_reg[0][38]  ( .D(block_next[38]), .E(n771), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFX1 \block_reg[0][37]  ( .D(block_next[37]), .E(n771), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFX1 \block_reg[0][36]  ( .D(block_next[36]), .E(n771), .CK(clk), .Q(
        \block[0][36] ) );
  EDFFX1 \block_reg[0][35]  ( .D(block_next[35]), .E(n771), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFX1 \block_reg[0][32]  ( .D(block_next[32]), .E(n771), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFX1 \block_reg[0][21]  ( .D(block_next[21]), .E(n770), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFX1 \block_reg[0][20]  ( .D(block_next[20]), .E(n770), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFX1 \block_reg[0][19]  ( .D(block_next[19]), .E(n770), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFX1 \block_reg[0][18]  ( .D(block_next[18]), .E(n770), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFX1 \block_reg[0][17]  ( .D(block_next[17]), .E(n770), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFX1 \block_reg[0][16]  ( .D(block_next[16]), .E(n770), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFX1 \block_reg[0][15]  ( .D(block_next[15]), .E(n770), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFX1 \block_reg[0][14]  ( .D(block_next[14]), .E(n770), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFX1 \block_reg[0][13]  ( .D(block_next[13]), .E(n769), .CK(clk), .Q(
        \block[0][13] ) );
  EDFFX1 \block_reg[0][12]  ( .D(block_next[12]), .E(n769), .CK(clk), .Q(
        \block[0][12] ) );
  EDFFX1 \block_reg[0][11]  ( .D(block_next[11]), .E(n769), .CK(clk), .Q(
        \block[0][11] ) );
  EDFFX1 \block_reg[0][10]  ( .D(block_next[10]), .E(n769), .CK(clk), .Q(
        \block[0][10] ) );
  EDFFX1 \block_reg[0][9]  ( .D(block_next[9]), .E(n769), .CK(clk), .Q(
        \block[0][9] ) );
  EDFFX1 \block_reg[0][8]  ( .D(block_next[8]), .E(n769), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFX1 \block_reg[0][7]  ( .D(block_next[7]), .E(n769), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFX1 \block_reg[0][0]  ( .D(block_next[0]), .E(n768), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFXL \block_reg[0][127]  ( .D(block_next[127]), .E(n778), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFXL \block_reg[0][126]  ( .D(block_next[126]), .E(n778), .CK(clk), .Q(
        \block[0][126] ) );
  EDFFXL \block_reg[0][125]  ( .D(block_next[125]), .E(n778), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFXL \block_reg[0][124]  ( .D(block_next[124]), .E(n778), .CK(clk), .Q(
        \block[0][124] ) );
  EDFFXL \block_reg[0][123]  ( .D(block_next[123]), .E(n778), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFXL \block_reg[0][122]  ( .D(block_next[122]), .E(n778), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFXL \block_reg[0][121]  ( .D(block_next[121]), .E(n778), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFXL \block_reg[0][120]  ( .D(block_next[120]), .E(n778), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFXL \block_reg[0][119]  ( .D(block_next[119]), .E(n778), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFXL \block_reg[0][118]  ( .D(block_next[118]), .E(n778), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFXL \block_reg[0][117]  ( .D(block_next[117]), .E(n777), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFXL \block_reg[6][116]  ( .D(block_next[116]), .E(n670), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFXL \block_reg[6][115]  ( .D(block_next[115]), .E(n670), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFXL \block_reg[6][114]  ( .D(block_next[114]), .E(n670), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFXL \block_reg[6][113]  ( .D(block_next[113]), .E(n670), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFXL \block_reg[6][112]  ( .D(block_next[112]), .E(n670), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFXL \block_reg[6][111]  ( .D(block_next[111]), .E(n670), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFXL \block_reg[6][110]  ( .D(block_next[110]), .E(n670), .CK(clk), .Q(
        \block[6][110] ) );
  EDFFXL \block_reg[6][109]  ( .D(block_next[109]), .E(n670), .CK(clk), .Q(
        \block[6][109] ) );
  EDFFXL \block_reg[6][108]  ( .D(block_next[108]), .E(n670), .CK(clk), .Q(
        \block[6][108] ) );
  EDFFXL \block_reg[6][107]  ( .D(block_next[107]), .E(n670), .CK(clk), .Q(
        \block[6][107] ) );
  EDFFXL \block_reg[6][106]  ( .D(block_next[106]), .E(n670), .CK(clk), .Q(
        \block[6][106] ) );
  EDFFXL \block_reg[6][105]  ( .D(block_next[105]), .E(n670), .CK(clk), .Q(
        \block[6][105] ) );
  EDFFXL \block_reg[6][104]  ( .D(block_next[104]), .E(n669), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFXL \block_reg[6][103]  ( .D(block_next[103]), .E(n669), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFXL \block_reg[6][102]  ( .D(block_next[102]), .E(n669), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFXL \block_reg[6][101]  ( .D(block_next[101]), .E(n669), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFXL \block_reg[6][100]  ( .D(block_next[100]), .E(n669), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFXL \block_reg[6][99]  ( .D(block_next[99]), .E(n669), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFXL \block_reg[6][98]  ( .D(block_next[98]), .E(n669), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFXL \block_reg[6][97]  ( .D(block_next[97]), .E(n669), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFXL \block_reg[6][96]  ( .D(block_next[96]), .E(n669), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFXL \block_reg[6][95]  ( .D(block_next[95]), .E(n669), .CK(clk), .Q(
        \block[6][95] ) );
  EDFFXL \block_reg[6][94]  ( .D(block_next[94]), .E(n669), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFXL \block_reg[6][93]  ( .D(block_next[93]), .E(n669), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFXL \block_reg[6][92]  ( .D(block_next[92]), .E(n669), .CK(clk), .Q(
        \block[6][92] ) );
  EDFFXL \block_reg[6][91]  ( .D(block_next[91]), .E(n668), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFXL \block_reg[6][90]  ( .D(block_next[90]), .E(n668), .CK(clk), .Q(
        \block[6][90] ) );
  EDFFXL \block_reg[6][89]  ( .D(block_next[89]), .E(n668), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFXL \block_reg[6][88]  ( .D(block_next[88]), .E(n668), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFXL \block_reg[6][87]  ( .D(block_next[87]), .E(n668), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFXL \block_reg[6][86]  ( .D(block_next[86]), .E(n668), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFXL \block_reg[6][85]  ( .D(block_next[85]), .E(n668), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFXL \block_reg[6][84]  ( .D(block_next[84]), .E(n668), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFXL \block_reg[6][83]  ( .D(block_next[83]), .E(n668), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFXL \block_reg[6][82]  ( .D(block_next[82]), .E(n668), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFXL \block_reg[6][81]  ( .D(block_next[81]), .E(n668), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFXL \block_reg[6][80]  ( .D(block_next[80]), .E(n668), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFXL \block_reg[6][79]  ( .D(block_next[79]), .E(n668), .CK(clk), .Q(
        \block[6][79] ) );
  EDFFXL \block_reg[6][78]  ( .D(block_next[78]), .E(n667), .CK(clk), .Q(
        \block[6][78] ) );
  EDFFXL \block_reg[6][77]  ( .D(block_next[77]), .E(n667), .CK(clk), .Q(
        \block[6][77] ) );
  EDFFXL \block_reg[6][76]  ( .D(block_next[76]), .E(n667), .CK(clk), .Q(
        \block[6][76] ) );
  EDFFXL \block_reg[6][75]  ( .D(block_next[75]), .E(n667), .CK(clk), .Q(
        \block[6][75] ) );
  EDFFXL \block_reg[6][74]  ( .D(block_next[74]), .E(n667), .CK(clk), .Q(
        \block[6][74] ) );
  EDFFXL \block_reg[6][73]  ( .D(block_next[73]), .E(n667), .CK(clk), .Q(
        \block[6][73] ) );
  EDFFXL \block_reg[6][72]  ( .D(block_next[72]), .E(n667), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFXL \block_reg[6][71]  ( .D(block_next[71]), .E(n667), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFXL \block_reg[6][70]  ( .D(block_next[70]), .E(n667), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFXL \block_reg[6][69]  ( .D(block_next[69]), .E(n667), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFXL \block_reg[6][68]  ( .D(block_next[68]), .E(n667), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFXL \block_reg[6][67]  ( .D(block_next[67]), .E(n667), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFXL \block_reg[6][66]  ( .D(block_next[66]), .E(n667), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFXL \block_reg[6][65]  ( .D(block_next[65]), .E(n666), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFXL \block_reg[6][64]  ( .D(block_next[64]), .E(n666), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFX1 \block_reg[6][53]  ( .D(block_next[53]), .E(n666), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFX1 \block_reg[6][52]  ( .D(block_next[52]), .E(n665), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFX1 \block_reg[6][41]  ( .D(block_next[41]), .E(n665), .CK(clk), .Q(
        \block[6][41] ) );
  EDFFX1 \block_reg[6][38]  ( .D(block_next[38]), .E(n664), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFX1 \block_reg[6][37]  ( .D(block_next[37]), .E(n664), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFX1 \block_reg[6][36]  ( .D(block_next[36]), .E(n664), .CK(clk), .Q(
        \block[6][36] ) );
  EDFFX1 \block_reg[6][35]  ( .D(block_next[35]), .E(n664), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFX1 \block_reg[6][32]  ( .D(block_next[32]), .E(n664), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFX1 \block_reg[6][20]  ( .D(block_next[20]), .E(n663), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFX1 \block_reg[6][19]  ( .D(block_next[19]), .E(n663), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFX1 \block_reg[6][18]  ( .D(block_next[18]), .E(n663), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFX1 \block_reg[6][17]  ( .D(block_next[17]), .E(n663), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFX1 \block_reg[6][16]  ( .D(block_next[16]), .E(n663), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFX1 \block_reg[6][15]  ( .D(block_next[15]), .E(n663), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFX1 \block_reg[6][14]  ( .D(block_next[14]), .E(n663), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFX1 \block_reg[6][13]  ( .D(block_next[13]), .E(n662), .CK(clk), .Q(
        \block[6][13] ) );
  EDFFX1 \block_reg[6][12]  ( .D(block_next[12]), .E(n662), .CK(clk), .Q(
        \block[6][12] ) );
  EDFFX1 \block_reg[6][11]  ( .D(block_next[11]), .E(n662), .CK(clk), .Q(
        \block[6][11] ) );
  EDFFX1 \block_reg[6][10]  ( .D(block_next[10]), .E(n662), .CK(clk), .Q(
        \block[6][10] ) );
  EDFFX1 \block_reg[6][9]  ( .D(block_next[9]), .E(n662), .CK(clk), .Q(
        \block[6][9] ) );
  EDFFX1 \block_reg[6][8]  ( .D(block_next[8]), .E(n662), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFX1 \block_reg[6][0]  ( .D(block_next[0]), .E(n661), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFXL \block_reg[6][127]  ( .D(block_next[127]), .E(n671), .CK(clk), .Q(
        \block[6][127] ) );
  EDFFXL \block_reg[6][126]  ( .D(block_next[126]), .E(n671), .CK(clk), .Q(
        \block[6][126] ) );
  EDFFXL \block_reg[6][125]  ( .D(block_next[125]), .E(n671), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFXL \block_reg[6][124]  ( .D(block_next[124]), .E(n671), .CK(clk), .Q(
        \block[6][124] ) );
  EDFFXL \block_reg[6][123]  ( .D(block_next[123]), .E(n671), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFXL \block_reg[6][122]  ( .D(block_next[122]), .E(n671), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFXL \block_reg[6][121]  ( .D(block_next[121]), .E(n671), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFXL \block_reg[6][120]  ( .D(block_next[120]), .E(n671), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFXL \block_reg[6][119]  ( .D(block_next[119]), .E(n671), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFXL \block_reg[6][118]  ( .D(block_next[118]), .E(n671), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFXL \block_reg[6][117]  ( .D(block_next[117]), .E(n670), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFXL \block_reg[2][116]  ( .D(block_next[116]), .E(n741), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFXL \block_reg[2][115]  ( .D(block_next[115]), .E(n741), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFXL \block_reg[2][114]  ( .D(block_next[114]), .E(n741), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFXL \block_reg[2][113]  ( .D(block_next[113]), .E(n741), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFXL \block_reg[2][112]  ( .D(block_next[112]), .E(n741), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFXL \block_reg[2][111]  ( .D(block_next[111]), .E(n741), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFXL \block_reg[2][110]  ( .D(block_next[110]), .E(n741), .CK(clk), .Q(
        \block[2][110] ) );
  EDFFXL \block_reg[2][109]  ( .D(block_next[109]), .E(n741), .CK(clk), .Q(
        \block[2][109] ) );
  EDFFXL \block_reg[2][108]  ( .D(block_next[108]), .E(n741), .CK(clk), .Q(
        \block[2][108] ) );
  EDFFXL \block_reg[2][107]  ( .D(block_next[107]), .E(n741), .CK(clk), .Q(
        \block[2][107] ) );
  EDFFXL \block_reg[2][106]  ( .D(block_next[106]), .E(n741), .CK(clk), .Q(
        \block[2][106] ) );
  EDFFXL \block_reg[2][105]  ( .D(block_next[105]), .E(n741), .CK(clk), .Q(
        \block[2][105] ) );
  EDFFXL \block_reg[2][104]  ( .D(block_next[104]), .E(n740), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFXL \block_reg[2][103]  ( .D(block_next[103]), .E(n740), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFXL \block_reg[2][102]  ( .D(block_next[102]), .E(n740), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFXL \block_reg[2][101]  ( .D(block_next[101]), .E(n740), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFXL \block_reg[2][100]  ( .D(block_next[100]), .E(n740), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFXL \block_reg[2][99]  ( .D(block_next[99]), .E(n740), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFXL \block_reg[2][98]  ( .D(block_next[98]), .E(n740), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFXL \block_reg[2][97]  ( .D(block_next[97]), .E(n740), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFXL \block_reg[2][96]  ( .D(block_next[96]), .E(n740), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFXL \block_reg[2][95]  ( .D(block_next[95]), .E(n740), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFXL \block_reg[2][94]  ( .D(block_next[94]), .E(n740), .CK(clk), .Q(
        \block[2][94] ) );
  EDFFXL \block_reg[2][93]  ( .D(block_next[93]), .E(n740), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFXL \block_reg[2][92]  ( .D(block_next[92]), .E(n740), .CK(clk), .Q(
        \block[2][92] ) );
  EDFFXL \block_reg[2][91]  ( .D(block_next[91]), .E(n739), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFXL \block_reg[2][90]  ( .D(block_next[90]), .E(n739), .CK(clk), .Q(
        \block[2][90] ) );
  EDFFXL \block_reg[2][89]  ( .D(block_next[89]), .E(n739), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFXL \block_reg[2][88]  ( .D(block_next[88]), .E(n739), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFXL \block_reg[2][87]  ( .D(block_next[87]), .E(n739), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFXL \block_reg[2][86]  ( .D(block_next[86]), .E(n739), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFXL \block_reg[2][85]  ( .D(block_next[85]), .E(n739), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFXL \block_reg[2][84]  ( .D(block_next[84]), .E(n739), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFXL \block_reg[2][83]  ( .D(block_next[83]), .E(n739), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFXL \block_reg[2][82]  ( .D(block_next[82]), .E(n739), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFXL \block_reg[2][81]  ( .D(block_next[81]), .E(n739), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFXL \block_reg[2][80]  ( .D(block_next[80]), .E(n739), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFXL \block_reg[2][79]  ( .D(block_next[79]), .E(n739), .CK(clk), .Q(
        \block[2][79] ) );
  EDFFXL \block_reg[2][78]  ( .D(block_next[78]), .E(n738), .CK(clk), .Q(
        \block[2][78] ) );
  EDFFXL \block_reg[2][77]  ( .D(block_next[77]), .E(n738), .CK(clk), .Q(
        \block[2][77] ) );
  EDFFXL \block_reg[2][76]  ( .D(block_next[76]), .E(n738), .CK(clk), .Q(
        \block[2][76] ) );
  EDFFXL \block_reg[2][75]  ( .D(block_next[75]), .E(n738), .CK(clk), .Q(
        \block[2][75] ) );
  EDFFXL \block_reg[2][74]  ( .D(block_next[74]), .E(n738), .CK(clk), .Q(
        \block[2][74] ) );
  EDFFXL \block_reg[2][73]  ( .D(block_next[73]), .E(n738), .CK(clk), .Q(
        \block[2][73] ) );
  EDFFXL \block_reg[2][72]  ( .D(block_next[72]), .E(n738), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFXL \block_reg[2][71]  ( .D(block_next[71]), .E(n738), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFXL \block_reg[2][70]  ( .D(block_next[70]), .E(n738), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFXL \block_reg[2][69]  ( .D(block_next[69]), .E(n738), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFXL \block_reg[2][68]  ( .D(block_next[68]), .E(n738), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFXL \block_reg[2][67]  ( .D(block_next[67]), .E(n738), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFXL \block_reg[2][66]  ( .D(block_next[66]), .E(n738), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFXL \block_reg[2][65]  ( .D(block_next[65]), .E(n737), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFXL \block_reg[2][64]  ( .D(block_next[64]), .E(n737), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFXL \block_reg[2][63]  ( .D(block_next[63]), .E(n737), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFXL \block_reg[2][62]  ( .D(block_next[62]), .E(n737), .CK(clk), .Q(
        \block[2][62] ) );
  EDFFXL \block_reg[2][61]  ( .D(block_next[61]), .E(n737), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFXL \block_reg[2][60]  ( .D(block_next[60]), .E(n737), .CK(clk), .Q(
        \block[2][60] ) );
  EDFFXL \block_reg[2][59]  ( .D(block_next[59]), .E(n737), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFXL \block_reg[2][58]  ( .D(block_next[58]), .E(n737), .CK(clk), .Q(
        \block[2][58] ) );
  EDFFXL \block_reg[2][57]  ( .D(block_next[57]), .E(n737), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFXL \block_reg[2][56]  ( .D(block_next[56]), .E(n737), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFXL \block_reg[2][55]  ( .D(block_next[55]), .E(n737), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFXL \block_reg[2][54]  ( .D(block_next[54]), .E(n737), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFXL \block_reg[2][53]  ( .D(block_next[53]), .E(n737), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFXL \block_reg[2][52]  ( .D(block_next[52]), .E(n736), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFXL \block_reg[2][51]  ( .D(block_next[51]), .E(n736), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFXL \block_reg[2][50]  ( .D(block_next[50]), .E(n736), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFXL \block_reg[2][49]  ( .D(block_next[49]), .E(n736), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFXL \block_reg[2][48]  ( .D(block_next[48]), .E(n736), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFXL \block_reg[2][47]  ( .D(block_next[47]), .E(n736), .CK(clk), .Q(
        \block[2][47] ) );
  EDFFXL \block_reg[2][46]  ( .D(block_next[46]), .E(n736), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFXL \block_reg[2][45]  ( .D(block_next[45]), .E(n736), .CK(clk), .Q(
        \block[2][45] ) );
  EDFFXL \block_reg[2][44]  ( .D(block_next[44]), .E(n736), .CK(clk), .Q(
        \block[2][44] ) );
  EDFFXL \block_reg[2][43]  ( .D(block_next[43]), .E(n736), .CK(clk), .Q(
        \block[2][43] ) );
  EDFFXL \block_reg[2][42]  ( .D(block_next[42]), .E(n736), .CK(clk), .Q(
        \block[2][42] ) );
  EDFFXL \block_reg[2][41]  ( .D(block_next[41]), .E(n736), .CK(clk), .Q(
        \block[2][41] ) );
  EDFFXL \block_reg[2][40]  ( .D(block_next[40]), .E(n736), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFXL \block_reg[2][39]  ( .D(block_next[39]), .E(n735), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFXL \block_reg[2][38]  ( .D(block_next[38]), .E(n735), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFXL \block_reg[2][37]  ( .D(block_next[37]), .E(n735), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFXL \block_reg[2][36]  ( .D(block_next[36]), .E(n735), .CK(clk), .Q(
        \block[2][36] ) );
  EDFFXL \block_reg[2][35]  ( .D(block_next[35]), .E(n735), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFXL \block_reg[2][34]  ( .D(block_next[34]), .E(n735), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFXL \block_reg[2][33]  ( .D(block_next[33]), .E(n735), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFXL \block_reg[2][32]  ( .D(block_next[32]), .E(n735), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFXL \block_reg[2][31]  ( .D(block_next[31]), .E(n735), .CK(clk), .Q(
        \block[2][31] ) );
  EDFFXL \block_reg[2][30]  ( .D(block_next[30]), .E(n735), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFXL \block_reg[2][29]  ( .D(block_next[29]), .E(n735), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFXL \block_reg[2][28]  ( .D(block_next[28]), .E(n735), .CK(clk), .Q(
        \block[2][28] ) );
  EDFFXL \block_reg[2][27]  ( .D(block_next[27]), .E(n735), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFXL \block_reg[2][26]  ( .D(block_next[26]), .E(n734), .CK(clk), .Q(
        \block[2][26] ) );
  EDFFXL \block_reg[2][25]  ( .D(block_next[25]), .E(n734), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFXL \block_reg[2][24]  ( .D(block_next[24]), .E(n734), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFXL \block_reg[2][23]  ( .D(block_next[23]), .E(n734), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFXL \block_reg[2][22]  ( .D(block_next[22]), .E(n734), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFXL \block_reg[2][21]  ( .D(block_next[21]), .E(n734), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFXL \block_reg[2][20]  ( .D(block_next[20]), .E(n734), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFXL \block_reg[2][19]  ( .D(block_next[19]), .E(n734), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFXL \block_reg[2][18]  ( .D(block_next[18]), .E(n734), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFXL \block_reg[2][17]  ( .D(block_next[17]), .E(n734), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFXL \block_reg[2][16]  ( .D(block_next[16]), .E(n734), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFXL \block_reg[2][15]  ( .D(block_next[15]), .E(n734), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFXL \block_reg[2][14]  ( .D(block_next[14]), .E(n734), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFXL \block_reg[2][13]  ( .D(block_next[13]), .E(n733), .CK(clk), .Q(
        \block[2][13] ) );
  EDFFXL \block_reg[2][12]  ( .D(block_next[12]), .E(n733), .CK(clk), .Q(
        \block[2][12] ) );
  EDFFXL \block_reg[2][11]  ( .D(block_next[11]), .E(n733), .CK(clk), .Q(
        \block[2][11] ) );
  EDFFXL \block_reg[2][10]  ( .D(block_next[10]), .E(n733), .CK(clk), .Q(
        \block[2][10] ) );
  EDFFXL \block_reg[2][9]  ( .D(block_next[9]), .E(n733), .CK(clk), .Q(
        \block[2][9] ) );
  EDFFXL \block_reg[2][8]  ( .D(block_next[8]), .E(n733), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFXL \block_reg[2][7]  ( .D(block_next[7]), .E(n733), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFXL \block_reg[2][6]  ( .D(block_next[6]), .E(n733), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFXL \block_reg[2][5]  ( .D(block_next[5]), .E(n733), .CK(clk), .QN(n132)
         );
  EDFFXL \block_reg[2][4]  ( .D(block_next[4]), .E(n733), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFXL \block_reg[2][3]  ( .D(block_next[3]), .E(n733), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFXL \block_reg[2][2]  ( .D(block_next[2]), .E(n733), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFXL \block_reg[2][1]  ( .D(block_next[1]), .E(n733), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFXL \block_reg[2][0]  ( .D(block_next[0]), .E(n732), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFXL \block_reg[2][127]  ( .D(block_next[127]), .E(n742), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFXL \block_reg[2][126]  ( .D(block_next[126]), .E(n742), .CK(clk), .Q(
        \block[2][126] ) );
  EDFFXL \block_reg[2][125]  ( .D(block_next[125]), .E(n742), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFXL \block_reg[2][124]  ( .D(block_next[124]), .E(n742), .CK(clk), .Q(
        \block[2][124] ) );
  EDFFXL \block_reg[2][123]  ( .D(block_next[123]), .E(n742), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFXL \block_reg[2][122]  ( .D(block_next[122]), .E(n742), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFXL \block_reg[2][121]  ( .D(block_next[121]), .E(n742), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFXL \block_reg[2][120]  ( .D(block_next[120]), .E(n742), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFXL \block_reg[2][119]  ( .D(block_next[119]), .E(n742), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFXL \block_reg[2][118]  ( .D(block_next[118]), .E(n742), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFXL \block_reg[2][117]  ( .D(block_next[117]), .E(n741), .CK(clk), .Q(
        \block[2][117] ) );
  DFFRX1 \blockvalid_reg[7]  ( .D(n503), .CK(clk), .RN(n792), .Q(blockvalid[7]), .QN(n486) );
  DFFRX1 \blockvalid_reg[3]  ( .D(n498), .CK(clk), .RN(n791), .Q(blockvalid[3]), .QN(n482) );
  DFFRX1 \blockvalid_reg[5]  ( .D(n500), .CK(clk), .RN(n791), .Q(blockvalid[5]), .QN(n484) );
  DFFRX1 \blockvalid_reg[1]  ( .D(n496), .CK(clk), .RN(n791), .Q(blockvalid[1]), .QN(n480) );
  DFFRX1 \blockvalid_reg[4]  ( .D(n499), .CK(clk), .RN(n791), .Q(blockvalid[4]), .QN(n483) );
  DFFRX1 \blockvalid_reg[0]  ( .D(n495), .CK(clk), .RN(n791), .Q(blockvalid[0]), .QN(n479) );
  DFFRX1 \blockvalid_reg[6]  ( .D(n501), .CK(clk), .RN(n792), .Q(blockvalid[6]), .QN(n485) );
  DFFRX1 \blockvalid_reg[2]  ( .D(n497), .CK(clk), .RN(n791), .Q(blockvalid[2]), .QN(n481) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][18] ) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][18] ) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(blocktag_next[17]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][17] ) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(blocktag_next[17]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][17] ) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(blocktag_next[0]), .E(n714), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(blocktag_next[0]), .E(n641), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(blocktag_next[14]), .E(n715), .CK(clk), 
        .QN(n109) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(blocktag_next[23]), .E(n715), .CK(clk), 
        .QN(n93) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(blocktag_next[14]), .E(n642), .CK(clk), 
        .QN(n113) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n715), .CK(clk), 
        .QN(n101) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(blocktag_next[23]), .E(n642), .CK(clk), 
        .QN(n97) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n642), .CK(clk), 
        .QN(n105) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n715), .CK(clk), 
        .QN(n117) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n642), .CK(clk), 
        .QN(n121) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][21] ) );
  EDFFX1 \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][21] ) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(n2), .E(n714), .CK(clk), .Q(
        \blocktag[3][5] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(n2), .E(n641), .CK(clk), .Q(
        \blocktag[7][5] ) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][16] ) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][16] ) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][20] ) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(blocktag_next[10]), .E(n714), .CK(clk), 
        .QN(n125) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(blocktag_next[10]), .E(n641), .CK(clk), 
        .QN(n129) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n714), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n641), .CK(clk), 
        .Q(\blocktag[7][11] ) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n715), .CK(clk), 
        .QN(n77) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n642), .CK(clk), 
        .QN(n81) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n714), .CK(clk), .QN(
        n61) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n641), .CK(clk), .QN(
        n65) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(blocktag_next[12]), .E(n714), .CK(clk), 
        .QN(n85) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(blocktag_next[12]), .E(n641), .CK(clk), 
        .QN(n89) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n714), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n641), .CK(clk), .Q(
        \blocktag[7][1] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n714), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n641), .CK(clk), .Q(
        \blocktag[7][2] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(n714), .CK(clk), .Q(
        \blocktag[3][8] ) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(n641), .CK(clk), .Q(
        \blocktag[7][8] ) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][13] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(blocktag_next[7]), .E(n714), .CK(clk), .Q(
        \blocktag[3][7] ) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(blocktag_next[7]), .E(n641), .CK(clk), .Q(
        \blocktag[7][7] ) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(n715), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(n642), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(n714), .CK(clk), .Q(
        \blocktag[3][6] ) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(n641), .CK(clk), .Q(
        \blocktag[7][6] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(n714), .CK(clk), .QN(
        n69) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(n641), .CK(clk), .QN(
        n73) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][18] ) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][18] ) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(blocktag_next[17]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][17] ) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(blocktag_next[17]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][17] ) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(blocktag_next[0]), .E(n748), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(blocktag_next[0]), .E(n679), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(blocktag_next[14]), .E(n749), .CK(clk), 
        .QN(n107) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(blocktag_next[23]), .E(n749), .CK(clk), 
        .QN(n91) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(blocktag_next[14]), .E(n680), .CK(clk), 
        .QN(n111) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n749), .CK(clk), 
        .QN(n99) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(blocktag_next[23]), .E(n680), .CK(clk), 
        .QN(n95) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n680), .CK(clk), 
        .QN(n103) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n749), .CK(clk), 
        .QN(n115) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n680), .CK(clk), 
        .QN(n119) );
  EDFFX1 \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][21] ) );
  EDFFX1 \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][21] ) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(n2), .E(n748), .CK(clk), .Q(
        \blocktag[1][5] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(n2), .E(n679), .CK(clk), .Q(
        \blocktag[5][5] ) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][16] ) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][16] ) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][20] ) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(blocktag_next[10]), .E(n748), .CK(clk), 
        .QN(n123) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(blocktag_next[10]), .E(n679), .CK(clk), 
        .QN(n127) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n748), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n679), .CK(clk), 
        .Q(\blocktag[5][11] ) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n749), .CK(clk), 
        .QN(n75) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n680), .CK(clk), 
        .QN(n79) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n748), .CK(clk), .QN(
        n59) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n679), .CK(clk), .QN(
        n63) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(blocktag_next[12]), .E(n748), .CK(clk), 
        .QN(n83) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(blocktag_next[12]), .E(n679), .CK(clk), 
        .QN(n87) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n748), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n679), .CK(clk), .Q(
        \blocktag[5][1] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n748), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n679), .CK(clk), .Q(
        \blocktag[5][2] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(n748), .CK(clk), .Q(
        \blocktag[1][8] ) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n679), .CK(clk), .Q(
        \blocktag[5][8] ) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][13] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(blocktag_next[7]), .E(n748), .CK(clk), .Q(
        \blocktag[1][7] ) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(blocktag_next[7]), .E(n679), .CK(clk), .Q(
        \blocktag[5][7] ) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n749), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(n680), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(n748), .CK(clk), .Q(
        \blocktag[1][6] ) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n679), .CK(clk), .Q(
        \blocktag[5][6] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(n748), .CK(clk), .QN(
        n67) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n679), .CK(clk), .QN(
        n71) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][18] ) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][18] ) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(blocktag_next[17]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][17] ) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(blocktag_next[17]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][17] ) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(blocktag_next[0]), .E(n767), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(blocktag_next[0]), .E(n696), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(blocktag_next[14]), .E(n768), .CK(clk), 
        .QN(n106) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(blocktag_next[23]), .E(n768), .CK(clk), 
        .QN(n90) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(blocktag_next[14]), .E(n697), .CK(clk), 
        .QN(n110) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n768), .CK(clk), 
        .QN(n98) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(blocktag_next[23]), .E(n697), .CK(clk), 
        .QN(n94) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n697), .CK(clk), 
        .QN(n102) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n768), .CK(clk), 
        .QN(n114) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n697), .CK(clk), 
        .QN(n118) );
  EDFFX1 \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][21] ) );
  EDFFX1 \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][21] ) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(n2), .E(n767), .CK(clk), .Q(
        \blocktag[0][5] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(n2), .E(n696), .CK(clk), .Q(
        \blocktag[4][5] ) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][16] ) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][16] ) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][20] ) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(blocktag_next[10]), .E(n767), .CK(clk), 
        .QN(n122) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(blocktag_next[10]), .E(n696), .CK(clk), 
        .QN(n126) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n767), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n696), .CK(clk), 
        .Q(\blocktag[4][11] ) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n768), .CK(clk), 
        .QN(n74) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n697), .CK(clk), 
        .QN(n78) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n767), .CK(clk), .QN(
        n58) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n696), .CK(clk), .QN(
        n62) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(blocktag_next[12]), .E(n767), .CK(clk), 
        .QN(n82) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(blocktag_next[12]), .E(n696), .CK(clk), 
        .QN(n86) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n767), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n696), .CK(clk), .Q(
        \blocktag[4][1] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n767), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n696), .CK(clk), .Q(
        \blocktag[4][2] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n767), .CK(clk), .Q(
        \blocktag[0][8] ) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n696), .CK(clk), .Q(
        \blocktag[4][8] ) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][13] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(blocktag_next[7]), .E(n767), .CK(clk), .Q(
        \blocktag[0][7] ) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(blocktag_next[7]), .E(n696), .CK(clk), .Q(
        \blocktag[4][7] ) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(n768), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(n697), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n767), .CK(clk), .Q(
        \blocktag[0][6] ) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n696), .CK(clk), .Q(
        \blocktag[4][6] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n767), .CK(clk), .QN(
        n66) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n696), .CK(clk), .QN(
        n70) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][18] ) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][18] ) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(blocktag_next[17]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][17] ) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(blocktag_next[17]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][17] ) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(blocktag_next[0]), .E(n731), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(blocktag_next[0]), .E(n660), .CK(clk), .Q(
        \blocktag[6][0] ) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(blocktag_next[14]), .E(n732), .CK(clk), 
        .QN(n108) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(blocktag_next[23]), .E(n732), .CK(clk), 
        .QN(n92) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(blocktag_next[14]), .E(n661), .CK(clk), 
        .QN(n112) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n732), .CK(clk), 
        .QN(n100) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(blocktag_next[23]), .E(n661), .CK(clk), 
        .QN(n96) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n661), .CK(clk), 
        .QN(n104) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n732), .CK(clk), 
        .QN(n116) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n661), .CK(clk), 
        .QN(n120) );
  EDFFX1 \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][21] ) );
  EDFFX1 \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][21] ) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(n2), .E(n731), .CK(clk), .Q(
        \blocktag[2][5] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(n2), .E(n660), .CK(clk), .Q(
        \blocktag[6][5] ) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][16] ) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][16] ) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][20] ) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(blocktag_next[10]), .E(n731), .CK(clk), 
        .QN(n124) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(blocktag_next[10]), .E(n660), .CK(clk), 
        .QN(n128) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n731), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n660), .CK(clk), 
        .Q(\blocktag[6][11] ) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n732), .CK(clk), 
        .QN(n76) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n661), .CK(clk), 
        .QN(n80) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n731), .CK(clk), .QN(
        n60) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n660), .CK(clk), .QN(
        n64) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(blocktag_next[12]), .E(n731), .CK(clk), 
        .QN(n84) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(blocktag_next[12]), .E(n660), .CK(clk), 
        .QN(n88) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n731), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n660), .CK(clk), .Q(
        \blocktag[6][1] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n731), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n660), .CK(clk), .Q(
        \blocktag[6][2] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n731), .CK(clk), .Q(
        \blocktag[2][8] ) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n660), .CK(clk), .Q(
        \blocktag[6][8] ) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][13] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(blocktag_next[7]), .E(n731), .CK(clk), .Q(
        \blocktag[2][7] ) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(blocktag_next[7]), .E(n660), .CK(clk), .Q(
        \blocktag[6][7] ) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(n732), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n661), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n731), .CK(clk), .Q(
        \blocktag[2][6] ) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n660), .CK(clk), .Q(
        \blocktag[6][6] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n731), .CK(clk), .QN(
        n68) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n660), .CK(clk), .QN(
        n72) );
  EDFFXL \block_reg[6][40]  ( .D(block_next[40]), .E(n665), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFXL \block_reg[0][40]  ( .D(block_next[40]), .E(n772), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFXL \block_reg[4][40]  ( .D(block_next[40]), .E(n701), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFXL \block_reg[1][40]  ( .D(block_next[40]), .E(n753), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFXL \block_reg[5][40]  ( .D(block_next[40]), .E(n684), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFXL \block_reg[3][40]  ( .D(block_next[40]), .E(n719), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFXL \block_reg[7][40]  ( .D(block_next[40]), .E(n646), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFXL \block_reg[6][22]  ( .D(block_next[22]), .E(n663), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFXL \block_reg[0][22]  ( .D(block_next[22]), .E(n770), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFXL \block_reg[4][22]  ( .D(block_next[22]), .E(n699), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFXL \block_reg[1][22]  ( .D(block_next[22]), .E(n751), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFXL \block_reg[5][22]  ( .D(block_next[22]), .E(n682), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFXL \block_reg[3][22]  ( .D(block_next[22]), .E(n717), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFXL \block_reg[7][22]  ( .D(block_next[22]), .E(n644), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFXL \block_reg[6][23]  ( .D(block_next[23]), .E(n663), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFXL \block_reg[0][23]  ( .D(block_next[23]), .E(n770), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFXL \block_reg[4][23]  ( .D(block_next[23]), .E(n699), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFXL \block_reg[1][23]  ( .D(block_next[23]), .E(n751), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFXL \block_reg[5][23]  ( .D(block_next[23]), .E(n682), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFXL \block_reg[3][23]  ( .D(block_next[23]), .E(n717), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFXL \block_reg[7][23]  ( .D(block_next[23]), .E(n644), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFXL \block_reg[6][24]  ( .D(block_next[24]), .E(n663), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFXL \block_reg[0][24]  ( .D(block_next[24]), .E(n770), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFXL \block_reg[4][24]  ( .D(block_next[24]), .E(n699), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFXL \block_reg[1][24]  ( .D(block_next[24]), .E(n751), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFXL \block_reg[5][24]  ( .D(block_next[24]), .E(n682), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFXL \block_reg[3][24]  ( .D(block_next[24]), .E(n717), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFXL \block_reg[7][24]  ( .D(block_next[24]), .E(n644), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFXL \block_reg[6][25]  ( .D(block_next[25]), .E(n663), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFXL \block_reg[0][25]  ( .D(block_next[25]), .E(n770), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFXL \block_reg[4][25]  ( .D(block_next[25]), .E(n699), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFXL \block_reg[1][25]  ( .D(block_next[25]), .E(n751), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFXL \block_reg[5][25]  ( .D(block_next[25]), .E(n682), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFXL \block_reg[3][25]  ( .D(block_next[25]), .E(n717), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFXL \block_reg[7][25]  ( .D(block_next[25]), .E(n644), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFXL \block_reg[6][26]  ( .D(block_next[26]), .E(n663), .CK(clk), .Q(
        \block[6][26] ) );
  EDFFXL \block_reg[0][26]  ( .D(block_next[26]), .E(n770), .CK(clk), .Q(
        \block[0][26] ) );
  EDFFXL \block_reg[4][26]  ( .D(block_next[26]), .E(n699), .CK(clk), .Q(
        \block[4][26] ) );
  EDFFXL \block_reg[1][26]  ( .D(block_next[26]), .E(n751), .CK(clk), .Q(
        \block[1][26] ) );
  EDFFXL \block_reg[5][26]  ( .D(block_next[26]), .E(n682), .CK(clk), .Q(
        \block[5][26] ) );
  EDFFXL \block_reg[3][26]  ( .D(block_next[26]), .E(n717), .CK(clk), .Q(
        \block[3][26] ) );
  EDFFXL \block_reg[7][26]  ( .D(block_next[26]), .E(n644), .CK(clk), .Q(
        \block[7][26] ) );
  EDFFXL \block_reg[6][29]  ( .D(block_next[29]), .E(n664), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFXL \block_reg[0][29]  ( .D(block_next[29]), .E(n771), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFXL \block_reg[4][29]  ( .D(block_next[29]), .E(n700), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFXL \block_reg[1][29]  ( .D(block_next[29]), .E(n752), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFXL \block_reg[5][29]  ( .D(block_next[29]), .E(n683), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFXL \block_reg[3][29]  ( .D(block_next[29]), .E(n718), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFXL \block_reg[7][29]  ( .D(block_next[29]), .E(n645), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFXL \block_reg[6][30]  ( .D(block_next[30]), .E(n664), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFXL \block_reg[0][30]  ( .D(block_next[30]), .E(n771), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFXL \block_reg[4][30]  ( .D(block_next[30]), .E(n700), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFXL \block_reg[1][30]  ( .D(block_next[30]), .E(n752), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFXL \block_reg[5][30]  ( .D(block_next[30]), .E(n683), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFXL \block_reg[3][30]  ( .D(block_next[30]), .E(n718), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFXL \block_reg[7][30]  ( .D(block_next[30]), .E(n645), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFXL \block_reg[6][31]  ( .D(block_next[31]), .E(n664), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFXL \block_reg[0][31]  ( .D(block_next[31]), .E(n771), .CK(clk), .Q(
        \block[0][31] ) );
  EDFFXL \block_reg[4][31]  ( .D(block_next[31]), .E(n700), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFXL \block_reg[1][31]  ( .D(block_next[31]), .E(n752), .CK(clk), .Q(
        \block[1][31] ) );
  EDFFXL \block_reg[5][31]  ( .D(block_next[31]), .E(n683), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFXL \block_reg[3][31]  ( .D(block_next[31]), .E(n718), .CK(clk), .Q(
        \block[3][31] ) );
  EDFFXL \block_reg[7][31]  ( .D(block_next[31]), .E(n645), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFXL \block_reg[6][27]  ( .D(block_next[27]), .E(n664), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFXL \block_reg[0][27]  ( .D(block_next[27]), .E(n771), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFXL \block_reg[4][27]  ( .D(block_next[27]), .E(n700), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFXL \block_reg[1][27]  ( .D(block_next[27]), .E(n752), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFXL \block_reg[5][27]  ( .D(block_next[27]), .E(n683), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFXL \block_reg[3][27]  ( .D(block_next[27]), .E(n718), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFXL \block_reg[7][27]  ( .D(block_next[27]), .E(n645), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFXL \block_reg[6][28]  ( .D(block_next[28]), .E(n664), .CK(clk), .Q(
        \block[6][28] ) );
  EDFFXL \block_reg[0][28]  ( .D(block_next[28]), .E(n771), .CK(clk), .Q(
        \block[0][28] ) );
  EDFFXL \block_reg[4][28]  ( .D(block_next[28]), .E(n700), .CK(clk), .Q(
        \block[4][28] ) );
  EDFFXL \block_reg[1][28]  ( .D(block_next[28]), .E(n752), .CK(clk), .Q(
        \block[1][28] ) );
  EDFFXL \block_reg[5][28]  ( .D(block_next[28]), .E(n683), .CK(clk), .Q(
        \block[5][28] ) );
  EDFFXL \block_reg[3][28]  ( .D(block_next[28]), .E(n718), .CK(clk), .Q(
        \block[3][28] ) );
  EDFFXL \block_reg[7][28]  ( .D(block_next[28]), .E(n645), .CK(clk), .Q(
        \block[7][28] ) );
  EDFFXL \block_reg[6][39]  ( .D(block_next[39]), .E(n664), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFXL \block_reg[0][39]  ( .D(block_next[39]), .E(n771), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFXL \block_reg[4][39]  ( .D(block_next[39]), .E(n700), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFXL \block_reg[1][39]  ( .D(block_next[39]), .E(n752), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFXL \block_reg[5][39]  ( .D(block_next[39]), .E(n683), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFXL \block_reg[3][39]  ( .D(block_next[39]), .E(n718), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFXL \block_reg[7][39]  ( .D(block_next[39]), .E(n645), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFXL \block_reg[6][33]  ( .D(block_next[33]), .E(n664), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFXL \block_reg[0][33]  ( .D(block_next[33]), .E(n771), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFXL \block_reg[4][33]  ( .D(block_next[33]), .E(n700), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFXL \block_reg[1][33]  ( .D(block_next[33]), .E(n752), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFXL \block_reg[5][33]  ( .D(block_next[33]), .E(n683), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFXL \block_reg[3][33]  ( .D(block_next[33]), .E(n718), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFXL \block_reg[7][33]  ( .D(block_next[33]), .E(n645), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFXL \block_reg[6][34]  ( .D(block_next[34]), .E(n664), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFXL \block_reg[0][34]  ( .D(block_next[34]), .E(n771), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFXL \block_reg[4][34]  ( .D(block_next[34]), .E(n700), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFXL \block_reg[1][34]  ( .D(block_next[34]), .E(n752), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFXL \block_reg[5][34]  ( .D(block_next[34]), .E(n683), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFXL \block_reg[6][42]  ( .D(block_next[42]), .E(n665), .CK(clk), .Q(
        \block[6][42] ) );
  EDFFXL \block_reg[0][42]  ( .D(block_next[42]), .E(n772), .CK(clk), .Q(
        \block[0][42] ) );
  EDFFXL \block_reg[4][42]  ( .D(block_next[42]), .E(n701), .CK(clk), .Q(
        \block[4][42] ) );
  EDFFXL \block_reg[1][42]  ( .D(block_next[42]), .E(n753), .CK(clk), .Q(
        \block[1][42] ) );
  EDFFXL \block_reg[5][42]  ( .D(block_next[42]), .E(n684), .CK(clk), .Q(
        \block[5][42] ) );
  EDFFXL \block_reg[3][42]  ( .D(block_next[42]), .E(n719), .CK(clk), .Q(
        \block[3][42] ) );
  EDFFXL \block_reg[7][42]  ( .D(block_next[42]), .E(n646), .CK(clk), .Q(
        \block[7][42] ) );
  EDFFXL \block_reg[6][54]  ( .D(block_next[54]), .E(n666), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFXL \block_reg[0][54]  ( .D(block_next[54]), .E(n773), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFXL \block_reg[4][54]  ( .D(block_next[54]), .E(n702), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFXL \block_reg[1][54]  ( .D(block_next[54]), .E(n754), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFXL \block_reg[5][54]  ( .D(block_next[54]), .E(n685), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFXL \block_reg[3][54]  ( .D(block_next[54]), .E(n720), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFXL \block_reg[7][54]  ( .D(block_next[54]), .E(n647), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFXL \block_reg[6][43]  ( .D(block_next[43]), .E(n665), .CK(clk), .Q(
        \block[6][43] ) );
  EDFFXL \block_reg[0][43]  ( .D(block_next[43]), .E(n772), .CK(clk), .Q(
        \block[0][43] ) );
  EDFFXL \block_reg[4][43]  ( .D(block_next[43]), .E(n701), .CK(clk), .Q(
        \block[4][43] ) );
  EDFFXL \block_reg[1][43]  ( .D(block_next[43]), .E(n753), .CK(clk), .Q(
        \block[1][43] ) );
  EDFFXL \block_reg[5][43]  ( .D(block_next[43]), .E(n684), .CK(clk), .Q(
        \block[5][43] ) );
  EDFFXL \block_reg[3][43]  ( .D(block_next[43]), .E(n719), .CK(clk), .Q(
        \block[3][43] ) );
  EDFFXL \block_reg[7][43]  ( .D(block_next[43]), .E(n646), .CK(clk), .Q(
        \block[7][43] ) );
  EDFFXL \block_reg[6][55]  ( .D(block_next[55]), .E(n666), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFXL \block_reg[0][55]  ( .D(block_next[55]), .E(n773), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFXL \block_reg[4][55]  ( .D(block_next[55]), .E(n702), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFXL \block_reg[1][55]  ( .D(block_next[55]), .E(n754), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFXL \block_reg[5][55]  ( .D(block_next[55]), .E(n685), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFXL \block_reg[3][55]  ( .D(block_next[55]), .E(n720), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFXL \block_reg[7][55]  ( .D(block_next[55]), .E(n647), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFXL \block_reg[6][1]  ( .D(block_next[1]), .E(n662), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFXL \block_reg[0][1]  ( .D(block_next[1]), .E(n769), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFXL \block_reg[4][1]  ( .D(block_next[1]), .E(n698), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFXL \block_reg[1][1]  ( .D(block_next[1]), .E(n750), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFXL \block_reg[5][1]  ( .D(block_next[1]), .E(n681), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFXL \block_reg[3][1]  ( .D(block_next[1]), .E(n716), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFXL \block_reg[7][1]  ( .D(block_next[1]), .E(n643), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFXL \block_reg[6][44]  ( .D(block_next[44]), .E(n665), .CK(clk), .Q(
        \block[6][44] ) );
  EDFFXL \block_reg[0][44]  ( .D(block_next[44]), .E(n772), .CK(clk), .Q(
        \block[0][44] ) );
  EDFFXL \block_reg[4][44]  ( .D(block_next[44]), .E(n701), .CK(clk), .Q(
        \block[4][44] ) );
  EDFFXL \block_reg[1][44]  ( .D(block_next[44]), .E(n753), .CK(clk), .Q(
        \block[1][44] ) );
  EDFFXL \block_reg[5][44]  ( .D(block_next[44]), .E(n684), .CK(clk), .Q(
        \block[5][44] ) );
  EDFFXL \block_reg[3][44]  ( .D(block_next[44]), .E(n719), .CK(clk), .Q(
        \block[3][44] ) );
  EDFFXL \block_reg[7][44]  ( .D(block_next[44]), .E(n646), .CK(clk), .Q(
        \block[7][44] ) );
  EDFFXL \block_reg[6][56]  ( .D(block_next[56]), .E(n666), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFXL \block_reg[0][56]  ( .D(block_next[56]), .E(n773), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFXL \block_reg[4][56]  ( .D(block_next[56]), .E(n702), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFXL \block_reg[1][56]  ( .D(block_next[56]), .E(n754), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFXL \block_reg[5][56]  ( .D(block_next[56]), .E(n685), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFXL \block_reg[3][56]  ( .D(block_next[56]), .E(n720), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFXL \block_reg[7][56]  ( .D(block_next[56]), .E(n647), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFXL \block_reg[6][21]  ( .D(block_next[21]), .E(n663), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFXL \block_reg[6][2]  ( .D(block_next[2]), .E(n662), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFXL \block_reg[0][2]  ( .D(block_next[2]), .E(n769), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFXL \block_reg[4][2]  ( .D(block_next[2]), .E(n698), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFXL \block_reg[1][2]  ( .D(block_next[2]), .E(n750), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFXL \block_reg[5][2]  ( .D(block_next[2]), .E(n681), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFXL \block_reg[3][2]  ( .D(block_next[2]), .E(n716), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFXL \block_reg[7][2]  ( .D(block_next[2]), .E(n643), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFXL \block_reg[6][45]  ( .D(block_next[45]), .E(n665), .CK(clk), .Q(
        \block[6][45] ) );
  EDFFXL \block_reg[0][45]  ( .D(block_next[45]), .E(n772), .CK(clk), .Q(
        \block[0][45] ) );
  EDFFXL \block_reg[4][45]  ( .D(block_next[45]), .E(n701), .CK(clk), .Q(
        \block[4][45] ) );
  EDFFXL \block_reg[1][45]  ( .D(block_next[45]), .E(n753), .CK(clk), .Q(
        \block[1][45] ) );
  EDFFXL \block_reg[5][45]  ( .D(block_next[45]), .E(n684), .CK(clk), .Q(
        \block[5][45] ) );
  EDFFXL \block_reg[3][45]  ( .D(block_next[45]), .E(n719), .CK(clk), .Q(
        \block[3][45] ) );
  EDFFXL \block_reg[7][45]  ( .D(block_next[45]), .E(n646), .CK(clk), .Q(
        \block[7][45] ) );
  EDFFXL \block_reg[6][57]  ( .D(block_next[57]), .E(n666), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFXL \block_reg[0][57]  ( .D(block_next[57]), .E(n773), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFXL \block_reg[4][57]  ( .D(block_next[57]), .E(n702), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFXL \block_reg[1][57]  ( .D(block_next[57]), .E(n754), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFXL \block_reg[5][57]  ( .D(block_next[57]), .E(n685), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFXL \block_reg[3][57]  ( .D(block_next[57]), .E(n720), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFXL \block_reg[7][57]  ( .D(block_next[57]), .E(n647), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFXL \block_reg[6][3]  ( .D(block_next[3]), .E(n662), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFXL \block_reg[0][3]  ( .D(block_next[3]), .E(n769), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFXL \block_reg[4][3]  ( .D(block_next[3]), .E(n698), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFXL \block_reg[1][3]  ( .D(block_next[3]), .E(n750), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFXL \block_reg[5][3]  ( .D(block_next[3]), .E(n681), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFXL \block_reg[3][3]  ( .D(block_next[3]), .E(n716), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFXL \block_reg[7][3]  ( .D(block_next[3]), .E(n643), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFXL \block_reg[6][46]  ( .D(block_next[46]), .E(n665), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFXL \block_reg[0][46]  ( .D(block_next[46]), .E(n772), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFXL \block_reg[4][46]  ( .D(block_next[46]), .E(n701), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFXL \block_reg[1][46]  ( .D(block_next[46]), .E(n753), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFXL \block_reg[5][46]  ( .D(block_next[46]), .E(n684), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFXL \block_reg[3][46]  ( .D(block_next[46]), .E(n719), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFXL \block_reg[7][46]  ( .D(block_next[46]), .E(n646), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFXL \block_reg[6][58]  ( .D(block_next[58]), .E(n666), .CK(clk), .Q(
        \block[6][58] ) );
  EDFFXL \block_reg[0][58]  ( .D(block_next[58]), .E(n773), .CK(clk), .Q(
        \block[0][58] ) );
  EDFFXL \block_reg[4][58]  ( .D(block_next[58]), .E(n702), .CK(clk), .Q(
        \block[4][58] ) );
  EDFFXL \block_reg[1][58]  ( .D(block_next[58]), .E(n754), .CK(clk), .Q(
        \block[1][58] ) );
  EDFFXL \block_reg[5][58]  ( .D(block_next[58]), .E(n685), .CK(clk), .Q(
        \block[5][58] ) );
  EDFFXL \block_reg[3][58]  ( .D(block_next[58]), .E(n720), .CK(clk), .Q(
        \block[3][58] ) );
  EDFFXL \block_reg[7][58]  ( .D(block_next[58]), .E(n647), .CK(clk), .Q(
        \block[7][58] ) );
  EDFFXL \block_reg[6][4]  ( .D(block_next[4]), .E(n662), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFXL \block_reg[0][4]  ( .D(block_next[4]), .E(n769), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFXL \block_reg[4][4]  ( .D(block_next[4]), .E(n698), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFXL \block_reg[1][4]  ( .D(block_next[4]), .E(n750), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFXL \block_reg[5][4]  ( .D(block_next[4]), .E(n681), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFXL \block_reg[3][4]  ( .D(block_next[4]), .E(n716), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFXL \block_reg[7][4]  ( .D(block_next[4]), .E(n643), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFXL \block_reg[6][47]  ( .D(block_next[47]), .E(n665), .CK(clk), .Q(
        \block[6][47] ) );
  EDFFXL \block_reg[0][47]  ( .D(block_next[47]), .E(n772), .CK(clk), .Q(
        \block[0][47] ) );
  EDFFXL \block_reg[4][47]  ( .D(block_next[47]), .E(n701), .CK(clk), .Q(
        \block[4][47] ) );
  EDFFXL \block_reg[1][47]  ( .D(block_next[47]), .E(n753), .CK(clk), .Q(
        \block[1][47] ) );
  EDFFXL \block_reg[5][47]  ( .D(block_next[47]), .E(n684), .CK(clk), .Q(
        \block[5][47] ) );
  EDFFXL \block_reg[3][47]  ( .D(block_next[47]), .E(n719), .CK(clk), .Q(
        \block[3][47] ) );
  EDFFXL \block_reg[7][47]  ( .D(block_next[47]), .E(n646), .CK(clk), .Q(
        \block[7][47] ) );
  EDFFXL \block_reg[6][59]  ( .D(block_next[59]), .E(n666), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFXL \block_reg[0][59]  ( .D(block_next[59]), .E(n773), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFXL \block_reg[4][59]  ( .D(block_next[59]), .E(n702), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFXL \block_reg[1][59]  ( .D(block_next[59]), .E(n754), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFXL \block_reg[5][59]  ( .D(block_next[59]), .E(n685), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFXL \block_reg[3][59]  ( .D(block_next[59]), .E(n720), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFXL \block_reg[7][59]  ( .D(block_next[59]), .E(n647), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFXL \block_reg[6][5]  ( .D(block_next[5]), .E(n662), .CK(clk), .Q(
        \block[6][5] ) );
  EDFFXL \block_reg[0][5]  ( .D(block_next[5]), .E(n769), .CK(clk), .QN(n130)
         );
  EDFFXL \block_reg[4][5]  ( .D(block_next[5]), .E(n698), .CK(clk), .Q(
        \block[4][5] ) );
  EDFFXL \block_reg[1][5]  ( .D(block_next[5]), .E(n750), .CK(clk), .QN(n131)
         );
  EDFFXL \block_reg[5][5]  ( .D(block_next[5]), .E(n681), .CK(clk), .Q(
        \block[5][5] ) );
  EDFFXL \block_reg[3][5]  ( .D(block_next[5]), .E(n716), .CK(clk), .QN(n133)
         );
  EDFFXL \block_reg[7][5]  ( .D(block_next[5]), .E(n643), .CK(clk), .Q(
        \block[7][5] ) );
  EDFFXL \block_reg[6][48]  ( .D(block_next[48]), .E(n665), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFXL \block_reg[0][48]  ( .D(block_next[48]), .E(n772), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFXL \block_reg[4][48]  ( .D(block_next[48]), .E(n701), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFXL \block_reg[1][48]  ( .D(block_next[48]), .E(n753), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFXL \block_reg[5][48]  ( .D(block_next[48]), .E(n684), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFXL \block_reg[3][48]  ( .D(block_next[48]), .E(n719), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFXL \block_reg[7][48]  ( .D(block_next[48]), .E(n646), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFXL \block_reg[6][60]  ( .D(block_next[60]), .E(n666), .CK(clk), .Q(
        \block[6][60] ) );
  EDFFXL \block_reg[0][60]  ( .D(block_next[60]), .E(n773), .CK(clk), .Q(
        \block[0][60] ) );
  EDFFXL \block_reg[4][60]  ( .D(block_next[60]), .E(n702), .CK(clk), .Q(
        \block[4][60] ) );
  EDFFXL \block_reg[1][60]  ( .D(block_next[60]), .E(n754), .CK(clk), .Q(
        \block[1][60] ) );
  EDFFXL \block_reg[5][60]  ( .D(block_next[60]), .E(n685), .CK(clk), .Q(
        \block[5][60] ) );
  EDFFXL \block_reg[3][60]  ( .D(block_next[60]), .E(n720), .CK(clk), .Q(
        \block[3][60] ) );
  EDFFXL \block_reg[7][60]  ( .D(block_next[60]), .E(n647), .CK(clk), .Q(
        \block[7][60] ) );
  EDFFXL \block_reg[6][6]  ( .D(block_next[6]), .E(n662), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFXL \block_reg[0][6]  ( .D(block_next[6]), .E(n769), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFXL \block_reg[4][6]  ( .D(block_next[6]), .E(n698), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFXL \block_reg[1][6]  ( .D(block_next[6]), .E(n750), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFXL \block_reg[5][6]  ( .D(block_next[6]), .E(n681), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFXL \block_reg[3][6]  ( .D(block_next[6]), .E(n716), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFXL \block_reg[7][6]  ( .D(block_next[6]), .E(n643), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFXL \block_reg[6][50]  ( .D(block_next[50]), .E(n665), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFXL \block_reg[0][50]  ( .D(block_next[50]), .E(n772), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFXL \block_reg[4][50]  ( .D(block_next[50]), .E(n701), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFXL \block_reg[1][50]  ( .D(block_next[50]), .E(n753), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFXL \block_reg[5][50]  ( .D(block_next[50]), .E(n684), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFXL \block_reg[3][50]  ( .D(block_next[50]), .E(n719), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFXL \block_reg[7][50]  ( .D(block_next[50]), .E(n646), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFXL \block_reg[6][61]  ( .D(block_next[61]), .E(n666), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFXL \block_reg[0][61]  ( .D(block_next[61]), .E(n773), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFXL \block_reg[4][61]  ( .D(block_next[61]), .E(n702), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFXL \block_reg[1][61]  ( .D(block_next[61]), .E(n754), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFXL \block_reg[5][61]  ( .D(block_next[61]), .E(n685), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFXL \block_reg[3][61]  ( .D(block_next[61]), .E(n720), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFXL \block_reg[7][61]  ( .D(block_next[61]), .E(n647), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFXL \block_reg[6][7]  ( .D(block_next[7]), .E(n662), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFXL \block_reg[6][51]  ( .D(block_next[51]), .E(n665), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFXL \block_reg[0][51]  ( .D(block_next[51]), .E(n772), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFXL \block_reg[4][51]  ( .D(block_next[51]), .E(n701), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFXL \block_reg[1][51]  ( .D(block_next[51]), .E(n753), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFXL \block_reg[5][51]  ( .D(block_next[51]), .E(n684), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFXL \block_reg[3][51]  ( .D(block_next[51]), .E(n719), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFXL \block_reg[7][51]  ( .D(block_next[51]), .E(n646), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFXL \block_reg[6][62]  ( .D(block_next[62]), .E(n666), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFXL \block_reg[0][62]  ( .D(block_next[62]), .E(n773), .CK(clk), .Q(
        \block[0][62] ) );
  EDFFXL \block_reg[4][62]  ( .D(block_next[62]), .E(n702), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFXL \block_reg[1][62]  ( .D(block_next[62]), .E(n754), .CK(clk), .Q(
        \block[1][62] ) );
  EDFFXL \block_reg[5][62]  ( .D(block_next[62]), .E(n685), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFXL \block_reg[3][62]  ( .D(block_next[62]), .E(n720), .CK(clk), .Q(
        \block[3][62] ) );
  EDFFXL \block_reg[7][62]  ( .D(block_next[62]), .E(n647), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFXL \block_reg[6][49]  ( .D(block_next[49]), .E(n665), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFXL \block_reg[6][63]  ( .D(block_next[63]), .E(n666), .CK(clk), .Q(
        \block[6][63] ) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n493), .CK(clk), .RN(n792), .Q(blockdirty[6]), .QN(n477) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n492), .CK(clk), .RN(n791), .Q(blockdirty[5]), .QN(n476) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n491), .CK(clk), .RN(n791), .Q(blockdirty[4]), .QN(n475) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n490), .CK(clk), .RN(n791), .Q(blockdirty[3]), .QN(n474) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n489), .CK(clk), .RN(n791), .Q(blockdirty[2]), .QN(n473) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n488), .CK(clk), .RN(n791), .Q(blockdirty[1]), .QN(n472) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n487), .CK(clk), .RN(n791), .Q(blockdirty[0]), .QN(n471) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n494), .CK(clk), .RN(n792), .Q(blockdirty[7]), .QN(n478) );
  EDFFXL \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n660), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFXL \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n731), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFXL \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n696), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFXL \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n767), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFXL \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n679), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFXL \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n748), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFXL \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n641), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFXL \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n714), .CK(clk), .Q(
        \blocktag[3][9] ) );
  XOR2X2 U3 ( .A(n1032), .B(proc_addr[21]), .Y(n803) );
  XNOR2X2 U4 ( .A(proc_addr[10]), .B(tag[5]), .Y(n795) );
  XOR2X1 U5 ( .A(n1041), .B(proc_addr[18]), .Y(n813) );
  XOR2X1 U6 ( .A(tag[9]), .B(proc_addr[14]), .Y(n800) );
  XOR2X1 U7 ( .A(tag[4]), .B(proc_addr[9]), .Y(n799) );
  XOR2X1 U8 ( .A(n1047), .B(proc_addr[16]), .Y(n802) );
  BUFX8 U9 ( .A(n868), .Y(n588) );
  NOR2X4 U10 ( .A(n808), .B(n807), .Y(n826) );
  AND2X6 U11 ( .A(n151), .B(n594), .Y(n147) );
  INVX1 U12 ( .A(mem_ready), .Y(n1086) );
  AND2X4 U13 ( .A(n1081), .B(n792), .Y(n138) );
  BUFX8 U14 ( .A(n1), .Y(n604) );
  CLKINVX2 U15 ( .A(n1095), .Y(n56) );
  CLKAND2X4 U16 ( .A(n147), .B(n608), .Y(n144) );
  CLKINVX4 U17 ( .A(tag[15]), .Y(n1035) );
  CLKINVX4 U18 ( .A(tag[7]), .Y(n1057) );
  CLKINVX4 U19 ( .A(tag[8]), .Y(n1054) );
  CLKINVX6 U20 ( .A(tag[21]), .Y(n1017) );
  INVX3 U21 ( .A(blockdata[3]), .Y(n1117) );
  INVX3 U22 ( .A(blockdata[4]), .Y(n1122) );
  INVX3 U23 ( .A(blockdata[5]), .Y(n1127) );
  INVX3 U24 ( .A(blockdata[6]), .Y(n1132) );
  INVX4 U25 ( .A(n1289), .Y(n21) );
  CLKAND2X3 U26 ( .A(mem_write), .B(blockdata[0]), .Y(n1289) );
  INVX4 U27 ( .A(n1288), .Y(n23) );
  CLKAND2X3 U28 ( .A(mem_write), .B(blockdata[121]), .Y(n1288) );
  INVX4 U29 ( .A(n1287), .Y(n25) );
  CLKAND2X3 U30 ( .A(mem_write), .B(blockdata[122]), .Y(n1287) );
  INVX4 U31 ( .A(n1286), .Y(n27) );
  CLKAND2X3 U32 ( .A(mem_write), .B(blockdata[123]), .Y(n1286) );
  INVX4 U33 ( .A(n1285), .Y(n29) );
  CLKAND2X3 U34 ( .A(mem_write), .B(blockdata[124]), .Y(n1285) );
  INVX4 U35 ( .A(n1284), .Y(n31) );
  CLKAND2X3 U36 ( .A(mem_write), .B(blockdata[125]), .Y(n1284) );
  INVX4 U37 ( .A(n1283), .Y(n33) );
  CLKAND2X3 U38 ( .A(mem_write), .B(blockdata[126]), .Y(n1283) );
  INVX4 U39 ( .A(n1282), .Y(n35) );
  CLKAND2X3 U40 ( .A(mem_write), .B(blockdata[127]), .Y(n1282) );
  OAI221X1 U41 ( .A0(n637), .A1(n1162), .B0(n633), .B1(n1161), .C0(n1160), .Y(
        proc_rdata[12]) );
  OAI221X1 U42 ( .A0(n637), .A1(n1167), .B0(n633), .B1(n1166), .C0(n1165), .Y(
        proc_rdata[13]) );
  OAI221X1 U43 ( .A0(n637), .A1(n1217), .B0(n633), .B1(n1216), .C0(n1215), .Y(
        proc_rdata[23]) );
  INVX4 U44 ( .A(n1060), .Y(blocktag_next[4]) );
  NAND2X2 U45 ( .A(mem_rdata[119]), .B(n616), .Y(n844) );
  NAND2X2 U46 ( .A(mem_rdata[77]), .B(n616), .Y(n889) );
  NAND2X2 U47 ( .A(mem_rdata[92]), .B(n616), .Y(n874) );
  NAND2X2 U48 ( .A(mem_rdata[97]), .B(n616), .Y(n866) );
  NAND2X2 U49 ( .A(mem_rdata[98]), .B(n616), .Y(n865) );
  CLKINVX4 U50 ( .A(N32), .Y(n784) );
  BUFX2 U51 ( .A(n583), .Y(n551) );
  BUFX4 U52 ( .A(n515), .Y(n523) );
  INVX4 U53 ( .A(N31), .Y(n783) );
  BUFX8 U54 ( .A(N31), .Y(n583) );
  BUFX2 U55 ( .A(n551), .Y(n556) );
  INVX3 U56 ( .A(n834), .Y(n1070) );
  AND2X4 U57 ( .A(n1077), .B(n792), .Y(n136) );
  BUFX2 U58 ( .A(n582), .Y(n550) );
  CLKBUFX3 U59 ( .A(n138), .Y(n710) );
  BUFX2 U60 ( .A(n547), .Y(n520) );
  BUFX2 U61 ( .A(n547), .Y(n521) );
  BUFX4 U62 ( .A(n1070), .Y(n620) );
  BUFX2 U63 ( .A(n547), .Y(n515) );
  INVX6 U64 ( .A(n870), .Y(n903) );
  NAND3X4 U65 ( .A(n57), .B(n832), .C(n1096), .Y(n1) );
  CLKMX2X12 U66 ( .A(tag[5]), .B(proc_addr[10]), .S0(n609), .Y(n2) );
  BUFX2 U67 ( .A(n551), .Y(n557) );
  INVX3 U68 ( .A(n1090), .Y(n1263) );
  BUFX8 U69 ( .A(n150), .Y(n585) );
  BUFX12 U70 ( .A(n150), .Y(n584) );
  AND3X4 U71 ( .A(n56), .B(n832), .C(n1096), .Y(n55) );
  INVX8 U72 ( .A(n1003), .Y(n832) );
  AND4X2 U73 ( .A(n869), .B(n594), .C(n600), .D(n606), .Y(n150) );
  CLKINVX12 U74 ( .A(n601), .Y(n600) );
  OAI221X1 U75 ( .A0(n636), .A1(n1102), .B0(n632), .B1(n1101), .C0(n1100), .Y(
        proc_rdata[0]) );
  OAI221X1 U76 ( .A0(n636), .A1(n1112), .B0(n632), .B1(n1111), .C0(n1110), .Y(
        proc_rdata[2]) );
  OAI221X1 U77 ( .A0(n636), .A1(n1117), .B0(n632), .B1(n1116), .C0(n1115), .Y(
        proc_rdata[3]) );
  OAI221X1 U78 ( .A0(n636), .A1(n1152), .B0(n632), .B1(n1151), .C0(n1150), .Y(
        proc_rdata[10]) );
  OAI221X1 U79 ( .A0(n635), .A1(n1237), .B0(n634), .B1(n1236), .C0(n1235), .Y(
        proc_rdata[27]) );
  OAI221XL U80 ( .A0(n635), .A1(n1260), .B0(n634), .B1(n1258), .C0(n1257), .Y(
        proc_rdata[31]) );
  OAI221XL U81 ( .A0(n635), .A1(n1242), .B0(n634), .B1(n1241), .C0(n1240), .Y(
        proc_rdata[28]) );
  OAI221X1 U82 ( .A0(n635), .A1(n1252), .B0(n634), .B1(n1251), .C0(n1250), .Y(
        proc_rdata[30]) );
  OAI221X1 U83 ( .A0(n635), .A1(n1222), .B0(n634), .B1(n1221), .C0(n1220), .Y(
        proc_rdata[24]) );
  BUFX2 U84 ( .A(n631), .Y(n634) );
  BUFX20 U85 ( .A(n630), .Y(n632) );
  OAI221X1 U86 ( .A0(n636), .A1(n1107), .B0(n632), .B1(n1106), .C0(n1105), .Y(
        proc_rdata[1]) );
  OAI221X1 U87 ( .A0(n636), .A1(n1147), .B0(n632), .B1(n1146), .C0(n1145), .Y(
        proc_rdata[9]) );
  OAI221X1 U88 ( .A0(n636), .A1(n1122), .B0(n632), .B1(n1121), .C0(n1120), .Y(
        proc_rdata[4]) );
  OAI221X1 U89 ( .A0(n636), .A1(n1157), .B0(n632), .B1(n1156), .C0(n1155), .Y(
        proc_rdata[11]) );
  OAI221X1 U90 ( .A0(n636), .A1(n1137), .B0(n632), .B1(n1136), .C0(n1135), .Y(
        proc_rdata[7]) );
  OAI221X1 U91 ( .A0(n636), .A1(n1142), .B0(n632), .B1(n1141), .C0(n1140), .Y(
        proc_rdata[8]) );
  OAI221X1 U92 ( .A0(n636), .A1(n1132), .B0(n632), .B1(n1131), .C0(n1130), .Y(
        proc_rdata[6]) );
  OAI221X1 U93 ( .A0(n636), .A1(n1127), .B0(n632), .B1(n1126), .C0(n1125), .Y(
        proc_rdata[5]) );
  BUFX20 U94 ( .A(n630), .Y(n633) );
  OAI221X1 U95 ( .A0(n637), .A1(n1202), .B0(n633), .B1(n1201), .C0(n1200), .Y(
        proc_rdata[20]) );
  OAI221X1 U96 ( .A0(n637), .A1(n1212), .B0(n633), .B1(n1211), .C0(n1210), .Y(
        proc_rdata[22]) );
  OAI221X1 U97 ( .A0(n637), .A1(n1182), .B0(n633), .B1(n1181), .C0(n1180), .Y(
        proc_rdata[16]) );
  OAI221X1 U98 ( .A0(n637), .A1(n1177), .B0(n633), .B1(n1176), .C0(n1175), .Y(
        proc_rdata[15]) );
  OAI221X1 U99 ( .A0(n637), .A1(n1172), .B0(n633), .B1(n1171), .C0(n1170), .Y(
        proc_rdata[14]) );
  OAI221X1 U100 ( .A0(n637), .A1(n1192), .B0(n633), .B1(n1191), .C0(n1190), 
        .Y(proc_rdata[18]) );
  OAI221X1 U101 ( .A0(n637), .A1(n1197), .B0(n633), .B1(n1196), .C0(n1195), 
        .Y(proc_rdata[19]) );
  OAI221X1 U102 ( .A0(n637), .A1(n1207), .B0(n633), .B1(n1206), .C0(n1205), 
        .Y(proc_rdata[21]) );
  INVX4 U103 ( .A(n1052), .Y(blocktag_next[9]) );
  CLKBUFX4 U104 ( .A(n627), .Y(n629) );
  OA22X2 U105 ( .A0(n629), .A1(n1184), .B0(n625), .B1(n1183), .Y(n1185) );
  OA22X2 U106 ( .A0(n629), .A1(n1199), .B0(n625), .B1(n1198), .Y(n1200) );
  OA22X2 U107 ( .A0(n629), .A1(n1179), .B0(n625), .B1(n1178), .Y(n1180) );
  OA22X2 U108 ( .A0(n629), .A1(n1209), .B0(n625), .B1(n1208), .Y(n1210) );
  OA22X2 U109 ( .A0(n629), .A1(n1174), .B0(n625), .B1(n1173), .Y(n1175) );
  OA22X2 U110 ( .A0(n629), .A1(n1194), .B0(n625), .B1(n1193), .Y(n1195) );
  OA22X2 U111 ( .A0(n629), .A1(n1189), .B0(n625), .B1(n1188), .Y(n1190) );
  OA22X2 U112 ( .A0(n629), .A1(n1169), .B0(n625), .B1(n1168), .Y(n1170) );
  OA22X2 U113 ( .A0(n629), .A1(n1204), .B0(n625), .B1(n1203), .Y(n1205) );
  OAI211X4 U114 ( .A0(mem_ready), .A1(valid), .B0(n829), .C0(n1087), .Y(n830)
         );
  CLKINVX8 U115 ( .A(n830), .Y(n869) );
  BUFX2 U116 ( .A(n627), .Y(n628) );
  OA22X1 U117 ( .A0(n628), .A1(n1124), .B0(n624), .B1(n1123), .Y(n1125) );
  OA22X1 U118 ( .A0(n628), .A1(n1104), .B0(n624), .B1(n1103), .Y(n1105) );
  OA22X1 U119 ( .A0(n628), .A1(n1144), .B0(n624), .B1(n1143), .Y(n1145) );
  OA22X1 U120 ( .A0(n628), .A1(n1119), .B0(n624), .B1(n1118), .Y(n1120) );
  OA22X1 U121 ( .A0(n628), .A1(n1149), .B0(n624), .B1(n1148), .Y(n1150) );
  OA22X1 U122 ( .A0(n628), .A1(n1154), .B0(n624), .B1(n1153), .Y(n1155) );
  OA22X1 U123 ( .A0(n628), .A1(n1129), .B0(n624), .B1(n1128), .Y(n1130) );
  OA22X1 U124 ( .A0(n628), .A1(n1134), .B0(n624), .B1(n1133), .Y(n1135) );
  OA22X1 U125 ( .A0(n628), .A1(n1139), .B0(n624), .B1(n1138), .Y(n1140) );
  BUFX20 U126 ( .A(n604), .Y(n606) );
  OAI221X4 U127 ( .A0(n585), .A1(n1171), .B0(n972), .B1(n587), .C0(n853), .Y(
        block_next[110]) );
  OAI221X4 U128 ( .A0(n584), .A1(n1201), .B0(n960), .B1(n586), .C0(n847), .Y(
        block_next[116]) );
  OAI221X4 U129 ( .A0(n585), .A1(n1166), .B0(n974), .B1(n587), .C0(n854), .Y(
        block_next[109]) );
  OAI221X4 U130 ( .A0(n585), .A1(n1161), .B0(n976), .B1(n587), .C0(n855), .Y(
        block_next[108]) );
  OAI221X4 U131 ( .A0(n637), .A1(n1187), .B0(n633), .B1(n1186), .C0(n1185), 
        .Y(proc_rdata[17]) );
  XOR2X4 U132 ( .A(n1029), .B(proc_addr[22]), .Y(n812) );
  OA22X2 U133 ( .A0(n626), .A1(n1229), .B0(n623), .B1(n1228), .Y(n1230) );
  OA22X2 U134 ( .A0(n626), .A1(n1234), .B0(n623), .B1(n1233), .Y(n1235) );
  OA22X2 U135 ( .A0(n626), .A1(n1239), .B0(n623), .B1(n1238), .Y(n1240) );
  OA22X2 U136 ( .A0(n626), .A1(n1244), .B0(n623), .B1(n1243), .Y(n1245) );
  OA22X2 U137 ( .A0(n626), .A1(n1249), .B0(n623), .B1(n1248), .Y(n1250) );
  OA22X2 U138 ( .A0(n626), .A1(n1255), .B0(n623), .B1(n1253), .Y(n1257) );
  OA22X2 U139 ( .A0(n626), .A1(n1224), .B0(n623), .B1(n1223), .Y(n1225) );
  MXI4X2 U140 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n577), .S1(n541), .Y(n454) );
  MXI4X2 U141 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n577), .S1(n541), .Y(n452) );
  MXI4X2 U142 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n577), .S1(n541), .Y(n453) );
  MXI4X2 U143 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n577), .S1(n541), .Y(n451) );
  MX4X1 U144 ( .A(n130), .B(n131), .C(n132), .D(n133), .S0(n577), .S1(n541), 
        .Y(n449) );
  BUFX20 U145 ( .A(n554), .Y(n577) );
  NAND2X4 U146 ( .A(mem_rdata[7]), .B(n611), .Y(n985) );
  NAND2X4 U147 ( .A(mem_rdata[12]), .B(n611), .Y(n975) );
  NAND2X4 U148 ( .A(mem_rdata[13]), .B(n611), .Y(n973) );
  NAND2X4 U149 ( .A(mem_rdata[8]), .B(n611), .Y(n983) );
  NAND2X4 U150 ( .A(mem_rdata[9]), .B(n611), .Y(n981) );
  NAND2X4 U151 ( .A(mem_rdata[10]), .B(n611), .Y(n979) );
  NAND2X4 U152 ( .A(mem_rdata[11]), .B(n611), .Y(n977) );
  NAND2X4 U153 ( .A(mem_rdata[1]), .B(n611), .Y(n997) );
  BUFX20 U154 ( .A(n621), .Y(n611) );
  NAND2X4 U155 ( .A(mem_rdata[21]), .B(n612), .Y(n957) );
  NAND2X4 U156 ( .A(mem_rdata[20]), .B(n612), .Y(n959) );
  NAND2X4 U157 ( .A(mem_rdata[19]), .B(n612), .Y(n961) );
  NAND2X4 U158 ( .A(mem_rdata[14]), .B(n612), .Y(n971) );
  NAND2X4 U159 ( .A(mem_rdata[15]), .B(n612), .Y(n969) );
  NAND2X4 U160 ( .A(mem_rdata[16]), .B(n612), .Y(n967) );
  NAND2X4 U161 ( .A(mem_rdata[17]), .B(n612), .Y(n965) );
  NAND2X4 U162 ( .A(mem_rdata[18]), .B(n612), .Y(n963) );
  BUFX20 U163 ( .A(n621), .Y(n612) );
  NAND2X4 U164 ( .A(mem_rdata[96]), .B(n611), .Y(n867) );
  NAND2X4 U165 ( .A(mem_rdata[99]), .B(n612), .Y(n864) );
  NAND2X4 U166 ( .A(mem_rdata[104]), .B(n611), .Y(n859) );
  NAND2X4 U167 ( .A(mem_rdata[93]), .B(n621), .Y(n873) );
  NAND2X4 U168 ( .A(mem_rdata[94]), .B(n612), .Y(n872) );
  OAI221X4 U169 ( .A0(n607), .A1(n964), .B0(n603), .B1(n1192), .C0(n963), .Y(
        block_next[18]) );
  OAI221X4 U170 ( .A0(n607), .A1(n966), .B0(n603), .B1(n1187), .C0(n965), .Y(
        block_next[17]) );
  OAI221X4 U171 ( .A0(n607), .A1(n968), .B0(n603), .B1(n1182), .C0(n967), .Y(
        block_next[16]) );
  OAI221X4 U172 ( .A0(n606), .A1(n978), .B0(n603), .B1(n1157), .C0(n977), .Y(
        block_next[11]) );
  OAI221X4 U173 ( .A0(n606), .A1(n980), .B0(n603), .B1(n1152), .C0(n979), .Y(
        block_next[10]) );
  OAI221X4 U174 ( .A0(n607), .A1(n970), .B0(n603), .B1(n1177), .C0(n969), .Y(
        block_next[15]) );
  OAI221X4 U175 ( .A0(n607), .A1(n972), .B0(n603), .B1(n1172), .C0(n971), .Y(
        block_next[14]) );
  OAI221X4 U176 ( .A0(n607), .A1(n962), .B0(n603), .B1(n1197), .C0(n961), .Y(
        block_next[19]) );
  OAI221X4 U177 ( .A0(n607), .A1(n974), .B0(n603), .B1(n1167), .C0(n973), .Y(
        block_next[13]) );
  OAI221X4 U178 ( .A0(n606), .A1(n976), .B0(n603), .B1(n1162), .C0(n975), .Y(
        block_next[12]) );
  OAI221X4 U179 ( .A0(n589), .A1(n1255), .B0(n938), .B1(n594), .C0(n871), .Y(
        block_next[95]) );
  NOR2BX2 U180 ( .AN(proc_read), .B(n833), .Y(n203) );
  NAND4X4 U181 ( .A(n819), .B(n818), .C(n817), .D(n816), .Y(n823) );
  XOR2X4 U182 ( .A(n1072), .B(proc_addr[5]), .Y(n819) );
  CLKINVX6 U183 ( .A(tag[0]), .Y(n1072) );
  BUFX8 U184 ( .A(n620), .Y(n619) );
  BUFX20 U185 ( .A(n620), .Y(n616) );
  CLKMX2X4 U186 ( .A(n177), .B(n178), .S0(n512), .Y(tag[20]) );
  BUFX20 U187 ( .A(n467), .Y(n512) );
  INVX8 U188 ( .A(n1273), .Y(n3) );
  INVX20 U189 ( .A(n3), .Y(mem_addr[18]) );
  INVX8 U190 ( .A(n1277), .Y(n5) );
  INVX20 U191 ( .A(n5), .Y(mem_addr[14]) );
  INVX8 U192 ( .A(n1276), .Y(n7) );
  INVX20 U193 ( .A(n7), .Y(mem_addr[15]) );
  INVX8 U194 ( .A(n1275), .Y(n9) );
  INVX20 U195 ( .A(n9), .Y(mem_addr[16]) );
  INVX8 U196 ( .A(n1274), .Y(n11) );
  INVX20 U197 ( .A(n11), .Y(mem_addr[17]) );
  INVX8 U198 ( .A(n1272), .Y(n13) );
  INVX20 U199 ( .A(n13), .Y(mem_addr[19]) );
  INVX8 U200 ( .A(n1268), .Y(n15) );
  INVX20 U201 ( .A(n15), .Y(mem_addr[23]) );
  INVX8 U202 ( .A(n1266), .Y(n17) );
  INVX20 U203 ( .A(n17), .Y(mem_addr[25]) );
  INVX8 U204 ( .A(n1265), .Y(n19) );
  INVX20 U205 ( .A(n19), .Y(mem_addr[26]) );
  CLKINVX20 U206 ( .A(n21), .Y(mem_wdata[0]) );
  CLKINVX20 U207 ( .A(n23), .Y(mem_wdata[121]) );
  CLKINVX20 U208 ( .A(n25), .Y(mem_wdata[122]) );
  CLKINVX20 U209 ( .A(n27), .Y(mem_wdata[123]) );
  CLKINVX20 U210 ( .A(n29), .Y(mem_wdata[124]) );
  CLKINVX20 U211 ( .A(n31), .Y(mem_wdata[125]) );
  CLKINVX20 U212 ( .A(n33), .Y(mem_wdata[126]) );
  CLKINVX20 U213 ( .A(n35), .Y(mem_wdata[127]) );
  XOR2X4 U214 ( .A(tag[14]), .B(n1037), .Y(n804) );
  CLKINVX4 U215 ( .A(tag[14]), .Y(n1038) );
  CLKMX2X3 U216 ( .A(n191), .B(n192), .S0(n512), .Y(tag[14]) );
  BUFX20 U217 ( .A(n518), .Y(n542) );
  XOR2X4 U218 ( .A(n1014), .B(proc_addr[27]), .Y(n811) );
  INVX4 U219 ( .A(tag[22]), .Y(n1014) );
  BUFX20 U220 ( .A(n553), .Y(n578) );
  BUFX20 U221 ( .A(N31), .Y(n553) );
  NAND3BX4 U222 ( .AN(n833), .B(proc_write), .C(n831), .Y(n1003) );
  NAND2X6 U223 ( .A(valid), .B(n828), .Y(n833) );
  OAI221X4 U224 ( .A0(n585), .A1(n1156), .B0(n978), .B1(n587), .C0(n856), .Y(
        block_next[107]) );
  NAND3BX4 U225 ( .AN(n1097), .B(proc_addr[0]), .C(n1096), .Y(n1254) );
  NAND2X4 U226 ( .A(n203), .B(n1093), .Y(n1097) );
  OA22X2 U227 ( .A0(n626), .A1(n1219), .B0(n623), .B1(n1218), .Y(n1220) );
  XNOR2X4 U228 ( .A(n1035), .B(proc_addr[20]), .Y(n148) );
  CLKMX2X3 U229 ( .A(n189), .B(n190), .S0(n512), .Y(tag[21]) );
  CLKMX2X3 U230 ( .A(n185), .B(n186), .S0(n512), .Y(tag[23]) );
  CLKMX2X3 U231 ( .A(n193), .B(n194), .S0(n512), .Y(tag[19]) );
  CLKMX2X3 U232 ( .A(n171), .B(n172), .S0(n512), .Y(tag[12]) );
  CLKMX2X3 U233 ( .A(n173), .B(n174), .S0(n512), .Y(tag[22]) );
  CLKMX2X3 U234 ( .A(n181), .B(n182), .S0(n512), .Y(tag[16]) );
  CLKMX2X2 U235 ( .A(n157), .B(n158), .S0(n512), .Y(tag[18]) );
  CLKMX2X3 U236 ( .A(n197), .B(n198), .S0(n512), .Y(tag[17]) );
  INVX6 U237 ( .A(n1002), .Y(proc_stall) );
  NAND2X4 U238 ( .A(n1087), .B(n833), .Y(n1002) );
  XOR2X4 U239 ( .A(n1020), .B(proc_addr[25]), .Y(n821) );
  CLKINVX6 U240 ( .A(tag[20]), .Y(n1020) );
  BUFX20 U241 ( .A(n517), .Y(n543) );
  BUFX12 U242 ( .A(N32), .Y(n517) );
  XOR2X1 U243 ( .A(n1023), .B(proc_addr[24]), .Y(n820) );
  OAI221X4 U244 ( .A0(n585), .A1(n1151), .B0(n980), .B1(n587), .C0(n857), .Y(
        block_next[106]) );
  XOR2X4 U245 ( .A(n1008), .B(proc_addr[29]), .Y(n817) );
  INVX4 U246 ( .A(tag[24]), .Y(n1008) );
  BUFX20 U247 ( .A(n619), .Y(n617) );
  BUFX20 U248 ( .A(n517), .Y(n545) );
  OAI221X4 U249 ( .A0(n584), .A1(n1136), .B0(n986), .B1(n588), .C0(n860), .Y(
        block_next[103]) );
  OAI221X4 U250 ( .A0(n585), .A1(n1146), .B0(n982), .B1(n587), .C0(n858), .Y(
        block_next[105]) );
  OAI221X4 U251 ( .A0(n585), .A1(n1141), .B0(n984), .B1(n587), .C0(n859), .Y(
        block_next[104]) );
  OAI221X4 U252 ( .A0(n585), .A1(n1191), .B0(n964), .B1(n587), .C0(n849), .Y(
        block_next[114]) );
  OAI221X4 U253 ( .A0(n585), .A1(n1181), .B0(n968), .B1(n587), .C0(n851), .Y(
        block_next[112]) );
  BUFX6 U254 ( .A(n55), .Y(n601) );
  BUFX20 U255 ( .A(n903), .Y(n590) );
  BUFX20 U256 ( .A(n903), .Y(n589) );
  OAI221X4 U257 ( .A0(n589), .A1(n1249), .B0(n940), .B1(n594), .C0(n872), .Y(
        block_next[94]) );
  OAI221X4 U258 ( .A0(n590), .A1(n1189), .B0(n964), .B1(n593), .C0(n884), .Y(
        block_next[82]) );
  AND2XL U259 ( .A(N31), .B(n1091), .Y(mem_addr[0]) );
  OAI221X4 U260 ( .A0(n589), .A1(n1244), .B0(n942), .B1(n594), .C0(n873), .Y(
        block_next[93]) );
  OAI221X4 U261 ( .A0(n590), .A1(n1184), .B0(n966), .B1(n593), .C0(n885), .Y(
        block_next[81]) );
  OAI221X4 U262 ( .A0(n589), .A1(n1239), .B0(n944), .B1(n594), .C0(n874), .Y(
        block_next[92]) );
  OAI221X4 U263 ( .A0(n590), .A1(n1179), .B0(n968), .B1(n593), .C0(n886), .Y(
        block_next[80]) );
  OAI221X4 U264 ( .A0(n589), .A1(n1234), .B0(n946), .B1(n594), .C0(n875), .Y(
        block_next[91]) );
  BUFX20 U265 ( .A(n622), .Y(n610) );
  CLKMX2X4 U266 ( .A(n1029), .B(n1028), .S0(n610), .Y(n1030) );
  CLKMX2X4 U267 ( .A(n1020), .B(n1019), .S0(n610), .Y(n1021) );
  CLKMX2X4 U268 ( .A(n1011), .B(n1010), .S0(n610), .Y(n1012) );
  CLKMX2X4 U269 ( .A(n1026), .B(n1025), .S0(n610), .Y(n1027) );
  CLKMX2X4 U270 ( .A(n1017), .B(n1016), .S0(n610), .Y(n1018) );
  CLKMX2X4 U271 ( .A(n1038), .B(n1037), .S0(n610), .Y(n1039) );
  CLKMX2X4 U272 ( .A(n1035), .B(n1034), .S0(n610), .Y(n1036) );
  CLKMX2X4 U273 ( .A(n1041), .B(n1040), .S0(n610), .Y(n1042) );
  OAI221X4 U274 ( .A0(n589), .A1(n1229), .B0(n948), .B1(n594), .C0(n876), .Y(
        block_next[90]) );
  OAI221X4 U275 ( .A0(n589), .A1(n1224), .B0(n950), .B1(n594), .C0(n877), .Y(
        block_next[89]) );
  OAI221X4 U276 ( .A0(n589), .A1(n1219), .B0(n952), .B1(n594), .C0(n878), .Y(
        block_next[88]) );
  OAI221X4 U277 ( .A0(n589), .A1(n1214), .B0(n954), .B1(n593), .C0(n879), .Y(
        block_next[87]) );
  OAI221X4 U278 ( .A0(n589), .A1(n1209), .B0(n956), .B1(n593), .C0(n880), .Y(
        block_next[86]) );
  OAI221X4 U279 ( .A0(n589), .A1(n1204), .B0(n958), .B1(n593), .C0(n881), .Y(
        block_next[85]) );
  OAI221X4 U280 ( .A0(n590), .A1(n1099), .B0(n1000), .B1(n592), .C0(n902), .Y(
        block_next[64]) );
  OAI221X4 U281 ( .A0(n590), .A1(n1174), .B0(n970), .B1(n593), .C0(n887), .Y(
        block_next[79]) );
  MXI2X1 U282 ( .A(tag[6]), .B(proc_addr[11]), .S0(n609), .Y(n1059) );
  CLKMX2X4 U283 ( .A(n1068), .B(n1067), .S0(n609), .Y(n1069) );
  CLKMX2X4 U284 ( .A(n1062), .B(n1061), .S0(n609), .Y(n1063) );
  CLKMX2X4 U285 ( .A(n1057), .B(n1056), .S0(n609), .Y(n1058) );
  CLKMX2X4 U286 ( .A(n1065), .B(n1064), .S0(n609), .Y(n1066) );
  CLKMX2X4 U287 ( .A(n1072), .B(n1071), .S0(n609), .Y(n1073) );
  CLKMX2X4 U288 ( .A(n1054), .B(n1053), .S0(n609), .Y(n1055) );
  CLKMX2X4 U289 ( .A(n1050), .B(n1049), .S0(n609), .Y(n1051) );
  BUFX20 U290 ( .A(n622), .Y(n609) );
  OAI221X4 U291 ( .A0(n589), .A1(n1199), .B0(n960), .B1(n593), .C0(n882), .Y(
        block_next[84]) );
  NAND4X4 U292 ( .A(n812), .B(n811), .C(n810), .D(n809), .Y(n815) );
  XOR2X4 U293 ( .A(n1054), .B(proc_addr[13]), .Y(n805) );
  XOR2X4 U294 ( .A(n1057), .B(proc_addr[12]), .Y(n806) );
  NAND2X2 U295 ( .A(n821), .B(n820), .Y(n822) );
  OA21X2 U296 ( .A0(n1002), .A1(n1086), .B0(dirty), .Y(n1004) );
  BUFX12 U297 ( .A(n517), .Y(n546) );
  NAND2X4 U298 ( .A(dirty), .B(valid), .Y(n1089) );
  AO21X2 U299 ( .A0(mem_ready), .A1(n1087), .B0(valid), .Y(n1001) );
  MXI2X4 U300 ( .A(n461), .B(n462), .S0(n511), .Y(valid) );
  XNOR2X2 U301 ( .A(proc_addr[23]), .B(tag[18]), .Y(n797) );
  NOR4X4 U302 ( .A(n801), .B(n800), .C(n799), .D(n798), .Y(n827) );
  XOR2X1 U303 ( .A(tag[6]), .B(proc_addr[11]), .Y(n798) );
  AND2XL U304 ( .A(N32), .B(n1091), .Y(mem_addr[1]) );
  AND2XL U305 ( .A(N33), .B(n1091), .Y(mem_addr[2]) );
  OAI221X4 U306 ( .A0(n584), .A1(n1221), .B0(n952), .B1(n586), .C0(n843), .Y(
        block_next[120]) );
  OAI221X4 U307 ( .A0(n584), .A1(n1216), .B0(n954), .B1(n586), .C0(n844), .Y(
        block_next[119]) );
  OAI221X4 U308 ( .A0(n584), .A1(n1211), .B0(n956), .B1(n586), .C0(n845), .Y(
        block_next[118]) );
  OAI221X4 U309 ( .A0(n584), .A1(n1231), .B0(n948), .B1(n586), .C0(n841), .Y(
        block_next[122]) );
  OAI221X4 U310 ( .A0(n584), .A1(n1226), .B0(n950), .B1(n586), .C0(n842), .Y(
        block_next[121]) );
  OAI221X4 U311 ( .A0(n584), .A1(n1258), .B0(n938), .B1(n586), .C0(n835), .Y(
        block_next[127]) );
  OAI221X4 U312 ( .A0(n584), .A1(n1251), .B0(n940), .B1(n586), .C0(n837), .Y(
        block_next[126]) );
  OAI221X4 U313 ( .A0(n584), .A1(n1246), .B0(n942), .B1(n586), .C0(n838), .Y(
        block_next[125]) );
  MXI2X1 U314 ( .A(tag[4]), .B(proc_addr[9]), .S0(n609), .Y(n1060) );
  OAI221X4 U315 ( .A0(n585), .A1(n1196), .B0(n962), .B1(n587), .C0(n848), .Y(
        block_next[115]) );
  OAI221X4 U316 ( .A0(n590), .A1(n1159), .B0(n976), .B1(n592), .C0(n890), .Y(
        block_next[76]) );
  NAND2X2 U317 ( .A(mem_rdata[76]), .B(n616), .Y(n890) );
  OAI221X4 U318 ( .A0(n590), .A1(n1154), .B0(n978), .B1(n592), .C0(n891), .Y(
        block_next[75]) );
  OAI221X4 U319 ( .A0(n590), .A1(n1149), .B0(n980), .B1(n592), .C0(n892), .Y(
        block_next[74]) );
  OAI221X4 U320 ( .A0(n590), .A1(n1144), .B0(n982), .B1(n592), .C0(n893), .Y(
        block_next[73]) );
  OAI221X4 U321 ( .A0(n590), .A1(n1139), .B0(n984), .B1(n592), .C0(n894), .Y(
        block_next[72]) );
  OAI221X4 U322 ( .A0(n590), .A1(n1129), .B0(n988), .B1(n592), .C0(n896), .Y(
        block_next[70]) );
  OAI221X4 U323 ( .A0(n589), .A1(n1124), .B0(n990), .B1(n592), .C0(n897), .Y(
        block_next[69]) );
  OAI221X4 U324 ( .A0(n590), .A1(n1169), .B0(n972), .B1(n593), .C0(n888), .Y(
        block_next[78]) );
  OAI221X4 U325 ( .A0(n590), .A1(n1119), .B0(n992), .B1(n592), .C0(n898), .Y(
        block_next[68]) );
  OAI221X4 U326 ( .A0(n590), .A1(n1164), .B0(n974), .B1(n593), .C0(n889), .Y(
        block_next[77]) );
  OAI221X4 U327 ( .A0(n589), .A1(n1114), .B0(n994), .B1(n592), .C0(n899), .Y(
        block_next[67]) );
  OAI221X4 U328 ( .A0(n903), .A1(n1134), .B0(n986), .B1(n593), .C0(n895), .Y(
        block_next[71]) );
  OAI221X4 U329 ( .A0(n903), .A1(n1109), .B0(n996), .B1(n592), .C0(n900), .Y(
        block_next[66]) );
  BUFX16 U330 ( .A(n622), .Y(n613) );
  AND2X8 U331 ( .A(n869), .B(n588), .Y(n151) );
  NAND2BXL U332 ( .AN(n1004), .B(n1003), .Y(n1005) );
  OAI221X4 U333 ( .A0(n585), .A1(n1106), .B0(n998), .B1(n588), .C0(n866), .Y(
        block_next[97]) );
  OAI221X4 U334 ( .A0(n585), .A1(n1111), .B0(n996), .B1(n588), .C0(n865), .Y(
        block_next[98]) );
  OAI221X4 U335 ( .A0(n584), .A1(n1116), .B0(n994), .B1(n588), .C0(n864), .Y(
        block_next[99]) );
  OAI221X4 U336 ( .A0(n585), .A1(n1121), .B0(n992), .B1(n588), .C0(n863), .Y(
        block_next[100]) );
  OAI221X4 U337 ( .A0(n584), .A1(n1126), .B0(n990), .B1(n588), .C0(n862), .Y(
        block_next[101]) );
  OAI221X4 U338 ( .A0(n585), .A1(n1131), .B0(n988), .B1(n588), .C0(n861), .Y(
        block_next[102]) );
  AND2XL U339 ( .A(n789), .B(blockdata[7]), .Y(mem_wdata[7]) );
  AND2XL U340 ( .A(n788), .B(blockdata[37]), .Y(mem_wdata[37]) );
  AND2XL U341 ( .A(n789), .B(blockdata[8]), .Y(mem_wdata[8]) );
  AND2XL U342 ( .A(n788), .B(blockdata[46]), .Y(mem_wdata[46]) );
  AND2XL U343 ( .A(n789), .B(blockdata[9]), .Y(mem_wdata[9]) );
  AND2XL U344 ( .A(n788), .B(blockdata[47]), .Y(mem_wdata[47]) );
  AND2XL U345 ( .A(n789), .B(blockdata[10]), .Y(mem_wdata[10]) );
  AND2XL U346 ( .A(n788), .B(blockdata[48]), .Y(mem_wdata[48]) );
  OAI221X4 U347 ( .A0(n595), .A1(n1253), .B0(n938), .B1(n600), .C0(n905), .Y(
        block_next[63]) );
  OAI221X4 U348 ( .A0(n596), .A1(n1183), .B0(n966), .B1(n599), .C0(n919), .Y(
        block_next[49]) );
  AND2XL U349 ( .A(n789), .B(blockdata[11]), .Y(mem_wdata[11]) );
  AND2XL U350 ( .A(n788), .B(blockdata[49]), .Y(mem_wdata[49]) );
  AND2XL U351 ( .A(n789), .B(blockdata[12]), .Y(mem_wdata[12]) );
  AND2XL U352 ( .A(n788), .B(blockdata[50]), .Y(mem_wdata[50]) );
  AND2XL U353 ( .A(n789), .B(blockdata[13]), .Y(mem_wdata[13]) );
  AND2XL U354 ( .A(n788), .B(blockdata[51]), .Y(mem_wdata[51]) );
  OAI221X4 U355 ( .A0(n595), .A1(n1248), .B0(n940), .B1(n600), .C0(n906), .Y(
        block_next[62]) );
  OAI221X4 U356 ( .A0(n596), .A1(n1193), .B0(n962), .B1(n599), .C0(n917), .Y(
        block_next[51]) );
  AND2XL U357 ( .A(n789), .B(blockdata[14]), .Y(mem_wdata[14]) );
  AND2XL U358 ( .A(n788), .B(blockdata[52]), .Y(mem_wdata[52]) );
  OAI221X4 U359 ( .A0(n606), .A1(n986), .B0(n603), .B1(n1137), .C0(n985), .Y(
        block_next[7]) );
  AND2XL U360 ( .A(n789), .B(blockdata[15]), .Y(mem_wdata[15]) );
  AND2XL U361 ( .A(n788), .B(blockdata[53]), .Y(mem_wdata[53]) );
  OAI221X4 U362 ( .A0(n595), .A1(n1243), .B0(n942), .B1(n600), .C0(n907), .Y(
        block_next[61]) );
  OAI221X4 U363 ( .A0(n596), .A1(n1188), .B0(n964), .B1(n599), .C0(n918), .Y(
        block_next[50]) );
  AND2XL U364 ( .A(n789), .B(blockdata[16]), .Y(mem_wdata[16]) );
  AND2XL U365 ( .A(n788), .B(blockdata[54]), .Y(mem_wdata[54]) );
  OAI221X4 U366 ( .A0(n606), .A1(n988), .B0(n603), .B1(n1132), .C0(n987), .Y(
        block_next[6]) );
  AND2XL U367 ( .A(n789), .B(blockdata[17]), .Y(mem_wdata[17]) );
  AND2XL U368 ( .A(n788), .B(blockdata[55]), .Y(mem_wdata[55]) );
  OAI221X4 U369 ( .A0(n595), .A1(n1238), .B0(n944), .B1(n600), .C0(n908), .Y(
        block_next[60]) );
  OAI221X4 U370 ( .A0(n596), .A1(n1178), .B0(n968), .B1(n599), .C0(n920), .Y(
        block_next[48]) );
  AND2XL U371 ( .A(n789), .B(blockdata[18]), .Y(mem_wdata[18]) );
  AND2XL U372 ( .A(n788), .B(blockdata[56]), .Y(mem_wdata[56]) );
  OAI221X4 U373 ( .A0(n606), .A1(n990), .B0(n603), .B1(n1127), .C0(n989), .Y(
        block_next[5]) );
  AND2XL U374 ( .A(n789), .B(blockdata[19]), .Y(mem_wdata[19]) );
  AND2XL U375 ( .A(n788), .B(blockdata[57]), .Y(mem_wdata[57]) );
  OAI221X4 U376 ( .A0(n595), .A1(n1233), .B0(n946), .B1(n600), .C0(n909), .Y(
        block_next[59]) );
  AND2XL U377 ( .A(n789), .B(blockdata[20]), .Y(mem_wdata[20]) );
  AND2XL U378 ( .A(n788), .B(blockdata[58]), .Y(mem_wdata[58]) );
  OAI221X4 U379 ( .A0(n596), .A1(n1173), .B0(n970), .B1(n599), .C0(n921), .Y(
        block_next[47]) );
  OAI221X4 U380 ( .A0(n606), .A1(n992), .B0(n603), .B1(n1122), .C0(n991), .Y(
        block_next[4]) );
  AND2XL U381 ( .A(n789), .B(blockdata[21]), .Y(mem_wdata[21]) );
  AND2XL U382 ( .A(n788), .B(blockdata[59]), .Y(mem_wdata[59]) );
  OAI221X4 U383 ( .A0(n595), .A1(n1228), .B0(n948), .B1(n600), .C0(n910), .Y(
        block_next[58]) );
  AND2XL U384 ( .A(n789), .B(blockdata[22]), .Y(mem_wdata[22]) );
  AND2XL U385 ( .A(n788), .B(blockdata[60]), .Y(mem_wdata[60]) );
  OAI221X4 U386 ( .A0(n596), .A1(n1168), .B0(n972), .B1(n599), .C0(n922), .Y(
        block_next[46]) );
  OAI221X4 U387 ( .A0(n606), .A1(n994), .B0(n603), .B1(n1117), .C0(n993), .Y(
        block_next[3]) );
  AND2XL U388 ( .A(n789), .B(blockdata[23]), .Y(mem_wdata[23]) );
  AND2XL U389 ( .A(n788), .B(blockdata[61]), .Y(mem_wdata[61]) );
  AND2XL U390 ( .A(n789), .B(blockdata[24]), .Y(mem_wdata[24]) );
  AND2XL U391 ( .A(n788), .B(blockdata[62]), .Y(mem_wdata[62]) );
  OAI221X4 U392 ( .A0(n595), .A1(n1223), .B0(n950), .B1(n600), .C0(n911), .Y(
        block_next[57]) );
  OAI221X4 U393 ( .A0(n596), .A1(n1163), .B0(n974), .B1(n599), .C0(n923), .Y(
        block_next[45]) );
  OAI221X4 U394 ( .A0(n606), .A1(n996), .B0(n603), .B1(n1112), .C0(n995), .Y(
        block_next[2]) );
  AND2XL U395 ( .A(n789), .B(blockdata[25]), .Y(mem_wdata[25]) );
  AND2XL U396 ( .A(n788), .B(blockdata[63]), .Y(mem_wdata[63]) );
  AND2XL U397 ( .A(mem_write), .B(blockdata[83]), .Y(mem_wdata[83]) );
  OAI221X4 U398 ( .A0(n607), .A1(n958), .B0(n602), .B1(n1207), .C0(n957), .Y(
        block_next[21]) );
  AND2XL U399 ( .A(n789), .B(blockdata[26]), .Y(mem_wdata[26]) );
  AND2XL U400 ( .A(n788), .B(blockdata[64]), .Y(mem_wdata[64]) );
  AND2XL U401 ( .A(mem_write), .B(blockdata[84]), .Y(mem_wdata[84]) );
  OAI221X4 U402 ( .A0(n595), .A1(n1218), .B0(n952), .B1(n600), .C0(n912), .Y(
        block_next[56]) );
  OAI221X4 U403 ( .A0(n596), .A1(n1158), .B0(n976), .B1(n598), .C0(n924), .Y(
        block_next[44]) );
  OAI221X4 U404 ( .A0(n606), .A1(n998), .B0(n603), .B1(n1107), .C0(n997), .Y(
        block_next[1]) );
  AND2XL U405 ( .A(n789), .B(blockdata[27]), .Y(mem_wdata[27]) );
  AND2XL U406 ( .A(n788), .B(blockdata[65]), .Y(mem_wdata[65]) );
  AND2XL U407 ( .A(mem_write), .B(blockdata[85]), .Y(mem_wdata[85]) );
  AND2XL U408 ( .A(n789), .B(blockdata[28]), .Y(mem_wdata[28]) );
  AND2XL U409 ( .A(n788), .B(blockdata[66]), .Y(mem_wdata[66]) );
  AND2XL U410 ( .A(mem_write), .B(blockdata[86]), .Y(mem_wdata[86]) );
  OAI221X4 U411 ( .A0(n595), .A1(n1213), .B0(n954), .B1(n599), .C0(n913), .Y(
        block_next[55]) );
  AND2XL U412 ( .A(n789), .B(blockdata[29]), .Y(mem_wdata[29]) );
  AND2XL U413 ( .A(n788), .B(blockdata[67]), .Y(mem_wdata[67]) );
  OAI221X4 U414 ( .A0(n596), .A1(n1153), .B0(n978), .B1(n598), .C0(n925), .Y(
        block_next[43]) );
  AND2XL U415 ( .A(mem_write), .B(blockdata[87]), .Y(mem_wdata[87]) );
  AND2XL U416 ( .A(n789), .B(blockdata[30]), .Y(mem_wdata[30]) );
  AND2XL U417 ( .A(n788), .B(blockdata[68]), .Y(mem_wdata[68]) );
  AND2XL U418 ( .A(mem_write), .B(blockdata[88]), .Y(mem_wdata[88]) );
  AND2XL U419 ( .A(n789), .B(blockdata[31]), .Y(mem_wdata[31]) );
  AND2XL U420 ( .A(n788), .B(blockdata[69]), .Y(mem_wdata[69]) );
  OAI221X4 U421 ( .A0(n595), .A1(n1208), .B0(n956), .B1(n599), .C0(n914), .Y(
        block_next[54]) );
  OAI221X4 U422 ( .A0(n596), .A1(n1148), .B0(n980), .B1(n598), .C0(n926), .Y(
        block_next[42]) );
  AND2XL U423 ( .A(mem_write), .B(blockdata[89]), .Y(mem_wdata[89]) );
  AND2XL U424 ( .A(n789), .B(blockdata[32]), .Y(mem_wdata[32]) );
  AND2XL U425 ( .A(n788), .B(blockdata[70]), .Y(mem_wdata[70]) );
  AND2XL U426 ( .A(mem_write), .B(blockdata[90]), .Y(mem_wdata[90]) );
  AND2XL U427 ( .A(n789), .B(blockdata[33]), .Y(mem_wdata[33]) );
  AND2XL U428 ( .A(n788), .B(blockdata[71]), .Y(mem_wdata[71]) );
  AND2XL U429 ( .A(mem_write), .B(blockdata[91]), .Y(mem_wdata[91]) );
  AND2XL U430 ( .A(n789), .B(blockdata[34]), .Y(mem_wdata[34]) );
  AND2XL U431 ( .A(n788), .B(blockdata[72]), .Y(mem_wdata[72]) );
  AND2XL U432 ( .A(mem_write), .B(blockdata[92]), .Y(mem_wdata[92]) );
  OAI221X4 U433 ( .A0(n597), .A1(n1128), .B0(n988), .B1(n598), .C0(n930), .Y(
        block_next[38]) );
  CLKBUFX4 U434 ( .A(n144), .Y(n597) );
  OAI221X4 U435 ( .A0(n597), .A1(n1123), .B0(n990), .B1(n598), .C0(n931), .Y(
        block_next[37]) );
  OAI221X4 U436 ( .A0(n597), .A1(n1118), .B0(n992), .B1(n598), .C0(n932), .Y(
        block_next[36]) );
  OAI221X4 U437 ( .A0(n597), .A1(n1113), .B0(n994), .B1(n598), .C0(n933), .Y(
        block_next[35]) );
  OAI221X4 U438 ( .A0(n597), .A1(n1108), .B0(n996), .B1(n598), .C0(n934), .Y(
        block_next[34]) );
  OAI221X4 U439 ( .A0(n597), .A1(n1103), .B0(n998), .B1(n598), .C0(n935), .Y(
        block_next[33]) );
  OAI221X4 U440 ( .A0(n597), .A1(n1133), .B0(n986), .B1(n599), .C0(n929), .Y(
        block_next[39]) );
  AND2XL U441 ( .A(n789), .B(blockdata[35]), .Y(mem_wdata[35]) );
  AND2XL U442 ( .A(n788), .B(blockdata[73]), .Y(mem_wdata[73]) );
  AND2XL U443 ( .A(mem_write), .B(blockdata[93]), .Y(mem_wdata[93]) );
  OAI221X4 U444 ( .A0(n608), .A1(n944), .B0(n602), .B1(n1242), .C0(n943), .Y(
        block_next[28]) );
  OAI221X4 U445 ( .A0(n608), .A1(n946), .B0(n602), .B1(n1237), .C0(n945), .Y(
        block_next[27]) );
  AND2XL U446 ( .A(n789), .B(blockdata[36]), .Y(mem_wdata[36]) );
  AND2XL U447 ( .A(n788), .B(blockdata[74]), .Y(mem_wdata[74]) );
  AND2XL U448 ( .A(mem_write), .B(blockdata[94]), .Y(mem_wdata[94]) );
  OAI221X4 U449 ( .A0(n608), .A1(n938), .B0(n602), .B1(n1260), .C0(n937), .Y(
        block_next[31]) );
  OAI221X4 U450 ( .A0(n608), .A1(n940), .B0(n602), .B1(n1252), .C0(n939), .Y(
        block_next[30]) );
  OAI221X4 U451 ( .A0(n608), .A1(n942), .B0(n602), .B1(n1247), .C0(n941), .Y(
        block_next[29]) );
  OAI221X4 U452 ( .A0(n608), .A1(n948), .B0(n602), .B1(n1232), .C0(n947), .Y(
        block_next[26]) );
  AND2XL U453 ( .A(n789), .B(blockdata[38]), .Y(mem_wdata[38]) );
  AND2XL U454 ( .A(n788), .B(blockdata[75]), .Y(mem_wdata[75]) );
  AND2XL U455 ( .A(mem_write), .B(blockdata[95]), .Y(mem_wdata[95]) );
  AND2XL U456 ( .A(n789), .B(blockdata[39]), .Y(mem_wdata[39]) );
  AND2XL U457 ( .A(n788), .B(blockdata[76]), .Y(mem_wdata[76]) );
  AND2XL U458 ( .A(mem_write), .B(blockdata[96]), .Y(mem_wdata[96]) );
  OAI221X4 U459 ( .A0(n608), .A1(n950), .B0(n602), .B1(n1227), .C0(n949), .Y(
        block_next[25]) );
  AND2XL U460 ( .A(n789), .B(blockdata[40]), .Y(mem_wdata[40]) );
  AND2XL U461 ( .A(n788), .B(blockdata[77]), .Y(mem_wdata[77]) );
  AND2XL U462 ( .A(mem_write), .B(blockdata[97]), .Y(mem_wdata[97]) );
  AND2XL U463 ( .A(n789), .B(blockdata[41]), .Y(mem_wdata[41]) );
  AND2XL U464 ( .A(n788), .B(blockdata[78]), .Y(mem_wdata[78]) );
  AND2XL U465 ( .A(mem_write), .B(blockdata[98]), .Y(mem_wdata[98]) );
  OAI221X4 U466 ( .A0(n607), .A1(n952), .B0(n602), .B1(n1222), .C0(n951), .Y(
        block_next[24]) );
  AND2XL U467 ( .A(n789), .B(blockdata[42]), .Y(mem_wdata[42]) );
  AND2XL U468 ( .A(n788), .B(blockdata[79]), .Y(mem_wdata[79]) );
  AND2XL U469 ( .A(mem_write), .B(blockdata[99]), .Y(mem_wdata[99]) );
  AND2XL U470 ( .A(n789), .B(blockdata[43]), .Y(mem_wdata[43]) );
  AND2XL U471 ( .A(n788), .B(blockdata[80]), .Y(mem_wdata[80]) );
  OAI221X4 U472 ( .A0(n607), .A1(n954), .B0(n602), .B1(n1217), .C0(n953), .Y(
        block_next[23]) );
  AND2XL U473 ( .A(mem_write), .B(blockdata[100]), .Y(mem_wdata[100]) );
  AND2XL U474 ( .A(n789), .B(blockdata[44]), .Y(mem_wdata[44]) );
  AND2XL U475 ( .A(n788), .B(blockdata[81]), .Y(mem_wdata[81]) );
  AND2XL U476 ( .A(mem_write), .B(blockdata[101]), .Y(mem_wdata[101]) );
  AND2XL U477 ( .A(n789), .B(blockdata[45]), .Y(mem_wdata[45]) );
  AND2XL U478 ( .A(n788), .B(blockdata[82]), .Y(mem_wdata[82]) );
  OAI221X4 U479 ( .A0(n607), .A1(n956), .B0(n602), .B1(n1212), .C0(n955), .Y(
        block_next[22]) );
  AND2XL U480 ( .A(mem_write), .B(blockdata[102]), .Y(mem_wdata[102]) );
  AND2XL U481 ( .A(mem_write), .B(blockdata[103]), .Y(mem_wdata[103]) );
  AND2XL U482 ( .A(mem_write), .B(blockdata[104]), .Y(mem_wdata[104]) );
  AND2XL U483 ( .A(mem_write), .B(blockdata[105]), .Y(mem_wdata[105]) );
  AND2XL U484 ( .A(mem_write), .B(blockdata[106]), .Y(mem_wdata[106]) );
  AND2XL U485 ( .A(mem_write), .B(blockdata[107]), .Y(mem_wdata[107]) );
  AND2XL U486 ( .A(mem_write), .B(blockdata[108]), .Y(mem_wdata[108]) );
  AND2XL U487 ( .A(mem_write), .B(blockdata[109]), .Y(mem_wdata[109]) );
  AND2XL U488 ( .A(mem_write), .B(blockdata[110]), .Y(mem_wdata[110]) );
  AND2XL U489 ( .A(mem_write), .B(blockdata[111]), .Y(mem_wdata[111]) );
  AND2XL U490 ( .A(mem_write), .B(blockdata[112]), .Y(mem_wdata[112]) );
  AND2XL U491 ( .A(mem_write), .B(blockdata[113]), .Y(mem_wdata[113]) );
  AND2XL U492 ( .A(mem_write), .B(blockdata[114]), .Y(mem_wdata[114]) );
  AND2XL U493 ( .A(mem_write), .B(blockdata[115]), .Y(mem_wdata[115]) );
  AND2XL U494 ( .A(mem_write), .B(blockdata[116]), .Y(mem_wdata[116]) );
  AND2XL U495 ( .A(mem_write), .B(blockdata[117]), .Y(mem_wdata[117]) );
  AND2XL U496 ( .A(mem_write), .B(blockdata[118]), .Y(mem_wdata[118]) );
  AND2XL U497 ( .A(mem_write), .B(blockdata[119]), .Y(mem_wdata[119]) );
  AND2XL U498 ( .A(mem_write), .B(blockdata[120]), .Y(mem_wdata[120]) );
  OAI221X4 U499 ( .A0(n597), .A1(n1098), .B0(n1000), .B1(n598), .C0(n936), .Y(
        block_next[32]) );
  OAI221X4 U500 ( .A0(n595), .A1(n1203), .B0(n958), .B1(n599), .C0(n915), .Y(
        block_next[53]) );
  CLKBUFX6 U501 ( .A(n144), .Y(n595) );
  OAI221X4 U502 ( .A0(n584), .A1(n1101), .B0(n1000), .B1(n588), .C0(n867), .Y(
        block_next[96]) );
  OAI221X4 U503 ( .A0(n607), .A1(n1000), .B0(n603), .B1(n1102), .C0(n999), .Y(
        block_next[0]) );
  OAI221X4 U504 ( .A0(n596), .A1(n1143), .B0(n982), .B1(n598), .C0(n927), .Y(
        block_next[41]) );
  CLKBUFX6 U505 ( .A(n144), .Y(n596) );
  OAI221X4 U506 ( .A0(n595), .A1(n1198), .B0(n960), .B1(n599), .C0(n916), .Y(
        block_next[52]) );
  OAI221X4 U507 ( .A0(n596), .A1(n1138), .B0(n984), .B1(n598), .C0(n928), .Y(
        block_next[40]) );
  XNOR2X1 U508 ( .A(proc_addr[7]), .B(tag[2]), .Y(n794) );
  MX2X6 U509 ( .A(n165), .B(n166), .S0(n513), .Y(tag[2]) );
  OAI221X4 U510 ( .A0(n606), .A1(n982), .B0(n603), .B1(n1147), .C0(n981), .Y(
        block_next[9]) );
  BUFX20 U511 ( .A(n145), .Y(n603) );
  XOR2X4 U512 ( .A(n1011), .B(proc_addr[28]), .Y(n818) );
  CLKINVX6 U513 ( .A(tag[23]), .Y(n1011) );
  OAI221X4 U514 ( .A0(n607), .A1(n960), .B0(n602), .B1(n1202), .C0(n959), .Y(
        block_next[20]) );
  CLKBUFX8 U515 ( .A(n145), .Y(n602) );
  BUFX20 U516 ( .A(n552), .Y(n580) );
  MX4X1 U517 ( .A(\blocktag[4][7] ), .B(\blocktag[5][7] ), .C(\blocktag[6][7] ), .D(\blocktag[7][7] ), .S0(n580), .S1(n545), .Y(n200) );
  MX4X1 U518 ( .A(\blocktag[4][8] ), .B(\blocktag[5][8] ), .C(\blocktag[6][8] ), .D(\blocktag[7][8] ), .S0(n580), .S1(n545), .Y(n170) );
  MX4X1 U519 ( .A(\blocktag[0][8] ), .B(\blocktag[1][8] ), .C(\blocktag[2][8] ), .D(\blocktag[3][8] ), .S0(n580), .S1(n545), .Y(n169) );
  OAI221X4 U520 ( .A0(n606), .A1(n984), .B0(n603), .B1(n1142), .C0(n983), .Y(
        block_next[8]) );
  OAI221X4 U521 ( .A0(n584), .A1(n1241), .B0(n944), .B1(n586), .C0(n839), .Y(
        block_next[124]) );
  XNOR2X4 U522 ( .A(proc_addr[8]), .B(tag[3]), .Y(n796) );
  MX2X6 U523 ( .A(n159), .B(n160), .S0(n513), .Y(tag[3]) );
  BUFX20 U524 ( .A(n552), .Y(n581) );
  BUFX8 U525 ( .A(N31), .Y(n552) );
  OAI221X4 U526 ( .A0(n585), .A1(n1186), .B0(n966), .B1(n587), .C0(n850), .Y(
        block_next[113]) );
  XOR2X2 U527 ( .A(n1068), .B(proc_addr[6]), .Y(n809) );
  CLKINVX4 U528 ( .A(tag[1]), .Y(n1068) );
  OAI221X4 U529 ( .A0(n584), .A1(n1236), .B0(n946), .B1(n586), .C0(n840), .Y(
        block_next[123]) );
  BUFX20 U530 ( .A(n553), .Y(n579) );
  NAND4BX4 U531 ( .AN(n1089), .B(n1088), .C(n1087), .D(n1086), .Y(n1090) );
  NAND4X6 U532 ( .A(n827), .B(n826), .C(n825), .D(n824), .Y(n1088) );
  AO22X4 U533 ( .A0(proc_addr[20]), .A1(mem_read), .B0(tag[15]), .B1(mem_write), .Y(n1273) );
  XOR2X4 U534 ( .A(n1017), .B(proc_addr[26]), .Y(n816) );
  CLKINVX8 U535 ( .A(n1088), .Y(n828) );
  BUFX20 U536 ( .A(n517), .Y(n544) );
  XNOR2X4 U537 ( .A(n1044), .B(proc_addr[17]), .Y(n149) );
  CLKINVX6 U538 ( .A(tag[12]), .Y(n1044) );
  MXI2X1 U539 ( .A(n447), .B(n448), .S0(n511), .Y(blockdata[6]) );
  INVX4 U540 ( .A(blockdata[2]), .Y(n1112) );
  MXI2X2 U541 ( .A(n455), .B(n456), .S0(n511), .Y(blockdata[2]) );
  MXI2X1 U542 ( .A(n449), .B(n450), .S0(n511), .Y(blockdata[5]) );
  CLKAND2X12 U543 ( .A(mem_write), .B(blockdata[6]), .Y(mem_wdata[6]) );
  MXI2X1 U544 ( .A(n451), .B(n452), .S0(n511), .Y(blockdata[4]) );
  CLKAND2X12 U545 ( .A(mem_write), .B(blockdata[5]), .Y(mem_wdata[5]) );
  MXI2X1 U546 ( .A(n453), .B(n454), .S0(n511), .Y(blockdata[3]) );
  CLKAND2X12 U547 ( .A(mem_write), .B(blockdata[4]), .Y(mem_wdata[4]) );
  INVX4 U548 ( .A(blockdata[1]), .Y(n1107) );
  MXI2X2 U549 ( .A(n457), .B(n458), .S0(n511), .Y(blockdata[1]) );
  CLKINVX6 U550 ( .A(n1267), .Y(n37) );
  INVX20 U551 ( .A(n37), .Y(mem_addr[24]) );
  AO22X1 U552 ( .A0(proc_addr[26]), .A1(mem_read), .B0(tag[21]), .B1(mem_write), .Y(n1267) );
  CLKINVX6 U553 ( .A(n1269), .Y(n39) );
  INVX20 U554 ( .A(n39), .Y(mem_addr[22]) );
  AO22X1 U555 ( .A0(proc_addr[24]), .A1(mem_read), .B0(tag[19]), .B1(mem_write), .Y(n1269) );
  CLKINVX6 U556 ( .A(n1270), .Y(n41) );
  INVX20 U557 ( .A(n41), .Y(mem_addr[21]) );
  AO22X1 U558 ( .A0(proc_addr[23]), .A1(mem_read), .B0(tag[18]), .B1(mem_write), .Y(n1270) );
  CLKAND2X12 U559 ( .A(mem_write), .B(blockdata[3]), .Y(mem_wdata[3]) );
  CLKINVX6 U560 ( .A(n1264), .Y(n43) );
  INVX20 U561 ( .A(n43), .Y(mem_addr[27]) );
  AO22X1 U562 ( .A0(proc_addr[29]), .A1(mem_read), .B0(tag[24]), .B1(mem_write), .Y(n1264) );
  CLKINVX6 U563 ( .A(n1278), .Y(n45) );
  INVX20 U564 ( .A(n45), .Y(mem_addr[11]) );
  AO22X1 U565 ( .A0(proc_addr[13]), .A1(mem_read), .B0(tag[8]), .B1(mem_write), 
        .Y(n1278) );
  CLKINVX6 U566 ( .A(n1279), .Y(n47) );
  INVX20 U567 ( .A(n47), .Y(mem_addr[9]) );
  AO22X1 U568 ( .A0(proc_addr[11]), .A1(mem_read), .B0(tag[6]), .B1(mem_write), 
        .Y(n1279) );
  CLKINVX6 U569 ( .A(n1280), .Y(n49) );
  INVX20 U570 ( .A(n49), .Y(mem_addr[6]) );
  AO22X1 U571 ( .A0(proc_addr[8]), .A1(mem_read), .B0(tag[3]), .B1(mem_write), 
        .Y(n1280) );
  CLKINVX6 U572 ( .A(n1281), .Y(n51) );
  INVX20 U573 ( .A(n51), .Y(mem_addr[3]) );
  AO22X1 U574 ( .A0(proc_addr[5]), .A1(mem_read), .B0(tag[0]), .B1(mem_write), 
        .Y(n1281) );
  CLKAND2X12 U575 ( .A(mem_write), .B(blockdata[2]), .Y(mem_wdata[2]) );
  CLKAND2X12 U576 ( .A(mem_write), .B(blockdata[1]), .Y(mem_wdata[1]) );
  INVX1 U577 ( .A(proc_wdata[16]), .Y(n968) );
  CLKINVX6 U578 ( .A(n1271), .Y(n53) );
  INVX20 U579 ( .A(n53), .Y(mem_addr[20]) );
  AO22X1 U580 ( .A0(proc_addr[22]), .A1(mem_read), .B0(tag[17]), .B1(mem_write), .Y(n1271) );
  INVXL U581 ( .A(proc_write), .Y(n1093) );
  CLKBUFX4 U582 ( .A(n465), .Y(n470) );
  BUFX4 U583 ( .A(n136), .Y(n744) );
  BUFX4 U584 ( .A(n639), .Y(n654) );
  BUFX4 U585 ( .A(n658), .Y(n673) );
  BUFX4 U586 ( .A(n765), .Y(n780) );
  BUFX4 U587 ( .A(n746), .Y(n761) );
  BUFX4 U588 ( .A(n677), .Y(n692) );
  BUFX4 U589 ( .A(n712), .Y(n727) );
  CLKBUFX3 U590 ( .A(n138), .Y(n709) );
  CLKBUFX2 U591 ( .A(n639), .Y(n653) );
  CLKBUFX2 U592 ( .A(n658), .Y(n672) );
  CLKBUFX2 U593 ( .A(n765), .Y(n779) );
  CLKBUFX2 U594 ( .A(n746), .Y(n760) );
  CLKBUFX2 U595 ( .A(n677), .Y(n691) );
  CLKBUFX2 U596 ( .A(n712), .Y(n726) );
  BUFX12 U597 ( .A(n619), .Y(n618) );
  BUFX12 U598 ( .A(n620), .Y(n615) );
  BUFX12 U599 ( .A(n620), .Y(n614) );
  BUFX8 U600 ( .A(n620), .Y(n621) );
  BUFX4 U601 ( .A(n1070), .Y(n622) );
  MXI4XL U602 ( .A(n82), .B(n83), .C(n84), .D(n85), .S0(n580), .S1(n544), .Y(
        n171) );
  MXI4X1 U603 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n580), .S1(n544), .Y(
        n172) );
  NAND2X1 U604 ( .A(mem_rdata[0]), .B(n610), .Y(n999) );
  AND2X4 U605 ( .A(n147), .B(n600), .Y(n145) );
  NAND2X1 U606 ( .A(n832), .B(n152), .Y(n868) );
  MXI4XL U607 ( .A(n62), .B(n63), .C(n64), .D(n65), .S0(n581), .S1(n546), .Y(
        n160) );
  MXI4XL U608 ( .A(n118), .B(n119), .C(n120), .D(n121), .S0(n578), .S1(N32), 
        .Y(n184) );
  CLKAND2X8 U609 ( .A(n1006), .B(n792), .Y(n134) );
  CLKAND2X8 U610 ( .A(n1075), .B(n792), .Y(n135) );
  CLKAND2X8 U611 ( .A(n1083), .B(n792), .Y(n139) );
  CLKAND2X8 U612 ( .A(n1079), .B(n792), .Y(n137) );
  BUFX20 U613 ( .A(n591), .Y(n594) );
  BUFX4 U614 ( .A(n793), .Y(n792) );
  INVX3 U615 ( .A(tag[19]), .Y(n1023) );
  MX4XL U616 ( .A(\blocktag[4][21] ), .B(\blocktag[5][21] ), .C(
        \blocktag[6][21] ), .D(\blocktag[7][21] ), .S0(n578), .S1(n543), .Y(
        n190) );
  MXI4XL U617 ( .A(n98), .B(n99), .C(n100), .D(n101), .S0(n579), .S1(n543), 
        .Y(n193) );
  MXI4XL U618 ( .A(n102), .B(n103), .C(n104), .D(n105), .S0(n578), .S1(n543), 
        .Y(n194) );
  AND2X6 U619 ( .A(n143), .B(n792), .Y(n141) );
  AND2X8 U620 ( .A(n146), .B(n792), .Y(n140) );
  BUFX8 U621 ( .A(n904), .Y(n591) );
  NOR2X4 U622 ( .A(n823), .B(n822), .Y(n824) );
  INVX3 U623 ( .A(tag[11]), .Y(n1047) );
  NAND2BX2 U624 ( .AN(n148), .B(n813), .Y(n814) );
  INVX3 U625 ( .A(tag[10]), .Y(n1050) );
  INVXL U626 ( .A(proc_addr[0]), .Y(n57) );
  CLKMX2X4 U627 ( .A(n153), .B(n154), .S0(n513), .Y(tag[6]) );
  CLKMX2X4 U628 ( .A(n201), .B(n202), .S0(n513), .Y(tag[1]) );
  MX4XL U629 ( .A(\blocktag[4][1] ), .B(\blocktag[5][1] ), .C(\blocktag[6][1] ), .D(\blocktag[7][1] ), .S0(n581), .S1(n546), .Y(n202) );
  MX4XL U630 ( .A(\blocktag[4][17] ), .B(\blocktag[5][17] ), .C(
        \blocktag[6][17] ), .D(\blocktag[7][17] ), .S0(n579), .S1(n544), .Y(
        n198) );
  MXI4XL U631 ( .A(n58), .B(n59), .C(n60), .D(n61), .S0(n581), .S1(n546), .Y(
        n159) );
  CLKMX2X4 U632 ( .A(n169), .B(n170), .S0(n513), .Y(tag[8]) );
  CLKMX2X4 U633 ( .A(n187), .B(n188), .S0(n513), .Y(tag[0]) );
  MXI4XL U634 ( .A(n94), .B(n95), .C(n96), .D(n97), .S0(n578), .S1(n543), .Y(
        n186) );
  MXI4XL U635 ( .A(n90), .B(n91), .C(n92), .D(n93), .S0(n578), .S1(n543), .Y(
        n185) );
  CLKMX2X4 U636 ( .A(n199), .B(n200), .S0(n513), .Y(tag[7]) );
  MXI4XL U637 ( .A(n78), .B(n79), .C(n80), .D(n81), .S0(n578), .S1(n543), .Y(
        n174) );
  MXI4XL U638 ( .A(n74), .B(n75), .C(n76), .D(n77), .S0(n578), .S1(n543), .Y(
        n173) );
  CLKMX2X4 U639 ( .A(n195), .B(n196), .S0(n512), .Y(tag[15]) );
  MXI4XL U640 ( .A(n114), .B(n115), .C(n116), .D(n117), .S0(n578), .S1(n542), 
        .Y(n183) );
  MXI4XL U641 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n580), .S1(n545), 
        .Y(n180) );
  MXI4XL U642 ( .A(n122), .B(n123), .C(n124), .D(n125), .S0(n580), .S1(n545), 
        .Y(n179) );
  BUFX8 U643 ( .A(n516), .Y(n518) );
  CLKBUFX4 U644 ( .A(n582), .Y(n559) );
  CLKBUFX2 U645 ( .A(n516), .Y(n519) );
  CLKBUFX4 U646 ( .A(n695), .Y(n706) );
  CLKBUFX4 U647 ( .A(n730), .Y(n741) );
  CLKBUFX4 U648 ( .A(n638), .Y(n651) );
  CLKBUFX4 U649 ( .A(n657), .Y(n670) );
  CLKBUFX4 U650 ( .A(n764), .Y(n777) );
  CLKBUFX4 U651 ( .A(n745), .Y(n758) );
  CLKBUFX4 U652 ( .A(n676), .Y(n689) );
  CLKBUFX4 U653 ( .A(n711), .Y(n724) );
  BUFX12 U654 ( .A(n468), .Y(n513) );
  BUFX4 U655 ( .A(N33), .Y(n468) );
  BUFX8 U656 ( .A(n583), .Y(n554) );
  CLKBUFX2 U657 ( .A(n551), .Y(n555) );
  BUFX8 U658 ( .A(N32), .Y(n549) );
  CLKBUFX2 U659 ( .A(N32), .Y(n548) );
  BUFX8 U660 ( .A(N33), .Y(n514) );
  BUFX20 U661 ( .A(n1263), .Y(mem_write) );
  CLKBUFX2 U662 ( .A(N31), .Y(n582) );
  AND2X1 U663 ( .A(n142), .B(N31), .Y(n143) );
  AND2XL U664 ( .A(N32), .B(N33), .Y(n142) );
  BUFX4 U665 ( .A(n1259), .Y(n630) );
  CLKINVX20 U666 ( .A(N33), .Y(n785) );
  NOR2X4 U667 ( .A(n815), .B(n814), .Y(n825) );
  INVX1 U668 ( .A(n1097), .Y(n1094) );
  MXI2XL U669 ( .A(tag[9]), .B(proc_addr[14]), .S0(n609), .Y(n1052) );
  INVXL U670 ( .A(tag[2]), .Y(n1065) );
  INVXL U671 ( .A(tag[3]), .Y(n1062) );
  INVXL U672 ( .A(blockdata[8]), .Y(n1142) );
  INVXL U673 ( .A(blockdata[0]), .Y(n1102) );
  INVXL U674 ( .A(blockdata[7]), .Y(n1137) );
  INVXL U675 ( .A(blockdata[16]), .Y(n1182) );
  INVXL U676 ( .A(blockdata[14]), .Y(n1172) );
  INVXL U677 ( .A(blockdata[15]), .Y(n1177) );
  INVXL U678 ( .A(blockdata[17]), .Y(n1187) );
  INVXL U679 ( .A(blockdata[18]), .Y(n1192) );
  INVXL U680 ( .A(blockdata[19]), .Y(n1197) );
  INVXL U681 ( .A(blockdata[20]), .Y(n1202) );
  INVXL U682 ( .A(blockdata[21]), .Y(n1207) );
  INVXL U683 ( .A(blockdata[22]), .Y(n1212) );
  INVXL U684 ( .A(blockdata[23]), .Y(n1217) );
  INVXL U685 ( .A(blockdata[24]), .Y(n1222) );
  INVXL U686 ( .A(blockdata[25]), .Y(n1227) );
  INVXL U687 ( .A(blockdata[26]), .Y(n1232) );
  INVXL U688 ( .A(blockdata[27]), .Y(n1237) );
  INVXL U689 ( .A(blockdata[28]), .Y(n1242) );
  INVXL U690 ( .A(blockdata[29]), .Y(n1247) );
  INVXL U691 ( .A(blockdata[30]), .Y(n1252) );
  INVXL U692 ( .A(blockdata[31]), .Y(n1260) );
  INVXL U693 ( .A(blockdata[9]), .Y(n1147) );
  INVXL U694 ( .A(blockdata[10]), .Y(n1152) );
  INVXL U695 ( .A(blockdata[11]), .Y(n1157) );
  INVXL U696 ( .A(blockdata[12]), .Y(n1162) );
  INVXL U697 ( .A(blockdata[13]), .Y(n1167) );
  INVXL U698 ( .A(blockdata[112]), .Y(n1181) );
  INVXL U699 ( .A(blockdata[104]), .Y(n1141) );
  INVXL U700 ( .A(blockdata[105]), .Y(n1146) );
  INVXL U701 ( .A(blockdata[106]), .Y(n1151) );
  INVXL U702 ( .A(blockdata[107]), .Y(n1156) );
  INVXL U703 ( .A(blockdata[108]), .Y(n1161) );
  INVXL U704 ( .A(blockdata[110]), .Y(n1171) );
  INVXL U705 ( .A(blockdata[111]), .Y(n1176) );
  INVXL U706 ( .A(blockdata[113]), .Y(n1186) );
  INVXL U707 ( .A(blockdata[114]), .Y(n1191) );
  INVXL U708 ( .A(blockdata[115]), .Y(n1196) );
  INVXL U709 ( .A(blockdata[116]), .Y(n1201) );
  INVXL U710 ( .A(blockdata[109]), .Y(n1166) );
  INVXL U711 ( .A(blockdata[97]), .Y(n1106) );
  INVXL U712 ( .A(blockdata[98]), .Y(n1111) );
  INVXL U713 ( .A(blockdata[99]), .Y(n1116) );
  INVXL U714 ( .A(blockdata[100]), .Y(n1121) );
  INVXL U715 ( .A(blockdata[101]), .Y(n1126) );
  INVXL U716 ( .A(blockdata[102]), .Y(n1131) );
  INVXL U717 ( .A(blockdata[103]), .Y(n1136) );
  INVXL U718 ( .A(blockdata[96]), .Y(n1101) );
  INVXL U719 ( .A(blockdata[118]), .Y(n1211) );
  INVXL U720 ( .A(blockdata[119]), .Y(n1216) );
  INVXL U721 ( .A(blockdata[120]), .Y(n1221) );
  INVXL U722 ( .A(blockdata[121]), .Y(n1226) );
  INVXL U723 ( .A(blockdata[122]), .Y(n1231) );
  INVXL U724 ( .A(blockdata[117]), .Y(n1206) );
  INVXL U725 ( .A(blockdata[123]), .Y(n1236) );
  INVXL U726 ( .A(blockdata[124]), .Y(n1241) );
  INVXL U727 ( .A(blockdata[125]), .Y(n1246) );
  INVXL U728 ( .A(blockdata[126]), .Y(n1251) );
  INVXL U729 ( .A(blockdata[127]), .Y(n1258) );
  INVXL U730 ( .A(blockdata[88]), .Y(n1219) );
  INVXL U731 ( .A(blockdata[89]), .Y(n1224) );
  INVXL U732 ( .A(blockdata[90]), .Y(n1229) );
  INVXL U733 ( .A(blockdata[91]), .Y(n1234) );
  INVXL U734 ( .A(blockdata[92]), .Y(n1239) );
  INVXL U735 ( .A(blockdata[93]), .Y(n1244) );
  INVXL U736 ( .A(blockdata[94]), .Y(n1249) );
  INVXL U737 ( .A(blockdata[95]), .Y(n1255) );
  INVXL U738 ( .A(blockdata[80]), .Y(n1179) );
  INVXL U739 ( .A(blockdata[72]), .Y(n1139) );
  INVXL U740 ( .A(blockdata[73]), .Y(n1144) );
  INVXL U741 ( .A(blockdata[74]), .Y(n1149) );
  INVXL U742 ( .A(blockdata[75]), .Y(n1154) );
  INVXL U743 ( .A(blockdata[76]), .Y(n1159) );
  INVXL U744 ( .A(blockdata[78]), .Y(n1169) );
  INVXL U745 ( .A(blockdata[79]), .Y(n1174) );
  INVXL U746 ( .A(blockdata[81]), .Y(n1184) );
  INVXL U747 ( .A(blockdata[82]), .Y(n1189) );
  INVXL U748 ( .A(blockdata[83]), .Y(n1194) );
  INVXL U749 ( .A(blockdata[84]), .Y(n1199) );
  INVXL U750 ( .A(blockdata[85]), .Y(n1204) );
  INVXL U751 ( .A(blockdata[86]), .Y(n1209) );
  INVXL U752 ( .A(blockdata[87]), .Y(n1214) );
  INVXL U753 ( .A(blockdata[66]), .Y(n1109) );
  INVXL U754 ( .A(blockdata[67]), .Y(n1114) );
  INVXL U755 ( .A(blockdata[68]), .Y(n1119) );
  INVXL U756 ( .A(blockdata[69]), .Y(n1124) );
  INVXL U757 ( .A(blockdata[70]), .Y(n1129) );
  INVXL U758 ( .A(blockdata[71]), .Y(n1134) );
  INVXL U759 ( .A(blockdata[65]), .Y(n1104) );
  INVXL U760 ( .A(blockdata[77]), .Y(n1164) );
  INVXL U761 ( .A(blockdata[64]), .Y(n1099) );
  INVXL U762 ( .A(blockdata[48]), .Y(n1178) );
  INVXL U763 ( .A(blockdata[40]), .Y(n1138) );
  INVXL U764 ( .A(blockdata[41]), .Y(n1143) );
  INVXL U765 ( .A(blockdata[42]), .Y(n1148) );
  INVXL U766 ( .A(blockdata[43]), .Y(n1153) );
  INVXL U767 ( .A(blockdata[44]), .Y(n1158) );
  INVXL U768 ( .A(blockdata[46]), .Y(n1168) );
  INVXL U769 ( .A(blockdata[47]), .Y(n1173) );
  INVXL U770 ( .A(blockdata[49]), .Y(n1183) );
  INVXL U771 ( .A(blockdata[50]), .Y(n1188) );
  INVXL U772 ( .A(blockdata[51]), .Y(n1193) );
  INVXL U773 ( .A(blockdata[52]), .Y(n1198) );
  INVXL U774 ( .A(blockdata[53]), .Y(n1203) );
  INVXL U775 ( .A(blockdata[54]), .Y(n1208) );
  INVXL U776 ( .A(blockdata[55]), .Y(n1213) );
  INVXL U777 ( .A(blockdata[56]), .Y(n1218) );
  INVXL U778 ( .A(blockdata[57]), .Y(n1223) );
  INVXL U779 ( .A(blockdata[58]), .Y(n1228) );
  INVXL U780 ( .A(blockdata[59]), .Y(n1233) );
  INVXL U781 ( .A(blockdata[60]), .Y(n1238) );
  INVXL U782 ( .A(blockdata[61]), .Y(n1243) );
  INVXL U783 ( .A(blockdata[62]), .Y(n1248) );
  INVXL U784 ( .A(blockdata[63]), .Y(n1253) );
  INVXL U785 ( .A(blockdata[45]), .Y(n1163) );
  INVXL U786 ( .A(blockdata[33]), .Y(n1103) );
  INVXL U787 ( .A(blockdata[34]), .Y(n1108) );
  INVXL U788 ( .A(blockdata[35]), .Y(n1113) );
  INVXL U789 ( .A(blockdata[36]), .Y(n1118) );
  INVXL U790 ( .A(blockdata[37]), .Y(n1123) );
  INVXL U791 ( .A(blockdata[38]), .Y(n1128) );
  INVXL U792 ( .A(blockdata[39]), .Y(n1133) );
  INVXL U793 ( .A(blockdata[32]), .Y(n1098) );
  CLKMX2X2 U794 ( .A(n155), .B(n156), .S0(n513), .Y(tag[5]) );
  MX4XL U795 ( .A(\blocktag[0][5] ), .B(\blocktag[1][5] ), .C(\blocktag[2][5] ), .D(\blocktag[3][5] ), .S0(n581), .S1(n546), .Y(n155) );
  MX4XL U796 ( .A(\blocktag[4][5] ), .B(\blocktag[5][5] ), .C(\blocktag[6][5] ), .D(\blocktag[7][5] ), .S0(n581), .S1(n546), .Y(n156) );
  MX4XL U797 ( .A(\blocktag[0][6] ), .B(\blocktag[1][6] ), .C(\blocktag[2][6] ), .D(\blocktag[3][6] ), .S0(n581), .S1(n545), .Y(n153) );
  MX4XL U798 ( .A(\blocktag[4][6] ), .B(\blocktag[5][6] ), .C(\blocktag[6][6] ), .D(\blocktag[7][6] ), .S0(n580), .S1(n545), .Y(n154) );
  MX4XL U799 ( .A(\blocktag[0][18] ), .B(\blocktag[1][18] ), .C(
        \blocktag[2][18] ), .D(\blocktag[3][18] ), .S0(n579), .S1(n543), .Y(
        n157) );
  MX4XL U800 ( .A(\blocktag[4][18] ), .B(\blocktag[5][18] ), .C(
        \blocktag[6][18] ), .D(\blocktag[7][18] ), .S0(n579), .S1(n543), .Y(
        n158) );
  MXI4XL U801 ( .A(n66), .B(n67), .C(n68), .D(n69), .S0(n581), .S1(n546), .Y(
        n161) );
  MXI4XL U802 ( .A(n70), .B(n71), .C(n72), .D(n73), .S0(n581), .S1(n546), .Y(
        n162) );
  CLKMX2X2 U803 ( .A(n163), .B(n164), .S0(n513), .Y(tag[9]) );
  MX4XL U804 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(\blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n580), .S1(n545), .Y(n163) );
  MX4XL U805 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(\blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n580), .S1(n545), .Y(n164) );
  MX2X2 U806 ( .A(n167), .B(n168), .S0(n512), .Y(tag[13]) );
  MX4XL U807 ( .A(\blocktag[0][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[3][13] ), .S0(n579), .S1(n544), .Y(
        n167) );
  MX4XL U808 ( .A(\blocktag[4][13] ), .B(\blocktag[5][13] ), .C(
        \blocktag[6][13] ), .D(\blocktag[7][13] ), .S0(n579), .S1(n544), .Y(
        n168) );
  MX4XL U809 ( .A(\blocktag[0][20] ), .B(\blocktag[1][20] ), .C(
        \blocktag[2][20] ), .D(\blocktag[3][20] ), .S0(n578), .S1(n543), .Y(
        n177) );
  MX4XL U810 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n578), .S1(n543), .Y(
        n178) );
  MX4XL U811 ( .A(\blocktag[0][16] ), .B(\blocktag[1][16] ), .C(
        \blocktag[2][16] ), .D(\blocktag[3][16] ), .S0(n579), .S1(n544), .Y(
        n181) );
  MX4XL U812 ( .A(\blocktag[4][16] ), .B(\blocktag[5][16] ), .C(
        \blocktag[6][16] ), .D(\blocktag[7][16] ), .S0(n579), .S1(n544), .Y(
        n182) );
  MX4XL U813 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(\blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n581), .S1(n546), .Y(n187) );
  MX4XL U814 ( .A(\blocktag[4][0] ), .B(\blocktag[5][0] ), .C(\blocktag[6][0] ), .D(\blocktag[7][0] ), .S0(n581), .S1(n546), .Y(n188) );
  MXI4X1 U815 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n579), .S1(n544), 
        .Y(n191) );
  MXI4X1 U816 ( .A(n110), .B(n111), .C(n112), .D(n113), .S0(n579), .S1(n544), 
        .Y(n192) );
  MX4XL U817 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n579), .S1(n544), .Y(
        n195) );
  MX4XL U818 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n579), .S1(n544), .Y(
        n196) );
  NAND2XL U819 ( .A(mem_rdata[105]), .B(n618), .Y(n858) );
  NAND2XL U820 ( .A(mem_rdata[118]), .B(n616), .Y(n845) );
  NAND2XL U821 ( .A(mem_rdata[72]), .B(n616), .Y(n894) );
  NAND2XL U822 ( .A(mem_rdata[79]), .B(n617), .Y(n887) );
  NAND2XL U823 ( .A(mem_rdata[40]), .B(n614), .Y(n928) );
  NAND2XL U824 ( .A(mem_rdata[53]), .B(n615), .Y(n915) );
  NAND2XL U825 ( .A(mem_rdata[32]), .B(n613), .Y(n936) );
  MXI4XL U826 ( .A(\block[4][9] ), .B(\block[5][9] ), .C(\block[6][9] ), .D(
        \block[7][9] ), .S0(n576), .S1(n540), .Y(n442) );
  MXI4XL U827 ( .A(\block[0][9] ), .B(\block[1][9] ), .C(\block[2][9] ), .D(
        \block[3][9] ), .S0(n576), .S1(n540), .Y(n441) );
  MXI4XL U828 ( .A(\block[4][10] ), .B(\block[5][10] ), .C(\block[6][10] ), 
        .D(\block[7][10] ), .S0(n576), .S1(n540), .Y(n440) );
  MXI4XL U829 ( .A(\block[0][10] ), .B(\block[1][10] ), .C(\block[2][10] ), 
        .D(\block[3][10] ), .S0(n576), .S1(n540), .Y(n439) );
  MXI4XL U830 ( .A(\block[4][11] ), .B(\block[5][11] ), .C(\block[6][11] ), 
        .D(\block[7][11] ), .S0(n576), .S1(n540), .Y(n438) );
  MXI4XL U831 ( .A(\block[0][11] ), .B(\block[1][11] ), .C(\block[2][11] ), 
        .D(\block[3][11] ), .S0(n576), .S1(n540), .Y(n437) );
  MXI2XL U832 ( .A(n471), .B(n1085), .S0(n1006), .Y(n487) );
  MXI2X1 U833 ( .A(n480), .B(n1084), .S0(n1075), .Y(n496) );
  MXI2X1 U834 ( .A(n481), .B(n1084), .S0(n1077), .Y(n497) );
  MXI2X1 U835 ( .A(n482), .B(n1084), .S0(n1079), .Y(n498) );
  MXI2X1 U836 ( .A(n483), .B(n1084), .S0(n1081), .Y(n499) );
  MXI2X1 U837 ( .A(n484), .B(n1084), .S0(n1083), .Y(n500) );
  MXI2X1 U838 ( .A(n485), .B(n1084), .S0(n146), .Y(n501) );
  MXI2X1 U839 ( .A(n486), .B(n1084), .S0(n143), .Y(n503) );
  CLKBUFX3 U840 ( .A(n520), .Y(n537) );
  CLKBUFX3 U841 ( .A(n548), .Y(n536) );
  CLKBUFX3 U842 ( .A(n548), .Y(n530) );
  CLKBUFX3 U843 ( .A(n521), .Y(n535) );
  CLKBUFX3 U844 ( .A(n548), .Y(n529) );
  CLKBUFX3 U845 ( .A(n515), .Y(n534) );
  CLKBUFX3 U846 ( .A(n521), .Y(n533) );
  CLKBUFX3 U847 ( .A(n548), .Y(n528) );
  CLKBUFX3 U848 ( .A(n521), .Y(n532) );
  CLKBUFX3 U849 ( .A(n520), .Y(n531) );
  CLKBUFX3 U850 ( .A(n521), .Y(n527) );
  CLKBUFX3 U851 ( .A(n518), .Y(n541) );
  CLKBUFX3 U852 ( .A(n521), .Y(n526) );
  CLKBUFX3 U853 ( .A(n519), .Y(n540) );
  CLKBUFX3 U854 ( .A(n515), .Y(n525) );
  CLKBUFX3 U855 ( .A(n519), .Y(n539) );
  CLKBUFX3 U856 ( .A(n515), .Y(n524) );
  CLKBUFX3 U857 ( .A(n520), .Y(n538) );
  CLKBUFX3 U858 ( .A(n514), .Y(n511) );
  CLKBUFX3 U859 ( .A(n556), .Y(n572) );
  CLKBUFX3 U860 ( .A(n550), .Y(n567) );
  CLKBUFX3 U861 ( .A(n557), .Y(n571) );
  CLKBUFX3 U862 ( .A(n582), .Y(n566) );
  CLKBUFX3 U863 ( .A(n557), .Y(n570) );
  CLKBUFX3 U864 ( .A(n557), .Y(n565) );
  CLKBUFX3 U865 ( .A(n556), .Y(n569) );
  CLKBUFX3 U866 ( .A(n550), .Y(n564) );
  CLKBUFX3 U867 ( .A(n550), .Y(n568) );
  CLKBUFX3 U868 ( .A(n557), .Y(n563) );
  CLKBUFX3 U869 ( .A(n555), .Y(n562) );
  CLKBUFX3 U870 ( .A(n554), .Y(n576) );
  CLKBUFX3 U871 ( .A(n557), .Y(n561) );
  CLKBUFX3 U872 ( .A(n555), .Y(n575) );
  CLKBUFX3 U873 ( .A(n550), .Y(n560) );
  CLKBUFX3 U874 ( .A(n555), .Y(n574) );
  CLKBUFX3 U875 ( .A(n556), .Y(n573) );
  CLKBUFX3 U876 ( .A(n550), .Y(n558) );
  CLKBUFX3 U877 ( .A(n467), .Y(n509) );
  CLKBUFX3 U878 ( .A(n466), .Y(n508) );
  CLKBUFX3 U879 ( .A(n466), .Y(n505) );
  CLKBUFX3 U880 ( .A(n466), .Y(n507) );
  CLKBUFX3 U881 ( .A(n465), .Y(n504) );
  CLKBUFX3 U882 ( .A(n466), .Y(n506) );
  CLKBUFX3 U883 ( .A(n465), .Y(n502) );
  CLKBUFX3 U884 ( .A(n467), .Y(n510) );
  CLKBUFX3 U885 ( .A(n781), .Y(n769) );
  CLKBUFX3 U886 ( .A(n781), .Y(n770) );
  CLKBUFX3 U887 ( .A(n780), .Y(n771) );
  CLKBUFX3 U888 ( .A(n780), .Y(n772) );
  CLKBUFX3 U889 ( .A(n779), .Y(n773) );
  CLKBUFX3 U890 ( .A(n779), .Y(n774) );
  CLKBUFX3 U891 ( .A(n764), .Y(n775) );
  CLKBUFX3 U892 ( .A(n764), .Y(n776) );
  CLKBUFX3 U893 ( .A(n762), .Y(n750) );
  CLKBUFX3 U894 ( .A(n762), .Y(n751) );
  CLKBUFX3 U895 ( .A(n761), .Y(n752) );
  CLKBUFX3 U896 ( .A(n761), .Y(n753) );
  CLKBUFX3 U897 ( .A(n760), .Y(n754) );
  CLKBUFX3 U898 ( .A(n760), .Y(n755) );
  CLKBUFX3 U899 ( .A(n745), .Y(n756) );
  CLKBUFX3 U900 ( .A(n745), .Y(n757) );
  CLKBUFX3 U901 ( .A(n744), .Y(n733) );
  CLKBUFX3 U902 ( .A(n744), .Y(n734) );
  CLKBUFX3 U903 ( .A(n730), .Y(n735) );
  CLKBUFX3 U904 ( .A(n730), .Y(n736) );
  CLKBUFX3 U905 ( .A(n743), .Y(n737) );
  CLKBUFX3 U906 ( .A(n743), .Y(n738) );
  CLKBUFX3 U907 ( .A(n743), .Y(n739) );
  CLKBUFX3 U908 ( .A(n743), .Y(n740) );
  CLKBUFX3 U909 ( .A(n728), .Y(n716) );
  CLKBUFX3 U910 ( .A(n728), .Y(n717) );
  CLKBUFX3 U911 ( .A(n727), .Y(n718) );
  CLKBUFX3 U912 ( .A(n727), .Y(n719) );
  CLKBUFX3 U913 ( .A(n726), .Y(n720) );
  CLKBUFX3 U914 ( .A(n726), .Y(n721) );
  CLKBUFX3 U915 ( .A(n711), .Y(n722) );
  CLKBUFX3 U916 ( .A(n711), .Y(n723) );
  CLKBUFX3 U917 ( .A(n708), .Y(n698) );
  CLKBUFX3 U918 ( .A(n708), .Y(n699) );
  CLKBUFX3 U919 ( .A(n710), .Y(n700) );
  CLKBUFX3 U920 ( .A(n710), .Y(n701) );
  CLKBUFX3 U921 ( .A(n709), .Y(n702) );
  CLKBUFX3 U922 ( .A(n709), .Y(n703) );
  CLKBUFX3 U923 ( .A(n708), .Y(n704) );
  CLKBUFX3 U924 ( .A(n708), .Y(n705) );
  CLKBUFX3 U925 ( .A(n693), .Y(n681) );
  CLKBUFX3 U926 ( .A(n693), .Y(n682) );
  CLKBUFX3 U927 ( .A(n692), .Y(n683) );
  CLKBUFX3 U928 ( .A(n692), .Y(n684) );
  CLKBUFX3 U929 ( .A(n691), .Y(n685) );
  CLKBUFX3 U930 ( .A(n691), .Y(n686) );
  CLKBUFX3 U931 ( .A(n676), .Y(n687) );
  CLKBUFX3 U932 ( .A(n676), .Y(n688) );
  CLKBUFX3 U933 ( .A(n674), .Y(n662) );
  CLKBUFX3 U934 ( .A(n674), .Y(n663) );
  CLKBUFX3 U935 ( .A(n673), .Y(n664) );
  CLKBUFX3 U936 ( .A(n673), .Y(n665) );
  CLKBUFX3 U937 ( .A(n672), .Y(n666) );
  CLKBUFX3 U938 ( .A(n672), .Y(n667) );
  CLKBUFX3 U939 ( .A(n657), .Y(n668) );
  CLKBUFX3 U940 ( .A(n657), .Y(n669) );
  CLKBUFX3 U941 ( .A(n655), .Y(n643) );
  CLKBUFX3 U942 ( .A(n655), .Y(n644) );
  CLKBUFX3 U943 ( .A(n654), .Y(n645) );
  CLKBUFX3 U944 ( .A(n654), .Y(n646) );
  CLKBUFX3 U945 ( .A(n653), .Y(n647) );
  CLKBUFX3 U946 ( .A(n653), .Y(n648) );
  CLKBUFX3 U947 ( .A(n638), .Y(n649) );
  CLKBUFX3 U948 ( .A(n638), .Y(n650) );
  CLKBUFX3 U949 ( .A(n782), .Y(n767) );
  CLKBUFX3 U950 ( .A(n782), .Y(n768) );
  CLKBUFX3 U951 ( .A(n763), .Y(n748) );
  CLKBUFX3 U952 ( .A(n763), .Y(n749) );
  CLKBUFX3 U953 ( .A(n744), .Y(n731) );
  CLKBUFX3 U954 ( .A(n744), .Y(n732) );
  CLKBUFX3 U955 ( .A(n729), .Y(n714) );
  CLKBUFX3 U956 ( .A(n729), .Y(n715) );
  CLKBUFX3 U957 ( .A(n695), .Y(n696) );
  CLKBUFX3 U958 ( .A(n695), .Y(n697) );
  CLKBUFX3 U959 ( .A(n694), .Y(n679) );
  CLKBUFX3 U960 ( .A(n694), .Y(n680) );
  CLKBUFX3 U961 ( .A(n675), .Y(n660) );
  CLKBUFX3 U962 ( .A(n675), .Y(n661) );
  CLKBUFX3 U963 ( .A(n656), .Y(n641) );
  CLKBUFX3 U964 ( .A(n656), .Y(n642) );
  CLKBUFX3 U965 ( .A(n764), .Y(n778) );
  CLKBUFX3 U966 ( .A(n745), .Y(n759) );
  CLKBUFX3 U967 ( .A(n730), .Y(n742) );
  CLKBUFX3 U968 ( .A(n711), .Y(n725) );
  CLKBUFX3 U969 ( .A(n695), .Y(n707) );
  CLKBUFX3 U970 ( .A(n676), .Y(n690) );
  CLKBUFX3 U971 ( .A(n657), .Y(n671) );
  CLKBUFX3 U972 ( .A(n638), .Y(n652) );
  CLKBUFX3 U973 ( .A(n549), .Y(n516) );
  CLKBUFX3 U974 ( .A(n465), .Y(n469) );
  CLKBUFX3 U975 ( .A(n515), .Y(n522) );
  CLKBUFX3 U976 ( .A(n766), .Y(n781) );
  CLKBUFX3 U977 ( .A(n747), .Y(n762) );
  CLKBUFX3 U978 ( .A(n136), .Y(n743) );
  CLKBUFX3 U979 ( .A(n713), .Y(n728) );
  CLKBUFX3 U980 ( .A(n138), .Y(n708) );
  CLKBUFX3 U981 ( .A(n678), .Y(n693) );
  CLKBUFX3 U982 ( .A(n659), .Y(n674) );
  CLKBUFX3 U983 ( .A(n640), .Y(n655) );
  CLKBUFX3 U984 ( .A(n766), .Y(n782) );
  CLKBUFX3 U985 ( .A(n747), .Y(n763) );
  CLKBUFX3 U986 ( .A(n713), .Y(n729) );
  CLKBUFX3 U987 ( .A(n678), .Y(n694) );
  CLKBUFX3 U988 ( .A(n659), .Y(n675) );
  CLKBUFX3 U989 ( .A(n640), .Y(n656) );
  CLKBUFX3 U990 ( .A(n134), .Y(n765) );
  CLKBUFX3 U991 ( .A(n135), .Y(n746) );
  CLKBUFX3 U992 ( .A(n137), .Y(n712) );
  CLKBUFX3 U993 ( .A(n139), .Y(n677) );
  CLKBUFX3 U994 ( .A(n140), .Y(n658) );
  CLKBUFX3 U995 ( .A(n141), .Y(n639) );
  CLKBUFX3 U996 ( .A(n134), .Y(n766) );
  CLKBUFX3 U997 ( .A(n135), .Y(n747) );
  CLKBUFX3 U998 ( .A(n137), .Y(n713) );
  CLKBUFX3 U999 ( .A(n138), .Y(n695) );
  CLKBUFX3 U1000 ( .A(n139), .Y(n678) );
  CLKBUFX3 U1001 ( .A(n140), .Y(n659) );
  CLKBUFX3 U1002 ( .A(n141), .Y(n640) );
  CLKBUFX3 U1003 ( .A(n134), .Y(n764) );
  CLKBUFX3 U1004 ( .A(n135), .Y(n745) );
  CLKBUFX3 U1005 ( .A(n136), .Y(n730) );
  CLKBUFX3 U1006 ( .A(n137), .Y(n711) );
  CLKBUFX3 U1007 ( .A(n139), .Y(n676) );
  CLKBUFX3 U1008 ( .A(n140), .Y(n657) );
  CLKBUFX3 U1009 ( .A(n141), .Y(n638) );
  CLKBUFX3 U1010 ( .A(n514), .Y(n467) );
  CLKBUFX3 U1011 ( .A(n514), .Y(n466) );
  CLKBUFX3 U1012 ( .A(n514), .Y(n465) );
  CLKBUFX3 U1013 ( .A(N32), .Y(n547) );
  CLKBUFX6 U1014 ( .A(n786), .Y(n789) );
  CLKBUFX6 U1015 ( .A(n786), .Y(n788) );
  CLKBUFX3 U1016 ( .A(n588), .Y(n586) );
  CLKBUFX3 U1017 ( .A(n588), .Y(n587) );
  CLKBUFX3 U1018 ( .A(n591), .Y(n593) );
  CLKBUFX3 U1019 ( .A(n591), .Y(n592) );
  INVX3 U1020 ( .A(n55), .Y(n599) );
  INVX3 U1021 ( .A(n601), .Y(n598) );
  CLKBUFX3 U1022 ( .A(n1263), .Y(n786) );
  CLKBUFX3 U1023 ( .A(n604), .Y(n607) );
  CLKBUFX3 U1024 ( .A(n1261), .Y(n636) );
  CLKBUFX3 U1025 ( .A(n1261), .Y(n637) );
  CLKBUFX3 U1026 ( .A(n1254), .Y(n624) );
  CLKBUFX3 U1027 ( .A(n1254), .Y(n625) );
  CLKBUFX3 U1028 ( .A(n1259), .Y(n631) );
  CLKINVX1 U1029 ( .A(n836), .Y(n1006) );
  NAND3BXL U1030 ( .AN(N32), .B(n783), .C(n785), .Y(n836) );
  CLKINVX1 U1031 ( .A(n1074), .Y(n1075) );
  NAND3BXL U1032 ( .AN(N32), .B(N31), .C(n785), .Y(n1074) );
  CLKINVX1 U1033 ( .A(n1076), .Y(n1077) );
  NAND3BXL U1034 ( .AN(N31), .B(N32), .C(n785), .Y(n1076) );
  CLKINVX1 U1035 ( .A(n1078), .Y(n1079) );
  NAND3BXL U1036 ( .AN(n784), .B(N31), .C(n785), .Y(n1078) );
  CLKINVX1 U1037 ( .A(n1080), .Y(n1081) );
  NAND3BXL U1038 ( .AN(N31), .B(N33), .C(n784), .Y(n1080) );
  CLKINVX1 U1039 ( .A(n1082), .Y(n1083) );
  NAND3BXL U1040 ( .AN(n785), .B(N31), .C(n784), .Y(n1082) );
  AND2X2 U1041 ( .A(n142), .B(n783), .Y(n146) );
  CLKBUFX3 U1042 ( .A(n793), .Y(n791) );
  CLKBUFX3 U1043 ( .A(n605), .Y(n608) );
  CLKBUFX3 U1044 ( .A(n1), .Y(n605) );
  NAND2X1 U1045 ( .A(n152), .B(n1094), .Y(n1259) );
  CLKBUFX3 U1046 ( .A(n1261), .Y(n635) );
  CLKBUFX3 U1047 ( .A(n627), .Y(n626) );
  CLKBUFX3 U1048 ( .A(n1254), .Y(n623) );
  CLKINVX1 U1049 ( .A(proc_reset), .Y(n793) );
  NAND2X2 U1050 ( .A(n806), .B(n805), .Y(n807) );
  NAND4X2 U1051 ( .A(n797), .B(n796), .C(n795), .D(n794), .Y(n801) );
  NAND4BX2 U1052 ( .AN(n149), .B(n804), .C(n803), .D(n802), .Y(n808) );
  XOR2X2 U1053 ( .A(n1050), .B(proc_addr[15]), .Y(n810) );
  CLKINVX1 U1054 ( .A(tag[16]), .Y(n1032) );
  CLKINVX1 U1055 ( .A(tag[13]), .Y(n1041) );
  CLKINVX1 U1056 ( .A(tag[17]), .Y(n1029) );
  CLKBUFX12 U1057 ( .A(n1262), .Y(mem_read) );
  NAND2XL U1058 ( .A(n1090), .B(n1092), .Y(n1091) );
  AO22X1 U1059 ( .A0(proc_addr[10]), .A1(mem_read), .B0(tag[5]), .B1(mem_write), .Y(mem_addr[8]) );
  AO22X1 U1060 ( .A0(proc_addr[15]), .A1(mem_read), .B0(tag[10]), .B1(
        mem_write), .Y(mem_addr[13]) );
  INVXL U1061 ( .A(proc_addr[18]), .Y(n1040) );
  MX2XL U1062 ( .A(n1032), .B(n1031), .S0(n610), .Y(n1033) );
  INVXL U1063 ( .A(proc_addr[21]), .Y(n1031) );
  INVXL U1064 ( .A(proc_addr[25]), .Y(n1019) );
  MX2XL U1065 ( .A(n1014), .B(n1013), .S0(n610), .Y(n1015) );
  INVXL U1066 ( .A(proc_addr[28]), .Y(n1010) );
  MX2XL U1067 ( .A(n1008), .B(n1007), .S0(n610), .Y(n1009) );
  INVXL U1068 ( .A(proc_addr[29]), .Y(n1007) );
  NAND2XL U1069 ( .A(n204), .B(proc_stall), .Y(n834) );
  INVXL U1070 ( .A(proc_addr[5]), .Y(n1071) );
  INVXL U1071 ( .A(proc_addr[13]), .Y(n1053) );
  INVXL U1072 ( .A(proc_addr[15]), .Y(n1049) );
  MX2XL U1073 ( .A(n1047), .B(n1046), .S0(n609), .Y(n1048) );
  INVXL U1074 ( .A(proc_addr[16]), .Y(n1046) );
  MX2XL U1075 ( .A(n1044), .B(n1043), .S0(n609), .Y(n1045) );
  INVXL U1076 ( .A(proc_addr[17]), .Y(n1043) );
  BUFX4 U1077 ( .A(n1256), .Y(n627) );
  INVX1 U1078 ( .A(proc_addr[1]), .Y(n1096) );
  AND2XL U1079 ( .A(proc_addr[0]), .B(proc_addr[1]), .Y(n152) );
  CLKMX2X4 U1080 ( .A(n161), .B(n162), .S0(n513), .Y(tag[4]) );
  MX4X1 U1081 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(
        \blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n581), .S1(n546), .Y(n165) );
  MX4X1 U1082 ( .A(\blocktag[4][2] ), .B(\blocktag[5][2] ), .C(
        \blocktag[6][2] ), .D(\blocktag[7][2] ), .S0(n581), .S1(n546), .Y(n166) );
  CLKMX2X4 U1083 ( .A(n175), .B(n176), .S0(n513), .Y(tag[11]) );
  MX4X1 U1084 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n580), .S1(n545), .Y(
        n175) );
  MX4X1 U1085 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n580), .S1(n545), .Y(
        n176) );
  CLKMX2X4 U1086 ( .A(n179), .B(n180), .S0(n513), .Y(tag[10]) );
  CLKMX2X4 U1087 ( .A(n183), .B(n184), .S0(n511), .Y(tag[24]) );
  MX4X1 U1088 ( .A(\blocktag[0][21] ), .B(\blocktag[1][21] ), .C(
        \blocktag[2][21] ), .D(\blocktag[3][21] ), .S0(n578), .S1(n543), .Y(
        n189) );
  MX4X1 U1089 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n579), .S1(n544), .Y(
        n197) );
  MX4X1 U1090 ( .A(\blocktag[0][7] ), .B(\blocktag[1][7] ), .C(
        \blocktag[2][7] ), .D(\blocktag[3][7] ), .S0(n580), .S1(n545), .Y(n199) );
  MX4X1 U1091 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(
        \blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n581), .S1(n546), .Y(n201) );
  NAND2XL U1092 ( .A(mem_rdata[41]), .B(n614), .Y(n927) );
  NAND2XL U1093 ( .A(mem_rdata[42]), .B(n614), .Y(n926) );
  NAND2XL U1094 ( .A(mem_rdata[43]), .B(n614), .Y(n925) );
  NAND2XL U1095 ( .A(mem_rdata[44]), .B(n614), .Y(n924) );
  NAND2XL U1096 ( .A(mem_rdata[45]), .B(n614), .Y(n923) );
  NAND2XL U1097 ( .A(mem_rdata[46]), .B(n614), .Y(n922) );
  NAND2XL U1098 ( .A(mem_rdata[47]), .B(n614), .Y(n921) );
  NAND2XL U1099 ( .A(mem_rdata[49]), .B(n614), .Y(n919) );
  NAND2XL U1100 ( .A(mem_rdata[50]), .B(n614), .Y(n918) );
  NAND2XL U1101 ( .A(mem_rdata[51]), .B(n614), .Y(n917) );
  NAND2XL U1102 ( .A(mem_rdata[52]), .B(n614), .Y(n916) );
  NAND2XL U1103 ( .A(mem_rdata[54]), .B(n615), .Y(n914) );
  NAND2XL U1104 ( .A(mem_rdata[55]), .B(n615), .Y(n913) );
  NAND2XL U1105 ( .A(mem_rdata[56]), .B(n615), .Y(n912) );
  NAND2XL U1106 ( .A(mem_rdata[57]), .B(n615), .Y(n911) );
  NAND2XL U1107 ( .A(mem_rdata[58]), .B(n615), .Y(n910) );
  NAND2XL U1108 ( .A(mem_rdata[59]), .B(n615), .Y(n909) );
  NAND2XL U1109 ( .A(mem_rdata[60]), .B(n615), .Y(n908) );
  NAND2XL U1110 ( .A(mem_rdata[61]), .B(n615), .Y(n907) );
  NAND2XL U1111 ( .A(mem_rdata[62]), .B(n615), .Y(n906) );
  NAND2XL U1112 ( .A(mem_rdata[63]), .B(n615), .Y(n905) );
  NAND2XL U1113 ( .A(mem_rdata[33]), .B(n613), .Y(n935) );
  NAND2XL U1114 ( .A(mem_rdata[34]), .B(n613), .Y(n934) );
  NAND2XL U1115 ( .A(mem_rdata[35]), .B(n613), .Y(n933) );
  NAND2XL U1116 ( .A(mem_rdata[36]), .B(n613), .Y(n932) );
  NAND2XL U1117 ( .A(mem_rdata[37]), .B(n613), .Y(n931) );
  NAND2XL U1118 ( .A(mem_rdata[38]), .B(n613), .Y(n930) );
  NAND2XL U1119 ( .A(mem_rdata[39]), .B(n613), .Y(n929) );
  NAND2XL U1120 ( .A(mem_rdata[73]), .B(n616), .Y(n893) );
  NAND2XL U1121 ( .A(mem_rdata[74]), .B(n616), .Y(n892) );
  NAND2XL U1122 ( .A(mem_rdata[75]), .B(n616), .Y(n891) );
  NAND2XL U1123 ( .A(mem_rdata[78]), .B(n616), .Y(n888) );
  NAND2XL U1124 ( .A(mem_rdata[81]), .B(n617), .Y(n885) );
  NAND2XL U1125 ( .A(mem_rdata[82]), .B(n617), .Y(n884) );
  NAND2XL U1126 ( .A(mem_rdata[83]), .B(n617), .Y(n883) );
  NAND2XL U1127 ( .A(mem_rdata[84]), .B(n617), .Y(n882) );
  NAND2XL U1128 ( .A(mem_rdata[85]), .B(n617), .Y(n881) );
  NAND2XL U1129 ( .A(mem_rdata[86]), .B(n617), .Y(n880) );
  NAND2XL U1130 ( .A(mem_rdata[87]), .B(n617), .Y(n879) );
  NAND2XL U1131 ( .A(mem_rdata[88]), .B(n617), .Y(n878) );
  NAND2XL U1132 ( .A(mem_rdata[89]), .B(n617), .Y(n877) );
  NAND2XL U1133 ( .A(mem_rdata[90]), .B(n617), .Y(n876) );
  NAND2XL U1134 ( .A(mem_rdata[91]), .B(n617), .Y(n875) );
  NAND2XL U1135 ( .A(mem_rdata[95]), .B(n612), .Y(n871) );
  NAND2XL U1136 ( .A(mem_rdata[64]), .B(n615), .Y(n902) );
  NAND2XL U1137 ( .A(mem_rdata[65]), .B(n615), .Y(n901) );
  NAND2XL U1138 ( .A(mem_rdata[66]), .B(n616), .Y(n900) );
  NAND2XL U1139 ( .A(mem_rdata[67]), .B(n616), .Y(n899) );
  NAND2XL U1140 ( .A(mem_rdata[68]), .B(n616), .Y(n898) );
  NAND2XL U1141 ( .A(mem_rdata[69]), .B(n616), .Y(n897) );
  NAND2XL U1142 ( .A(mem_rdata[70]), .B(n616), .Y(n896) );
  NAND2XL U1143 ( .A(mem_rdata[71]), .B(n616), .Y(n895) );
  NAND2XL U1144 ( .A(mem_rdata[106]), .B(n618), .Y(n857) );
  NAND2XL U1145 ( .A(mem_rdata[107]), .B(n618), .Y(n856) );
  NAND2XL U1146 ( .A(mem_rdata[108]), .B(n618), .Y(n855) );
  NAND2XL U1147 ( .A(mem_rdata[109]), .B(n618), .Y(n854) );
  NAND2XL U1148 ( .A(mem_rdata[110]), .B(n618), .Y(n853) );
  NAND2XL U1149 ( .A(mem_rdata[111]), .B(n618), .Y(n852) );
  NAND2XL U1150 ( .A(mem_rdata[113]), .B(n618), .Y(n850) );
  NAND2XL U1151 ( .A(mem_rdata[114]), .B(n618), .Y(n849) );
  NAND2XL U1152 ( .A(mem_rdata[115]), .B(n618), .Y(n848) );
  NAND2XL U1153 ( .A(mem_rdata[116]), .B(n618), .Y(n847) );
  NAND2XL U1154 ( .A(mem_rdata[117]), .B(n618), .Y(n846) );
  NAND2XL U1155 ( .A(mem_rdata[120]), .B(n616), .Y(n843) );
  NAND2XL U1156 ( .A(mem_rdata[121]), .B(n616), .Y(n842) );
  NAND2XL U1157 ( .A(mem_rdata[122]), .B(n616), .Y(n841) );
  NAND2XL U1158 ( .A(mem_rdata[123]), .B(n616), .Y(n840) );
  NAND2XL U1159 ( .A(mem_rdata[124]), .B(n616), .Y(n839) );
  NAND2XL U1160 ( .A(mem_rdata[125]), .B(n616), .Y(n838) );
  NAND2XL U1161 ( .A(mem_rdata[126]), .B(n616), .Y(n837) );
  NAND2XL U1162 ( .A(mem_rdata[127]), .B(n616), .Y(n835) );
  NAND2XL U1163 ( .A(mem_rdata[100]), .B(n616), .Y(n863) );
  NAND2XL U1164 ( .A(mem_rdata[101]), .B(n616), .Y(n862) );
  NAND2XL U1165 ( .A(mem_rdata[102]), .B(n616), .Y(n861) );
  NAND2XL U1166 ( .A(mem_rdata[103]), .B(n611), .Y(n860) );
  NAND2XL U1167 ( .A(mem_rdata[48]), .B(n614), .Y(n920) );
  NAND2XL U1168 ( .A(mem_rdata[80]), .B(n617), .Y(n886) );
  NAND2XL U1169 ( .A(mem_rdata[112]), .B(n618), .Y(n851) );
  NAND2XL U1170 ( .A(mem_rdata[22]), .B(n612), .Y(n955) );
  NAND2XL U1171 ( .A(mem_rdata[23]), .B(n612), .Y(n953) );
  NAND2XL U1172 ( .A(mem_rdata[24]), .B(n612), .Y(n951) );
  NAND2XL U1173 ( .A(mem_rdata[25]), .B(n612), .Y(n949) );
  NAND2XL U1174 ( .A(mem_rdata[26]), .B(n612), .Y(n947) );
  NAND2XL U1175 ( .A(mem_rdata[27]), .B(n613), .Y(n945) );
  NAND2XL U1176 ( .A(mem_rdata[28]), .B(n613), .Y(n943) );
  NAND2XL U1177 ( .A(mem_rdata[29]), .B(n613), .Y(n941) );
  NAND2XL U1178 ( .A(mem_rdata[30]), .B(n613), .Y(n939) );
  NAND2XL U1179 ( .A(mem_rdata[31]), .B(n613), .Y(n937) );
  NAND2XL U1180 ( .A(mem_rdata[2]), .B(n611), .Y(n995) );
  NAND2XL U1181 ( .A(mem_rdata[3]), .B(n611), .Y(n993) );
  NAND2XL U1182 ( .A(mem_rdata[4]), .B(n611), .Y(n991) );
  NAND2XL U1183 ( .A(mem_rdata[5]), .B(n611), .Y(n989) );
  NAND2XL U1184 ( .A(mem_rdata[6]), .B(n611), .Y(n987) );
  MXI4XL U1185 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n577), .S1(n542), .Y(n461) );
  MXI4XL U1186 ( .A(blockvalid[4]), .B(blockvalid[5]), .C(blockvalid[6]), .D(
        blockvalid[7]), .S0(n577), .S1(n542), .Y(n462) );
  MXI2X1 U1187 ( .A(n463), .B(n464), .S0(n511), .Y(dirty) );
  MXI4XL U1188 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n578), .S1(n542), .Y(n463) );
  MXI4XL U1189 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n578), .S1(n542), .Y(n464) );
  AOI2BB1XL U1190 ( .A0N(n828), .A1N(n204), .B0(n203), .Y(n829) );
  INVXL U1191 ( .A(tag[18]), .Y(n1026) );
  INVXL U1192 ( .A(proc_addr[23]), .Y(n1025) );
  INVXL U1193 ( .A(proc_addr[26]), .Y(n1016) );
  INVXL U1194 ( .A(proc_addr[22]), .Y(n1028) );
  MXI2XL U1195 ( .A(n472), .B(n1085), .S0(n1075), .Y(n488) );
  MXI2XL U1196 ( .A(n473), .B(n1085), .S0(n1077), .Y(n489) );
  MXI2XL U1197 ( .A(n474), .B(n1085), .S0(n1079), .Y(n490) );
  MXI2XL U1198 ( .A(n475), .B(n1085), .S0(n1081), .Y(n491) );
  MXI2XL U1199 ( .A(n476), .B(n1085), .S0(n1083), .Y(n492) );
  MXI2XL U1200 ( .A(n477), .B(n1085), .S0(n146), .Y(n493) );
  MXI2XL U1201 ( .A(n478), .B(n1085), .S0(n143), .Y(n494) );
  MXI2X1 U1202 ( .A(n225), .B(n226), .S0(n469), .Y(blockdata[117]) );
  MXI4X1 U1203 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n559), .S1(n523), .Y(n226) );
  MXI4X1 U1204 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n559), .S1(n523), .Y(n225) );
  MXI2X1 U1205 ( .A(n223), .B(n224), .S0(n469), .Y(blockdata[118]) );
  MXI4X1 U1206 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n559), .S1(n523), .Y(n224) );
  MXI4X1 U1207 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n559), .S1(n523), .Y(n223) );
  MXI2X1 U1208 ( .A(n221), .B(n222), .S0(n469), .Y(blockdata[119]) );
  MXI4X1 U1209 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n559), .S1(n523), .Y(n222) );
  MXI4X1 U1210 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n559), .S1(n523), .Y(n221) );
  MXI2X1 U1211 ( .A(n219), .B(n220), .S0(n469), .Y(blockdata[120]) );
  MXI4X1 U1212 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n559), .S1(n523), .Y(n220) );
  MXI4X1 U1213 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n559), .S1(n523), .Y(n219) );
  MXI2X1 U1214 ( .A(n217), .B(n218), .S0(n469), .Y(blockdata[121]) );
  MXI4X1 U1215 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n559), .S1(n523), .Y(n218) );
  MXI4X1 U1216 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n559), .S1(n523), .Y(n217) );
  MXI2X1 U1217 ( .A(n215), .B(n216), .S0(n469), .Y(blockdata[122]) );
  MXI4X1 U1218 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n558), .S1(n523), .Y(n216) );
  MXI4X1 U1219 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n559), .S1(n523), .Y(n215) );
  AND2XL U1220 ( .A(mem_ready), .B(n1089), .Y(n204) );
  INVXL U1221 ( .A(proc_addr[19]), .Y(n1037) );
  MX2XL U1222 ( .A(n1023), .B(n1022), .S0(n610), .Y(n1024) );
  INVXL U1223 ( .A(proc_addr[24]), .Y(n1022) );
  MXI2X1 U1224 ( .A(n427), .B(n428), .S0(n510), .Y(blockdata[16]) );
  MXI4X1 U1225 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n575), .S1(n539), .Y(n428) );
  MXI4X1 U1226 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n575), .S1(n539), .Y(n427) );
  MXI2X1 U1227 ( .A(n433), .B(n434), .S0(n510), .Y(blockdata[13]) );
  MXI4X1 U1228 ( .A(\block[4][13] ), .B(\block[5][13] ), .C(\block[6][13] ), 
        .D(\block[7][13] ), .S0(n575), .S1(n540), .Y(n434) );
  MXI4X1 U1229 ( .A(\block[0][13] ), .B(\block[1][13] ), .C(\block[2][13] ), 
        .D(\block[3][13] ), .S0(n575), .S1(n540), .Y(n433) );
  MXI2X1 U1230 ( .A(n431), .B(n432), .S0(n510), .Y(blockdata[14]) );
  MXI4X1 U1231 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), 
        .D(\block[7][14] ), .S0(n575), .S1(n540), .Y(n432) );
  MXI4X1 U1232 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), 
        .D(\block[3][14] ), .S0(n575), .S1(n540), .Y(n431) );
  MXI2X1 U1233 ( .A(n429), .B(n430), .S0(n510), .Y(blockdata[15]) );
  MXI4X1 U1234 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n575), .S1(n539), .Y(n430) );
  MXI4X1 U1235 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n575), .S1(n539), .Y(n429) );
  MXI2X1 U1236 ( .A(n425), .B(n426), .S0(n510), .Y(blockdata[17]) );
  MXI4X1 U1237 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n575), .S1(n539), .Y(n426) );
  MXI4X1 U1238 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n575), .S1(n539), .Y(n425) );
  MXI2X1 U1239 ( .A(n423), .B(n424), .S0(n510), .Y(blockdata[18]) );
  MXI4X1 U1240 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n574), .S1(n539), .Y(n424) );
  MXI4X1 U1241 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n575), .S1(n539), .Y(n423) );
  MXI2X1 U1242 ( .A(n421), .B(n422), .S0(n510), .Y(blockdata[19]) );
  MXI4X1 U1243 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n574), .S1(n539), .Y(n422) );
  MXI4X1 U1244 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n574), .S1(n539), .Y(n421) );
  MXI2X1 U1245 ( .A(n419), .B(n420), .S0(n510), .Y(blockdata[20]) );
  MXI4X1 U1246 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n574), .S1(n539), .Y(n420) );
  MXI4X1 U1247 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n574), .S1(n539), .Y(n419) );
  MXI2X1 U1248 ( .A(n417), .B(n418), .S0(n509), .Y(blockdata[21]) );
  MXI4X1 U1249 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n574), .S1(n538), .Y(n418) );
  MXI4X1 U1250 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n574), .S1(n538), .Y(n417) );
  MXI2X1 U1251 ( .A(n415), .B(n416), .S0(n509), .Y(blockdata[22]) );
  MXI4X1 U1252 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n574), .S1(n538), .Y(n416) );
  MXI4X1 U1253 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n574), .S1(n538), .Y(n415) );
  MXI2X1 U1254 ( .A(n413), .B(n414), .S0(n509), .Y(blockdata[23]) );
  MXI4X1 U1255 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n574), .S1(n538), .Y(n414) );
  MXI4X1 U1256 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n574), .S1(n538), .Y(n413) );
  MXI2X1 U1257 ( .A(n411), .B(n412), .S0(n509), .Y(blockdata[24]) );
  MXI4X1 U1258 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n574), .S1(n538), .Y(n412) );
  MXI4X1 U1259 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n574), .S1(n538), .Y(n411) );
  MXI2XL U1260 ( .A(n459), .B(n460), .S0(n511), .Y(blockdata[0]) );
  MXI4XL U1261 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n577), .S1(n542), .Y(n460) );
  MXI4XL U1262 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n577), .S1(n542), .Y(n459) );
  MXI2X1 U1263 ( .A(n405), .B(n406), .S0(n509), .Y(blockdata[27]) );
  MXI4X1 U1264 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), 
        .D(\block[7][27] ), .S0(n573), .S1(n537), .Y(n406) );
  MXI4X1 U1265 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), 
        .D(\block[3][27] ), .S0(n573), .S1(n537), .Y(n405) );
  MXI2X1 U1266 ( .A(n403), .B(n404), .S0(n509), .Y(blockdata[28]) );
  MXI4X1 U1267 ( .A(\block[4][28] ), .B(\block[5][28] ), .C(\block[6][28] ), 
        .D(\block[7][28] ), .S0(n573), .S1(n537), .Y(n404) );
  MXI4X1 U1268 ( .A(\block[0][28] ), .B(\block[1][28] ), .C(\block[2][28] ), 
        .D(\block[3][28] ), .S0(n573), .S1(n537), .Y(n403) );
  MXI2X1 U1269 ( .A(n401), .B(n402), .S0(n509), .Y(blockdata[29]) );
  MXI4X1 U1270 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n573), .S1(n537), .Y(n402) );
  MXI4X1 U1271 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n573), .S1(n537), .Y(n401) );
  MXI2X1 U1272 ( .A(n399), .B(n400), .S0(n509), .Y(blockdata[30]) );
  MXI4X1 U1273 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n573), .S1(n537), .Y(n400) );
  MXI4X1 U1274 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n573), .S1(n537), .Y(n399) );
  MXI2X1 U1275 ( .A(n397), .B(n398), .S0(n509), .Y(blockdata[31]) );
  MXI4X1 U1276 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n572), .S1(n537), .Y(n398) );
  MXI4X1 U1277 ( .A(\block[0][31] ), .B(\block[1][31] ), .C(\block[2][31] ), 
        .D(\block[3][31] ), .S0(n573), .S1(n537), .Y(n397) );
  MXI2X1 U1278 ( .A(n409), .B(n410), .S0(n509), .Y(blockdata[25]) );
  MXI4X1 U1279 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n573), .S1(n538), .Y(n410) );
  MXI4X1 U1280 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n573), .S1(n538), .Y(n409) );
  MXI2X1 U1281 ( .A(n407), .B(n408), .S0(n509), .Y(blockdata[26]) );
  MXI4X1 U1282 ( .A(\block[4][26] ), .B(\block[5][26] ), .C(\block[6][26] ), 
        .D(\block[7][26] ), .S0(n573), .S1(n538), .Y(n408) );
  MXI4X1 U1283 ( .A(\block[0][26] ), .B(\block[1][26] ), .C(\block[2][26] ), 
        .D(\block[3][26] ), .S0(n573), .S1(n538), .Y(n407) );
  MXI2XL U1284 ( .A(n443), .B(n444), .S0(n511), .Y(blockdata[8]) );
  MXI4X1 U1285 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n576), .S1(n541), .Y(n444) );
  MXI4X1 U1286 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n576), .S1(n541), .Y(n443) );
  MXI2X1 U1287 ( .A(n441), .B(n442), .S0(n510), .Y(blockdata[9]) );
  MXI2X1 U1288 ( .A(n439), .B(n440), .S0(n510), .Y(blockdata[10]) );
  MXI2X1 U1289 ( .A(n437), .B(n438), .S0(n510), .Y(blockdata[11]) );
  MXI2X1 U1290 ( .A(n435), .B(n436), .S0(n510), .Y(blockdata[12]) );
  MXI4X1 U1291 ( .A(\block[4][12] ), .B(\block[5][12] ), .C(\block[6][12] ), 
        .D(\block[7][12] ), .S0(n575), .S1(n540), .Y(n436) );
  MXI4X1 U1292 ( .A(\block[0][12] ), .B(\block[1][12] ), .C(\block[2][12] ), 
        .D(\block[3][12] ), .S0(n575), .S1(n540), .Y(n435) );
  MXI4XL U1293 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n577), .S1(n542), .Y(n458) );
  MXI4XL U1294 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n577), .S1(n542), .Y(n457) );
  MXI4XL U1295 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n577), .S1(n542), .Y(n456) );
  MXI4XL U1296 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n577), .S1(n542), .Y(n455) );
  MXI4X1 U1297 ( .A(\block[4][5] ), .B(\block[5][5] ), .C(\block[6][5] ), .D(
        \block[7][5] ), .S0(n576), .S1(n541), .Y(n450) );
  MXI4X1 U1298 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n576), .S1(n541), .Y(n448) );
  MXI4X1 U1299 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n576), .S1(n541), .Y(n447) );
  MXI2XL U1300 ( .A(n445), .B(n446), .S0(n511), .Y(blockdata[7]) );
  MXI4X1 U1301 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n576), .S1(n541), .Y(n446) );
  MXI4X1 U1302 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n576), .S1(n541), .Y(n445) );
  MXI2X1 U1303 ( .A(n395), .B(n396), .S0(n509), .Y(blockdata[32]) );
  MXI4X1 U1304 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n572), .S1(n537), .Y(n396) );
  MXI4X1 U1305 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n572), .S1(n537), .Y(n395) );
  MXI2X1 U1306 ( .A(n331), .B(n332), .S0(n506), .Y(blockdata[64]) );
  MXI4X1 U1307 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n567), .S1(n531), .Y(n332) );
  MXI4X1 U1308 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n567), .S1(n531), .Y(n331) );
  MXI2X1 U1309 ( .A(n393), .B(n394), .S0(n508), .Y(blockdata[33]) );
  MXI4X1 U1310 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n572), .S1(n536), .Y(n394) );
  MXI4X1 U1311 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n572), .S1(n536), .Y(n393) );
  MXI2X1 U1312 ( .A(n329), .B(n330), .S0(n506), .Y(blockdata[65]) );
  MXI4X1 U1313 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n567), .S1(n531), .Y(n330) );
  MXI4X1 U1314 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n567), .S1(n531), .Y(n329) );
  MXI2X1 U1315 ( .A(n391), .B(n392), .S0(n508), .Y(blockdata[34]) );
  MXI4X1 U1316 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n572), .S1(n536), .Y(n392) );
  MXI4X1 U1317 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n572), .S1(n536), .Y(n391) );
  MXI2X1 U1318 ( .A(n327), .B(n328), .S0(n506), .Y(blockdata[66]) );
  MXI4X1 U1319 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n567), .S1(n531), .Y(n328) );
  MXI4X1 U1320 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n567), .S1(n531), .Y(n327) );
  MXI2X1 U1321 ( .A(n389), .B(n390), .S0(n508), .Y(blockdata[35]) );
  MXI4X1 U1322 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n572), .S1(n536), .Y(n390) );
  MXI4X1 U1323 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n572), .S1(n536), .Y(n389) );
  MXI2X1 U1324 ( .A(n325), .B(n326), .S0(n506), .Y(blockdata[67]) );
  MXI4X1 U1325 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n567), .S1(n531), .Y(n326) );
  MXI4X1 U1326 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n567), .S1(n531), .Y(n325) );
  MXI2X1 U1327 ( .A(n387), .B(n388), .S0(n508), .Y(blockdata[36]) );
  MXI4X1 U1328 ( .A(\block[4][36] ), .B(\block[5][36] ), .C(\block[6][36] ), 
        .D(\block[7][36] ), .S0(n572), .S1(n536), .Y(n388) );
  MXI4X1 U1329 ( .A(\block[0][36] ), .B(\block[1][36] ), .C(\block[2][36] ), 
        .D(\block[3][36] ), .S0(n572), .S1(n536), .Y(n387) );
  MXI2X1 U1330 ( .A(n323), .B(n324), .S0(n506), .Y(blockdata[68]) );
  MXI4X1 U1331 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n567), .S1(n531), .Y(n324) );
  MXI4X1 U1332 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n567), .S1(n531), .Y(n323) );
  MXI2X1 U1333 ( .A(n385), .B(n386), .S0(n508), .Y(blockdata[37]) );
  MXI4X1 U1334 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n572), .S1(n536), .Y(n386) );
  MXI4X1 U1335 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n572), .S1(n536), .Y(n385) );
  MXI2X1 U1336 ( .A(n321), .B(n322), .S0(n505), .Y(blockdata[69]) );
  MXI4X1 U1337 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), 
        .D(\block[7][69] ), .S0(n567), .S1(n530), .Y(n322) );
  MXI4X1 U1338 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), 
        .D(\block[3][69] ), .S0(n567), .S1(n530), .Y(n321) );
  MXI2X1 U1339 ( .A(n383), .B(n384), .S0(n508), .Y(blockdata[38]) );
  MXI4X1 U1340 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), 
        .D(\block[7][38] ), .S0(n571), .S1(n536), .Y(n384) );
  MXI4X1 U1341 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), 
        .D(\block[3][38] ), .S0(n571), .S1(n536), .Y(n383) );
  MXI2X1 U1342 ( .A(n319), .B(n320), .S0(n505), .Y(blockdata[70]) );
  MXI4X1 U1343 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), 
        .D(\block[7][70] ), .S0(n566), .S1(n530), .Y(n320) );
  MXI4X1 U1344 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), 
        .D(\block[3][70] ), .S0(n567), .S1(n530), .Y(n319) );
  MXI2X1 U1345 ( .A(n381), .B(n382), .S0(n508), .Y(blockdata[39]) );
  MXI4X1 U1346 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), 
        .D(\block[7][39] ), .S0(n571), .S1(n535), .Y(n382) );
  MXI4X1 U1347 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), 
        .D(\block[3][39] ), .S0(n571), .S1(n535), .Y(n381) );
  MXI2X1 U1348 ( .A(n317), .B(n318), .S0(n505), .Y(blockdata[71]) );
  MXI4X1 U1349 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), 
        .D(\block[7][71] ), .S0(n566), .S1(n530), .Y(n318) );
  MXI4X1 U1350 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), 
        .D(\block[3][71] ), .S0(n566), .S1(n530), .Y(n317) );
  MXI2X1 U1351 ( .A(n379), .B(n380), .S0(n508), .Y(blockdata[40]) );
  MXI4X1 U1352 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), 
        .D(\block[7][40] ), .S0(n571), .S1(n535), .Y(n380) );
  MXI4X1 U1353 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n571), .S1(n535), .Y(n379) );
  MXI2X1 U1354 ( .A(n315), .B(n316), .S0(n505), .Y(blockdata[72]) );
  MXI4X1 U1355 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), 
        .D(\block[7][72] ), .S0(n566), .S1(n530), .Y(n316) );
  MXI4X1 U1356 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n566), .S1(n530), .Y(n315) );
  MXI2X1 U1357 ( .A(n377), .B(n378), .S0(n508), .Y(blockdata[41]) );
  MXI4X1 U1358 ( .A(\block[4][41] ), .B(\block[5][41] ), .C(\block[6][41] ), 
        .D(\block[7][41] ), .S0(n571), .S1(n535), .Y(n378) );
  MXI4X1 U1359 ( .A(\block[0][41] ), .B(\block[1][41] ), .C(\block[2][41] ), 
        .D(\block[3][41] ), .S0(n571), .S1(n535), .Y(n377) );
  MXI2X1 U1360 ( .A(n313), .B(n314), .S0(n505), .Y(blockdata[73]) );
  MXI4X1 U1361 ( .A(\block[4][73] ), .B(\block[5][73] ), .C(\block[6][73] ), 
        .D(\block[7][73] ), .S0(n566), .S1(n530), .Y(n314) );
  MXI4X1 U1362 ( .A(\block[0][73] ), .B(\block[1][73] ), .C(\block[2][73] ), 
        .D(\block[3][73] ), .S0(n566), .S1(n530), .Y(n313) );
  MXI2X1 U1363 ( .A(n375), .B(n376), .S0(n508), .Y(blockdata[42]) );
  MXI4X1 U1364 ( .A(\block[4][42] ), .B(\block[5][42] ), .C(\block[6][42] ), 
        .D(\block[7][42] ), .S0(n571), .S1(n535), .Y(n376) );
  MXI4X1 U1365 ( .A(\block[0][42] ), .B(\block[1][42] ), .C(\block[2][42] ), 
        .D(\block[3][42] ), .S0(n571), .S1(n535), .Y(n375) );
  MXI2X1 U1366 ( .A(n311), .B(n312), .S0(n505), .Y(blockdata[74]) );
  MXI4X1 U1367 ( .A(\block[4][74] ), .B(\block[5][74] ), .C(\block[6][74] ), 
        .D(\block[7][74] ), .S0(n566), .S1(n530), .Y(n312) );
  MXI4X1 U1368 ( .A(\block[0][74] ), .B(\block[1][74] ), .C(\block[2][74] ), 
        .D(\block[3][74] ), .S0(n566), .S1(n530), .Y(n311) );
  MXI2X1 U1369 ( .A(n373), .B(n374), .S0(n508), .Y(blockdata[43]) );
  MXI4X1 U1370 ( .A(\block[4][43] ), .B(\block[5][43] ), .C(\block[6][43] ), 
        .D(\block[7][43] ), .S0(n571), .S1(n535), .Y(n374) );
  MXI4X1 U1371 ( .A(\block[0][43] ), .B(\block[1][43] ), .C(\block[2][43] ), 
        .D(\block[3][43] ), .S0(n571), .S1(n535), .Y(n373) );
  MXI2X1 U1372 ( .A(n309), .B(n310), .S0(n505), .Y(blockdata[75]) );
  MXI4X1 U1373 ( .A(\block[4][75] ), .B(\block[5][75] ), .C(\block[6][75] ), 
        .D(\block[7][75] ), .S0(n566), .S1(n529), .Y(n310) );
  MXI4X1 U1374 ( .A(\block[0][75] ), .B(\block[1][75] ), .C(\block[2][75] ), 
        .D(\block[3][75] ), .S0(n566), .S1(n529), .Y(n309) );
  MXI2X1 U1375 ( .A(n371), .B(n372), .S0(n508), .Y(blockdata[44]) );
  MXI4X1 U1376 ( .A(\block[4][44] ), .B(\block[5][44] ), .C(\block[6][44] ), 
        .D(\block[7][44] ), .S0(n570), .S1(n535), .Y(n372) );
  MXI4X1 U1377 ( .A(\block[0][44] ), .B(\block[1][44] ), .C(\block[2][44] ), 
        .D(\block[3][44] ), .S0(n571), .S1(n535), .Y(n371) );
  MXI2X1 U1378 ( .A(n307), .B(n308), .S0(n505), .Y(blockdata[76]) );
  MXI4X1 U1379 ( .A(\block[4][76] ), .B(\block[5][76] ), .C(\block[6][76] ), 
        .D(\block[7][76] ), .S0(n566), .S1(n529), .Y(n308) );
  MXI4X1 U1380 ( .A(\block[0][76] ), .B(\block[1][76] ), .C(\block[2][76] ), 
        .D(\block[3][76] ), .S0(n566), .S1(n529), .Y(n307) );
  MXI2X1 U1381 ( .A(n369), .B(n370), .S0(n507), .Y(blockdata[45]) );
  MXI4X1 U1382 ( .A(\block[4][45] ), .B(\block[5][45] ), .C(\block[6][45] ), 
        .D(\block[7][45] ), .S0(n570), .S1(n534), .Y(n370) );
  MXI4X1 U1383 ( .A(\block[0][45] ), .B(\block[1][45] ), .C(\block[2][45] ), 
        .D(\block[3][45] ), .S0(n570), .S1(n534), .Y(n369) );
  MXI2X1 U1384 ( .A(n305), .B(n306), .S0(n505), .Y(blockdata[77]) );
  MXI4X1 U1385 ( .A(\block[4][77] ), .B(\block[5][77] ), .C(\block[6][77] ), 
        .D(\block[7][77] ), .S0(n565), .S1(n529), .Y(n306) );
  MXI4X1 U1386 ( .A(\block[0][77] ), .B(\block[1][77] ), .C(\block[2][77] ), 
        .D(\block[3][77] ), .S0(n565), .S1(n529), .Y(n305) );
  MXI2X1 U1387 ( .A(n367), .B(n368), .S0(n507), .Y(blockdata[46]) );
  MXI4X1 U1388 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), 
        .D(\block[7][46] ), .S0(n570), .S1(n534), .Y(n368) );
  MXI4X1 U1389 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n570), .S1(n534), .Y(n367) );
  MXI2X1 U1390 ( .A(n303), .B(n304), .S0(n505), .Y(blockdata[78]) );
  MXI4X1 U1391 ( .A(\block[4][78] ), .B(\block[5][78] ), .C(\block[6][78] ), 
        .D(\block[7][78] ), .S0(n565), .S1(n529), .Y(n304) );
  MXI4X1 U1392 ( .A(\block[0][78] ), .B(\block[1][78] ), .C(\block[2][78] ), 
        .D(\block[3][78] ), .S0(n565), .S1(n529), .Y(n303) );
  MXI2X1 U1393 ( .A(n365), .B(n366), .S0(n507), .Y(blockdata[47]) );
  MXI4X1 U1394 ( .A(\block[4][47] ), .B(\block[5][47] ), .C(\block[6][47] ), 
        .D(\block[7][47] ), .S0(n570), .S1(n534), .Y(n366) );
  MXI4X1 U1395 ( .A(\block[0][47] ), .B(\block[1][47] ), .C(\block[2][47] ), 
        .D(\block[3][47] ), .S0(n570), .S1(n534), .Y(n365) );
  MXI2X1 U1396 ( .A(n301), .B(n302), .S0(n505), .Y(blockdata[79]) );
  MXI4X1 U1397 ( .A(\block[4][79] ), .B(\block[5][79] ), .C(\block[6][79] ), 
        .D(\block[7][79] ), .S0(n565), .S1(n529), .Y(n302) );
  MXI4X1 U1398 ( .A(\block[0][79] ), .B(\block[1][79] ), .C(\block[2][79] ), 
        .D(\block[3][79] ), .S0(n565), .S1(n529), .Y(n301) );
  MXI2X1 U1399 ( .A(n363), .B(n364), .S0(n507), .Y(blockdata[48]) );
  MXI4X1 U1400 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n570), .S1(n534), .Y(n364) );
  MXI4X1 U1401 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n570), .S1(n534), .Y(n363) );
  MXI2X1 U1402 ( .A(n299), .B(n300), .S0(n505), .Y(blockdata[80]) );
  MXI4X1 U1403 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n565), .S1(n529), .Y(n300) );
  MXI4X1 U1404 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n565), .S1(n529), .Y(n299) );
  MXI2X1 U1405 ( .A(n361), .B(n362), .S0(n507), .Y(blockdata[49]) );
  MXI4X1 U1406 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n570), .S1(n534), .Y(n362) );
  MXI4X1 U1407 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n570), .S1(n534), .Y(n361) );
  MXI2X1 U1408 ( .A(n297), .B(n298), .S0(n504), .Y(blockdata[81]) );
  MXI4X1 U1409 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n565), .S1(n528), .Y(n298) );
  MXI4X1 U1410 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n565), .S1(n523), .Y(n297) );
  MXI2X1 U1411 ( .A(n359), .B(n360), .S0(n507), .Y(blockdata[50]) );
  MXI4X1 U1412 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n570), .S1(n534), .Y(n360) );
  MXI4X1 U1413 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n570), .S1(n534), .Y(n359) );
  MXI2X1 U1414 ( .A(n295), .B(n296), .S0(n504), .Y(blockdata[82]) );
  MXI4X1 U1415 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n565), .S1(n523), .Y(n296) );
  MXI4X1 U1416 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n565), .S1(n525), .Y(n295) );
  MXI2X1 U1417 ( .A(n357), .B(n358), .S0(n507), .Y(blockdata[51]) );
  MXI4X1 U1418 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n569), .S1(n533), .Y(n358) );
  MXI4X1 U1419 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n569), .S1(n533), .Y(n357) );
  MXI2X1 U1420 ( .A(n293), .B(n294), .S0(n504), .Y(blockdata[83]) );
  MXI4X1 U1421 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n564), .S1(n530), .Y(n294) );
  MXI4X1 U1422 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n565), .S1(n529), .Y(n293) );
  MXI2X1 U1423 ( .A(n355), .B(n356), .S0(n507), .Y(blockdata[52]) );
  MXI4X1 U1424 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n569), .S1(n533), .Y(n356) );
  MXI4X1 U1425 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n569), .S1(n533), .Y(n355) );
  MXI2X1 U1426 ( .A(n291), .B(n292), .S0(n504), .Y(blockdata[84]) );
  MXI4X1 U1427 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n564), .S1(n529), .Y(n292) );
  MXI4X1 U1428 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n564), .S1(n522), .Y(n291) );
  MXI2X1 U1429 ( .A(n353), .B(n354), .S0(n507), .Y(blockdata[53]) );
  MXI4X1 U1430 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n569), .S1(n533), .Y(n354) );
  MXI4X1 U1431 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n569), .S1(n533), .Y(n353) );
  MXI2X1 U1432 ( .A(n289), .B(n290), .S0(n504), .Y(blockdata[85]) );
  MXI4X1 U1433 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n564), .S1(n530), .Y(n290) );
  MXI4X1 U1434 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n564), .S1(n523), .Y(n289) );
  MXI2X1 U1435 ( .A(n351), .B(n352), .S0(n507), .Y(blockdata[54]) );
  MXI4X1 U1436 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n569), .S1(n533), .Y(n352) );
  MXI4X1 U1437 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n569), .S1(n533), .Y(n351) );
  MXI2X1 U1438 ( .A(n287), .B(n288), .S0(n504), .Y(blockdata[86]) );
  MXI4X1 U1439 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n564), .S1(n528), .Y(n288) );
  MXI4X1 U1440 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n564), .S1(n526), .Y(n287) );
  MXI2X1 U1441 ( .A(n349), .B(n350), .S0(n507), .Y(blockdata[55]) );
  MXI4X1 U1442 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n569), .S1(n533), .Y(n350) );
  MXI4X1 U1443 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n569), .S1(n533), .Y(n349) );
  MXI2X1 U1444 ( .A(n285), .B(n286), .S0(n504), .Y(blockdata[87]) );
  MXI4X1 U1445 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n564), .S1(n528), .Y(n286) );
  MXI4X1 U1446 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n564), .S1(n528), .Y(n285) );
  MXI2X1 U1447 ( .A(n347), .B(n348), .S0(n507), .Y(blockdata[56]) );
  MXI4X1 U1448 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n569), .S1(n533), .Y(n348) );
  MXI4X1 U1449 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n569), .S1(n533), .Y(n347) );
  MXI2X1 U1450 ( .A(n283), .B(n284), .S0(n504), .Y(blockdata[88]) );
  MXI4X1 U1451 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n564), .S1(n528), .Y(n284) );
  MXI4X1 U1452 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n564), .S1(n528), .Y(n283) );
  MXI2X1 U1453 ( .A(n345), .B(n346), .S0(n506), .Y(blockdata[57]) );
  MXI4X1 U1454 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n568), .S1(n532), .Y(n346) );
  MXI4X1 U1455 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n569), .S1(n532), .Y(n345) );
  MXI2X1 U1456 ( .A(n281), .B(n282), .S0(n504), .Y(blockdata[89]) );
  MXI4X1 U1457 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n564), .S1(n528), .Y(n282) );
  MXI4X1 U1458 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n564), .S1(n528), .Y(n281) );
  MXI2X1 U1459 ( .A(n343), .B(n344), .S0(n506), .Y(blockdata[58]) );
  MXI4X1 U1460 ( .A(\block[4][58] ), .B(\block[5][58] ), .C(\block[6][58] ), 
        .D(\block[7][58] ), .S0(n568), .S1(n532), .Y(n344) );
  MXI4X1 U1461 ( .A(\block[0][58] ), .B(\block[1][58] ), .C(\block[2][58] ), 
        .D(\block[3][58] ), .S0(n568), .S1(n532), .Y(n343) );
  MXI2X1 U1462 ( .A(n279), .B(n280), .S0(n504), .Y(blockdata[90]) );
  MXI4X1 U1463 ( .A(\block[4][90] ), .B(\block[5][90] ), .C(\block[6][90] ), 
        .D(\block[7][90] ), .S0(n563), .S1(n528), .Y(n280) );
  MXI4X1 U1464 ( .A(\block[0][90] ), .B(\block[1][90] ), .C(\block[2][90] ), 
        .D(\block[3][90] ), .S0(n563), .S1(n528), .Y(n279) );
  MXI2X1 U1465 ( .A(n341), .B(n342), .S0(n506), .Y(blockdata[59]) );
  MXI4X1 U1466 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), 
        .D(\block[7][59] ), .S0(n568), .S1(n532), .Y(n342) );
  MXI4X1 U1467 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), 
        .D(\block[3][59] ), .S0(n568), .S1(n532), .Y(n341) );
  MXI2X1 U1468 ( .A(n277), .B(n278), .S0(n504), .Y(blockdata[91]) );
  MXI4X1 U1469 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), 
        .D(\block[7][91] ), .S0(n563), .S1(n528), .Y(n278) );
  MXI4X1 U1470 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), 
        .D(\block[3][91] ), .S0(n563), .S1(n528), .Y(n277) );
  MXI2X1 U1471 ( .A(n339), .B(n340), .S0(n506), .Y(blockdata[60]) );
  MXI4X1 U1472 ( .A(\block[4][60] ), .B(\block[5][60] ), .C(\block[6][60] ), 
        .D(\block[7][60] ), .S0(n568), .S1(n532), .Y(n340) );
  MXI4X1 U1473 ( .A(\block[0][60] ), .B(\block[1][60] ), .C(\block[2][60] ), 
        .D(\block[3][60] ), .S0(n568), .S1(n532), .Y(n339) );
  MXI2X1 U1474 ( .A(n275), .B(n276), .S0(n504), .Y(blockdata[92]) );
  MXI4X1 U1475 ( .A(\block[4][92] ), .B(\block[5][92] ), .C(\block[6][92] ), 
        .D(\block[7][92] ), .S0(n563), .S1(n528), .Y(n276) );
  MXI4X1 U1476 ( .A(\block[0][92] ), .B(\block[1][92] ), .C(\block[2][92] ), 
        .D(\block[3][92] ), .S0(n563), .S1(n528), .Y(n275) );
  MXI2X1 U1477 ( .A(n337), .B(n338), .S0(n506), .Y(blockdata[61]) );
  MXI4X1 U1478 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n568), .S1(n532), .Y(n338) );
  MXI4X1 U1479 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n568), .S1(n532), .Y(n337) );
  MXI2X1 U1480 ( .A(n273), .B(n274), .S0(n502), .Y(blockdata[93]) );
  MXI4X1 U1481 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n563), .S1(n527), .Y(n274) );
  MXI4X1 U1482 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n563), .S1(n527), .Y(n273) );
  MXI2X1 U1483 ( .A(n335), .B(n336), .S0(n506), .Y(blockdata[62]) );
  MXI4X1 U1484 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n568), .S1(n532), .Y(n336) );
  MXI4X1 U1485 ( .A(\block[0][62] ), .B(\block[1][62] ), .C(\block[2][62] ), 
        .D(\block[3][62] ), .S0(n568), .S1(n532), .Y(n335) );
  MXI2X1 U1486 ( .A(n271), .B(n272), .S0(n502), .Y(blockdata[94]) );
  MXI4X1 U1487 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), 
        .D(\block[7][94] ), .S0(n563), .S1(n527), .Y(n272) );
  MXI4X1 U1488 ( .A(\block[0][94] ), .B(\block[1][94] ), .C(\block[2][94] ), 
        .D(\block[3][94] ), .S0(n563), .S1(n527), .Y(n271) );
  MXI2X1 U1489 ( .A(n333), .B(n334), .S0(n506), .Y(blockdata[63]) );
  MXI4X1 U1490 ( .A(\block[4][63] ), .B(\block[5][63] ), .C(\block[6][63] ), 
        .D(\block[7][63] ), .S0(n568), .S1(n531), .Y(n334) );
  MXI4X1 U1491 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n568), .S1(n531), .Y(n333) );
  MXI2X1 U1492 ( .A(n269), .B(n270), .S0(n502), .Y(blockdata[95]) );
  MXI4X1 U1493 ( .A(\block[4][95] ), .B(\block[5][95] ), .C(\block[6][95] ), 
        .D(\block[7][95] ), .S0(n563), .S1(n527), .Y(n270) );
  MXI4X1 U1494 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n563), .S1(n527), .Y(n269) );
  MXI2X1 U1495 ( .A(n267), .B(n268), .S0(n502), .Y(blockdata[96]) );
  MXI4X1 U1496 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n562), .S1(n527), .Y(n268) );
  MXI4X1 U1497 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n563), .S1(n527), .Y(n267) );
  MXI2X1 U1498 ( .A(n265), .B(n266), .S0(n502), .Y(blockdata[97]) );
  MXI4X1 U1499 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n562), .S1(n527), .Y(n266) );
  MXI4X1 U1500 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n562), .S1(n527), .Y(n265) );
  MXI2X1 U1501 ( .A(n263), .B(n264), .S0(n502), .Y(blockdata[98]) );
  MXI4X1 U1502 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n562), .S1(n527), .Y(n264) );
  MXI4X1 U1503 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n562), .S1(n527), .Y(n263) );
  MXI2X1 U1504 ( .A(n261), .B(n262), .S0(n502), .Y(blockdata[99]) );
  MXI4X1 U1505 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), 
        .D(\block[7][99] ), .S0(n562), .S1(n526), .Y(n262) );
  MXI4X1 U1506 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), 
        .D(\block[3][99] ), .S0(n562), .S1(n526), .Y(n261) );
  MXI2X1 U1507 ( .A(n259), .B(n260), .S0(n502), .Y(blockdata[100]) );
  MXI4X1 U1508 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n562), .S1(n526), .Y(n260) );
  MXI4X1 U1509 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n562), .S1(n526), .Y(n259) );
  MXI2X1 U1510 ( .A(n257), .B(n258), .S0(n502), .Y(blockdata[101]) );
  MXI4X1 U1511 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n562), .S1(n526), .Y(n258) );
  MXI4X1 U1512 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n562), .S1(n526), .Y(n257) );
  MXI2X1 U1513 ( .A(n255), .B(n256), .S0(n502), .Y(blockdata[102]) );
  MXI4X1 U1514 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n562), .S1(n526), .Y(n256) );
  MXI4X1 U1515 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n562), .S1(n526), .Y(n255) );
  MXI2X1 U1516 ( .A(n253), .B(n254), .S0(n502), .Y(blockdata[103]) );
  MXI4X1 U1517 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n561), .S1(n526), .Y(n254) );
  MXI4X1 U1518 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n561), .S1(n526), .Y(n253) );
  MXI2X1 U1519 ( .A(n251), .B(n252), .S0(n502), .Y(blockdata[104]) );
  MXI4X1 U1520 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n561), .S1(n526), .Y(n252) );
  MXI4X1 U1521 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n561), .S1(n526), .Y(n251) );
  MXI2X1 U1522 ( .A(n249), .B(n250), .S0(n470), .Y(blockdata[105]) );
  MXI4X1 U1523 ( .A(\block[4][105] ), .B(\block[5][105] ), .C(\block[6][105] ), 
        .D(\block[7][105] ), .S0(n561), .S1(n525), .Y(n250) );
  MXI4X1 U1524 ( .A(\block[0][105] ), .B(\block[1][105] ), .C(\block[2][105] ), 
        .D(\block[3][105] ), .S0(n561), .S1(n525), .Y(n249) );
  MXI2X1 U1525 ( .A(n247), .B(n248), .S0(n470), .Y(blockdata[106]) );
  MXI4X1 U1526 ( .A(\block[4][106] ), .B(\block[5][106] ), .C(\block[6][106] ), 
        .D(\block[7][106] ), .S0(n561), .S1(n525), .Y(n248) );
  MXI4X1 U1527 ( .A(\block[0][106] ), .B(\block[1][106] ), .C(\block[2][106] ), 
        .D(\block[3][106] ), .S0(n561), .S1(n525), .Y(n247) );
  MXI2X1 U1528 ( .A(n245), .B(n246), .S0(n470), .Y(blockdata[107]) );
  MXI4X1 U1529 ( .A(\block[4][107] ), .B(\block[5][107] ), .C(\block[6][107] ), 
        .D(\block[7][107] ), .S0(n561), .S1(n525), .Y(n246) );
  MXI4X1 U1530 ( .A(\block[0][107] ), .B(\block[1][107] ), .C(\block[2][107] ), 
        .D(\block[3][107] ), .S0(n561), .S1(n525), .Y(n245) );
  MXI2X1 U1531 ( .A(n243), .B(n244), .S0(n470), .Y(blockdata[108]) );
  MXI4X1 U1532 ( .A(\block[4][108] ), .B(\block[5][108] ), .C(\block[6][108] ), 
        .D(\block[7][108] ), .S0(n561), .S1(n525), .Y(n244) );
  MXI4X1 U1533 ( .A(\block[0][108] ), .B(\block[1][108] ), .C(\block[2][108] ), 
        .D(\block[3][108] ), .S0(n561), .S1(n525), .Y(n243) );
  MXI2X1 U1534 ( .A(n241), .B(n242), .S0(n470), .Y(blockdata[109]) );
  MXI4X1 U1535 ( .A(\block[4][109] ), .B(\block[5][109] ), .C(\block[6][109] ), 
        .D(\block[7][109] ), .S0(n560), .S1(n525), .Y(n242) );
  MXI4X1 U1536 ( .A(\block[0][109] ), .B(\block[1][109] ), .C(\block[2][109] ), 
        .D(\block[3][109] ), .S0(n561), .S1(n525), .Y(n241) );
  MXI2X1 U1537 ( .A(n239), .B(n240), .S0(n470), .Y(blockdata[110]) );
  MXI4X1 U1538 ( .A(\block[4][110] ), .B(\block[5][110] ), .C(\block[6][110] ), 
        .D(\block[7][110] ), .S0(n560), .S1(n525), .Y(n240) );
  MXI4X1 U1539 ( .A(\block[0][110] ), .B(\block[1][110] ), .C(\block[2][110] ), 
        .D(\block[3][110] ), .S0(n560), .S1(n525), .Y(n239) );
  MXI2X1 U1540 ( .A(n237), .B(n238), .S0(n470), .Y(blockdata[111]) );
  MXI4X1 U1541 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n560), .S1(n524), .Y(n238) );
  MXI4X1 U1542 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n560), .S1(n524), .Y(n237) );
  MXI2X1 U1543 ( .A(n235), .B(n236), .S0(n470), .Y(blockdata[112]) );
  MXI4X1 U1544 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n560), .S1(n524), .Y(n236) );
  MXI4X1 U1545 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n560), .S1(n524), .Y(n235) );
  MXI2X1 U1546 ( .A(n233), .B(n234), .S0(n470), .Y(blockdata[113]) );
  MXI4X1 U1547 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n560), .S1(n524), .Y(n234) );
  MXI4X1 U1548 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n560), .S1(n524), .Y(n233) );
  MXI2X1 U1549 ( .A(n231), .B(n232), .S0(n470), .Y(blockdata[114]) );
  MXI4X1 U1550 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n560), .S1(n524), .Y(n232) );
  MXI4X1 U1551 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n560), .S1(n524), .Y(n231) );
  MXI2X1 U1552 ( .A(n229), .B(n230), .S0(n470), .Y(blockdata[115]) );
  MXI4X1 U1553 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n560), .S1(n524), .Y(n230) );
  MXI4X1 U1554 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n560), .S1(n524), .Y(n229) );
  MXI2X1 U1555 ( .A(n227), .B(n228), .S0(n470), .Y(blockdata[116]) );
  MXI4X1 U1556 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n559), .S1(n524), .Y(n228) );
  MXI4X1 U1557 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n559), .S1(n524), .Y(n227) );
  MXI2X1 U1558 ( .A(n213), .B(n214), .S0(n469), .Y(blockdata[123]) );
  MXI4X1 U1559 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n558), .S1(n522), .Y(n214) );
  MXI4X1 U1560 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n558), .S1(n522), .Y(n213) );
  MXI2X1 U1561 ( .A(n211), .B(n212), .S0(n469), .Y(blockdata[124]) );
  MXI4X1 U1562 ( .A(\block[4][124] ), .B(\block[5][124] ), .C(\block[6][124] ), 
        .D(\block[7][124] ), .S0(n558), .S1(n522), .Y(n212) );
  MXI4X1 U1563 ( .A(\block[0][124] ), .B(\block[1][124] ), .C(\block[2][124] ), 
        .D(\block[3][124] ), .S0(n558), .S1(n522), .Y(n211) );
  MXI2X1 U1564 ( .A(n209), .B(n210), .S0(n469), .Y(blockdata[125]) );
  MXI4X1 U1565 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n558), .S1(n522), .Y(n210) );
  MXI4X1 U1566 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n558), .S1(n522), .Y(n209) );
  MXI2X1 U1567 ( .A(n207), .B(n208), .S0(n469), .Y(blockdata[126]) );
  MXI4X1 U1568 ( .A(\block[4][126] ), .B(\block[5][126] ), .C(\block[6][126] ), 
        .D(\block[7][126] ), .S0(n558), .S1(n522), .Y(n208) );
  MXI4X1 U1569 ( .A(\block[0][126] ), .B(\block[1][126] ), .C(\block[2][126] ), 
        .D(\block[3][126] ), .S0(n558), .S1(n522), .Y(n207) );
  MXI2X1 U1570 ( .A(n205), .B(n206), .S0(n469), .Y(blockdata[127]) );
  MXI4X1 U1571 ( .A(\block[4][127] ), .B(\block[5][127] ), .C(\block[6][127] ), 
        .D(\block[7][127] ), .S0(n558), .S1(n522), .Y(n206) );
  MXI4X1 U1572 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n558), .S1(n522), .Y(n205) );
  OAI221XL U1573 ( .A0(n635), .A1(n1232), .B0(n634), .B1(n1231), .C0(n1230), 
        .Y(proc_rdata[26]) );
  OAI221XL U1574 ( .A0(n635), .A1(n1247), .B0(n634), .B1(n1246), .C0(n1245), 
        .Y(proc_rdata[29]) );
  OA22XL U1575 ( .A0(n628), .A1(n1099), .B0(n624), .B1(n1098), .Y(n1100) );
  OA22XL U1576 ( .A0(n628), .A1(n1109), .B0(n624), .B1(n1108), .Y(n1110) );
  OA22XL U1577 ( .A0(n628), .A1(n1114), .B0(n624), .B1(n1113), .Y(n1115) );
  OA22XL U1578 ( .A0(n629), .A1(n1159), .B0(n625), .B1(n1158), .Y(n1160) );
  OA22XL U1579 ( .A0(n629), .A1(n1164), .B0(n625), .B1(n1163), .Y(n1165) );
  OA22XL U1580 ( .A0(n629), .A1(n1214), .B0(n625), .B1(n1213), .Y(n1215) );
  OAI221XL U1581 ( .A0(n635), .A1(n1227), .B0(n634), .B1(n1226), .C0(n1225), 
        .Y(proc_rdata[25]) );
  INVX1 U1582 ( .A(proc_wdata[22]), .Y(n956) );
  INVX1 U1583 ( .A(proc_wdata[23]), .Y(n954) );
  INVX1 U1584 ( .A(proc_wdata[13]), .Y(n974) );
  INVX1 U1585 ( .A(proc_wdata[14]), .Y(n972) );
  INVX1 U1586 ( .A(proc_wdata[15]), .Y(n970) );
  INVX1 U1587 ( .A(proc_wdata[17]), .Y(n966) );
  INVX1 U1588 ( .A(proc_wdata[18]), .Y(n964) );
  INVX1 U1589 ( .A(proc_wdata[19]), .Y(n962) );
  INVX1 U1590 ( .A(proc_wdata[20]), .Y(n960) );
  INVX1 U1591 ( .A(proc_wdata[21]), .Y(n958) );
  INVX1 U1592 ( .A(proc_wdata[8]), .Y(n984) );
  INVX1 U1593 ( .A(proc_wdata[9]), .Y(n982) );
  INVX1 U1594 ( .A(proc_wdata[10]), .Y(n980) );
  INVX1 U1595 ( .A(proc_wdata[11]), .Y(n978) );
  INVX1 U1596 ( .A(proc_wdata[12]), .Y(n976) );
  INVX1 U1597 ( .A(proc_wdata[0]), .Y(n1000) );
  INVX1 U1598 ( .A(proc_wdata[24]), .Y(n952) );
  INVX1 U1599 ( .A(proc_wdata[1]), .Y(n998) );
  INVX1 U1600 ( .A(proc_wdata[2]), .Y(n996) );
  INVX1 U1601 ( .A(proc_wdata[3]), .Y(n994) );
  INVX1 U1602 ( .A(proc_wdata[4]), .Y(n992) );
  INVX1 U1603 ( .A(proc_wdata[5]), .Y(n990) );
  INVX1 U1604 ( .A(proc_wdata[6]), .Y(n988) );
  INVX1 U1605 ( .A(proc_wdata[7]), .Y(n986) );
  INVX1 U1606 ( .A(proc_wdata[27]), .Y(n946) );
  INVX1 U1607 ( .A(proc_wdata[28]), .Y(n944) );
  INVX1 U1608 ( .A(proc_wdata[29]), .Y(n942) );
  INVX1 U1609 ( .A(proc_wdata[30]), .Y(n940) );
  INVX1 U1610 ( .A(proc_wdata[31]), .Y(n938) );
  INVX1 U1611 ( .A(proc_wdata[26]), .Y(n948) );
  INVX1 U1612 ( .A(proc_wdata[25]), .Y(n950) );
  MXI2X1 U1613 ( .A(n479), .B(n1084), .S0(n1006), .Y(n495) );
  INVXL U1614 ( .A(proc_addr[20]), .Y(n1034) );
  INVXL U1615 ( .A(proc_addr[8]), .Y(n1061) );
  INVX1 U1616 ( .A(proc_addr[27]), .Y(n1013) );
  INVXL U1617 ( .A(proc_addr[6]), .Y(n1067) );
  INVXL U1618 ( .A(proc_addr[12]), .Y(n1056) );
  AO22XL U1619 ( .A0(proc_addr[12]), .A1(mem_read), .B0(tag[7]), .B1(mem_write), .Y(mem_addr[10]) );
  AO22XL U1620 ( .A0(proc_addr[6]), .A1(mem_read), .B0(tag[1]), .B1(mem_write), 
        .Y(mem_addr[4]) );
  AO22X1 U1621 ( .A0(proc_addr[7]), .A1(mem_read), .B0(tag[2]), .B1(mem_write), 
        .Y(mem_addr[5]) );
  AO22X1 U1622 ( .A0(proc_addr[9]), .A1(mem_read), .B0(tag[4]), .B1(mem_write), 
        .Y(mem_addr[7]) );
  AO22X1 U1623 ( .A0(proc_addr[14]), .A1(mem_read), .B0(tag[9]), .B1(mem_write), .Y(mem_addr[12]) );
  INVXL U1624 ( .A(proc_addr[7]), .Y(n1064) );
  NAND3BXL U1625 ( .AN(n1097), .B(proc_addr[1]), .C(n1095), .Y(n1256) );
  CLKINVX3 U1626 ( .A(proc_read), .Y(n831) );
  NAND2X2 U1627 ( .A(n831), .B(n1093), .Y(n1087) );
  CLKINVX3 U1628 ( .A(proc_addr[0]), .Y(n1095) );
  NAND3BX2 U1629 ( .AN(n1096), .B(n832), .C(n1095), .Y(n904) );
  OAI221X2 U1630 ( .A0(n584), .A1(n1206), .B0(n958), .B1(n586), .C0(n846), .Y(
        block_next[117]) );
  OAI221X2 U1631 ( .A0(n585), .A1(n1176), .B0(n970), .B1(n587), .C0(n852), .Y(
        block_next[111]) );
  NAND3BX2 U1632 ( .AN(n601), .B(n151), .C(n608), .Y(n870) );
  OAI221X2 U1633 ( .A0(n590), .A1(n1194), .B0(n962), .B1(n593), .C0(n883), .Y(
        block_next[83]) );
  OAI221X2 U1634 ( .A0(n589), .A1(n1104), .B0(n998), .B1(n592), .C0(n901), .Y(
        block_next[65]) );
  CLKINVX3 U1635 ( .A(n1001), .Y(n1084) );
  CLKINVX3 U1636 ( .A(n1005), .Y(n1085) );
  CLKINVX3 U1637 ( .A(n1009), .Y(blocktag_next[24]) );
  CLKINVX3 U1638 ( .A(n1012), .Y(blocktag_next[23]) );
  CLKINVX3 U1639 ( .A(n1015), .Y(blocktag_next[22]) );
  CLKINVX3 U1640 ( .A(n1018), .Y(blocktag_next[21]) );
  CLKINVX3 U1641 ( .A(n1021), .Y(blocktag_next[20]) );
  CLKINVX3 U1642 ( .A(n1024), .Y(blocktag_next[19]) );
  CLKINVX3 U1643 ( .A(n1027), .Y(blocktag_next[18]) );
  CLKINVX3 U1644 ( .A(n1030), .Y(blocktag_next[17]) );
  CLKINVX3 U1645 ( .A(n1033), .Y(blocktag_next[16]) );
  CLKINVX3 U1646 ( .A(n1036), .Y(blocktag_next[15]) );
  CLKINVX3 U1647 ( .A(n1039), .Y(blocktag_next[14]) );
  CLKINVX3 U1648 ( .A(n1042), .Y(blocktag_next[13]) );
  CLKINVX3 U1649 ( .A(n1045), .Y(blocktag_next[12]) );
  CLKINVX3 U1650 ( .A(n1048), .Y(blocktag_next[11]) );
  CLKINVX3 U1651 ( .A(n1051), .Y(blocktag_next[10]) );
  CLKINVX3 U1652 ( .A(n1055), .Y(blocktag_next[8]) );
  CLKINVX3 U1653 ( .A(n1058), .Y(blocktag_next[7]) );
  CLKINVX3 U1654 ( .A(n1059), .Y(blocktag_next[6]) );
  CLKINVX3 U1655 ( .A(n1063), .Y(blocktag_next[3]) );
  CLKINVX3 U1656 ( .A(n1066), .Y(blocktag_next[2]) );
  CLKINVX3 U1657 ( .A(n1069), .Y(blocktag_next[1]) );
  CLKINVX3 U1658 ( .A(n1073), .Y(blocktag_next[0]) );
  NAND3BX2 U1659 ( .AN(mem_ready), .B(proc_stall), .C(n1089), .Y(n1092) );
  CLKINVX3 U1660 ( .A(n1092), .Y(n1262) );
  AO22X4 U1661 ( .A0(proc_addr[16]), .A1(mem_read), .B0(tag[11]), .B1(
        mem_write), .Y(n1277) );
  AO22X4 U1662 ( .A0(proc_addr[17]), .A1(mem_read), .B0(tag[12]), .B1(
        mem_write), .Y(n1276) );
  AO22X4 U1663 ( .A0(proc_addr[18]), .A1(mem_read), .B0(tag[13]), .B1(
        mem_write), .Y(n1275) );
  AO22X4 U1664 ( .A0(proc_addr[19]), .A1(mem_read), .B0(tag[14]), .B1(
        mem_write), .Y(n1274) );
  AO22X4 U1665 ( .A0(proc_addr[21]), .A1(mem_read), .B0(tag[16]), .B1(
        mem_write), .Y(n1272) );
  AO22X4 U1666 ( .A0(proc_addr[25]), .A1(mem_read), .B0(tag[20]), .B1(
        mem_write), .Y(n1268) );
  AO22X4 U1667 ( .A0(proc_addr[27]), .A1(mem_read), .B0(tag[22]), .B1(
        mem_write), .Y(n1266) );
  AO22X4 U1668 ( .A0(proc_addr[28]), .A1(mem_read), .B0(tag[23]), .B1(
        mem_write), .Y(n1265) );
  NAND3BX2 U1669 ( .AN(proc_addr[0]), .B(n1094), .C(n1096), .Y(n1261) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   N31, N32, N33, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, \blocktag[7][24] , \blocktag[7][23] , \blocktag[7][22] ,
         \blocktag[7][20] , \blocktag[7][19] , \blocktag[7][17] ,
         \blocktag[7][15] , \blocktag[7][14] , \blocktag[7][13] ,
         \blocktag[7][11] , \blocktag[7][10] , \blocktag[7][9] ,
         \blocktag[7][4] , \blocktag[7][2] , \blocktag[7][0] ,
         \blocktag[6][24] , \blocktag[6][23] , \blocktag[6][22] ,
         \blocktag[6][20] , \blocktag[6][19] , \blocktag[6][17] ,
         \blocktag[6][15] , \blocktag[6][14] , \blocktag[6][13] ,
         \blocktag[6][11] , \blocktag[6][10] , \blocktag[6][9] ,
         \blocktag[6][4] , \blocktag[6][2] , \blocktag[6][0] ,
         \blocktag[5][24] , \blocktag[5][23] , \blocktag[5][22] ,
         \blocktag[5][20] , \blocktag[5][19] , \blocktag[5][17] ,
         \blocktag[5][15] , \blocktag[5][14] , \blocktag[5][13] ,
         \blocktag[5][11] , \blocktag[5][10] , \blocktag[5][9] ,
         \blocktag[5][4] , \blocktag[5][2] , \blocktag[5][0] ,
         \blocktag[4][24] , \blocktag[4][23] , \blocktag[4][22] ,
         \blocktag[4][20] , \blocktag[4][19] , \blocktag[4][17] ,
         \blocktag[4][15] , \blocktag[4][14] , \blocktag[4][13] ,
         \blocktag[4][11] , \blocktag[4][10] , \blocktag[4][9] ,
         \blocktag[4][4] , \blocktag[4][2] , \blocktag[4][0] ,
         \blocktag[3][24] , \blocktag[3][23] , \blocktag[3][22] ,
         \blocktag[3][21] , \blocktag[3][19] , \blocktag[3][17] ,
         \blocktag[3][16] , \blocktag[3][15] , \blocktag[3][14] ,
         \blocktag[3][13] , \blocktag[3][11] , \blocktag[3][10] ,
         \blocktag[3][9] , \blocktag[3][4] , \blocktag[3][2] ,
         \blocktag[3][1] , \blocktag[3][0] , \blocktag[2][24] ,
         \blocktag[2][23] , \blocktag[2][22] , \blocktag[2][21] ,
         \blocktag[2][19] , \blocktag[2][17] , \blocktag[2][16] ,
         \blocktag[2][15] , \blocktag[2][14] , \blocktag[2][13] ,
         \blocktag[2][11] , \blocktag[2][10] , \blocktag[2][9] ,
         \blocktag[2][4] , \blocktag[2][2] , \blocktag[2][1] ,
         \blocktag[2][0] , \blocktag[1][24] , \blocktag[1][23] ,
         \blocktag[1][22] , \blocktag[1][21] , \blocktag[1][19] ,
         \blocktag[1][17] , \blocktag[1][16] , \blocktag[1][15] ,
         \blocktag[1][14] , \blocktag[1][13] , \blocktag[1][11] ,
         \blocktag[1][10] , \blocktag[1][9] , \blocktag[1][4] ,
         \blocktag[1][2] , \blocktag[1][1] , \blocktag[1][0] ,
         \blocktag[0][24] , \blocktag[0][23] , \blocktag[0][22] ,
         \blocktag[0][21] , \blocktag[0][19] , \blocktag[0][17] ,
         \blocktag[0][16] , \blocktag[0][15] , \blocktag[0][14] ,
         \blocktag[0][13] , \blocktag[0][11] , \blocktag[0][10] ,
         \blocktag[0][9] , \blocktag[0][4] , \blocktag[0][2] ,
         \blocktag[0][1] , \blocktag[0][0] , valid, dirty, \block[7][125] ,
         \block[7][123] , \block[7][122] , \block[7][121] , \block[7][120] ,
         \block[7][119] , \block[7][118] , \block[7][117] , \block[7][116] ,
         \block[7][115] , \block[7][114] , \block[7][113] , \block[7][112] ,
         \block[7][111] , \block[7][104] , \block[7][103] , \block[7][102] ,
         \block[7][101] , \block[7][100] , \block[7][99] , \block[7][98] ,
         \block[7][97] , \block[7][96] , \block[7][94] , \block[7][93] ,
         \block[7][91] , \block[7][89] , \block[7][88] , \block[7][87] ,
         \block[7][86] , \block[7][85] , \block[7][84] , \block[7][83] ,
         \block[7][82] , \block[7][81] , \block[7][80] , \block[7][72] ,
         \block[7][71] , \block[7][70] , \block[7][69] , \block[7][68] ,
         \block[7][67] , \block[7][66] , \block[7][65] , \block[7][64] ,
         \block[7][62] , \block[7][61] , \block[7][59] , \block[7][57] ,
         \block[7][56] , \block[7][55] , \block[7][54] , \block[7][53] ,
         \block[7][52] , \block[7][51] , \block[7][50] , \block[7][49] ,
         \block[7][48] , \block[7][46] , \block[7][40] , \block[7][39] ,
         \block[7][38] , \block[7][37] , \block[7][35] , \block[7][34] ,
         \block[7][33] , \block[7][32] , \block[7][31] , \block[7][30] ,
         \block[7][29] , \block[7][27] , \block[7][25] , \block[7][24] ,
         \block[7][23] , \block[7][22] , \block[7][21] , \block[7][20] ,
         \block[7][19] , \block[7][18] , \block[7][17] , \block[7][16] ,
         \block[7][15] , \block[7][14] , \block[7][8] , \block[7][7] ,
         \block[7][6] , \block[7][4] , \block[7][3] , \block[7][2] ,
         \block[7][1] , \block[7][0] , \block[6][125] , \block[6][123] ,
         \block[6][122] , \block[6][121] , \block[6][120] , \block[6][119] ,
         \block[6][118] , \block[6][117] , \block[6][116] , \block[6][115] ,
         \block[6][114] , \block[6][113] , \block[6][112] , \block[6][111] ,
         \block[6][104] , \block[6][103] , \block[6][102] , \block[6][101] ,
         \block[6][100] , \block[6][99] , \block[6][98] , \block[6][97] ,
         \block[6][96] , \block[6][94] , \block[6][93] , \block[6][91] ,
         \block[6][89] , \block[6][88] , \block[6][87] , \block[6][86] ,
         \block[6][85] , \block[6][84] , \block[6][83] , \block[6][82] ,
         \block[6][81] , \block[6][80] , \block[6][72] , \block[6][71] ,
         \block[6][70] , \block[6][69] , \block[6][68] , \block[6][67] ,
         \block[6][66] , \block[6][65] , \block[6][64] , \block[6][62] ,
         \block[6][61] , \block[6][59] , \block[6][57] , \block[6][56] ,
         \block[6][55] , \block[6][54] , \block[6][53] , \block[6][52] ,
         \block[6][51] , \block[6][50] , \block[6][49] , \block[6][48] ,
         \block[6][46] , \block[6][40] , \block[6][39] , \block[6][38] ,
         \block[6][37] , \block[6][35] , \block[6][34] , \block[6][33] ,
         \block[6][32] , \block[6][31] , \block[6][30] , \block[6][29] ,
         \block[6][27] , \block[6][25] , \block[6][24] , \block[6][23] ,
         \block[6][22] , \block[6][21] , \block[6][20] , \block[6][19] ,
         \block[6][18] , \block[6][17] , \block[6][16] , \block[6][15] ,
         \block[6][14] , \block[6][8] , \block[6][7] , \block[6][6] ,
         \block[6][4] , \block[6][3] , \block[6][2] , \block[6][1] ,
         \block[6][0] , \block[5][125] , \block[5][123] , \block[5][122] ,
         \block[5][121] , \block[5][120] , \block[5][119] , \block[5][118] ,
         \block[5][117] , \block[5][116] , \block[5][115] , \block[5][114] ,
         \block[5][113] , \block[5][112] , \block[5][111] , \block[5][104] ,
         \block[5][103] , \block[5][102] , \block[5][101] , \block[5][100] ,
         \block[5][99] , \block[5][98] , \block[5][97] , \block[5][96] ,
         \block[5][94] , \block[5][93] , \block[5][91] , \block[5][89] ,
         \block[5][88] , \block[5][87] , \block[5][86] , \block[5][85] ,
         \block[5][84] , \block[5][83] , \block[5][82] , \block[5][81] ,
         \block[5][80] , \block[5][72] , \block[5][71] , \block[5][70] ,
         \block[5][69] , \block[5][68] , \block[5][67] , \block[5][66] ,
         \block[5][65] , \block[5][64] , \block[5][62] , \block[5][61] ,
         \block[5][59] , \block[5][57] , \block[5][56] , \block[5][55] ,
         \block[5][54] , \block[5][53] , \block[5][52] , \block[5][51] ,
         \block[5][50] , \block[5][49] , \block[5][48] , \block[5][46] ,
         \block[5][40] , \block[5][39] , \block[5][38] , \block[5][37] ,
         \block[5][35] , \block[5][34] , \block[5][33] , \block[5][32] ,
         \block[5][31] , \block[5][30] , \block[5][29] , \block[5][27] ,
         \block[5][25] , \block[5][24] , \block[5][23] , \block[5][22] ,
         \block[5][21] , \block[5][20] , \block[5][19] , \block[5][18] ,
         \block[5][17] , \block[5][16] , \block[5][15] , \block[5][14] ,
         \block[5][8] , \block[5][7] , \block[5][6] , \block[5][4] ,
         \block[5][3] , \block[5][2] , \block[5][1] , \block[5][0] ,
         \block[4][125] , \block[4][123] , \block[4][122] , \block[4][121] ,
         \block[4][120] , \block[4][119] , \block[4][118] , \block[4][117] ,
         \block[4][116] , \block[4][115] , \block[4][114] , \block[4][113] ,
         \block[4][112] , \block[4][111] , \block[4][104] , \block[4][103] ,
         \block[4][102] , \block[4][101] , \block[4][100] , \block[4][99] ,
         \block[4][98] , \block[4][97] , \block[4][96] , \block[4][94] ,
         \block[4][93] , \block[4][91] , \block[4][89] , \block[4][88] ,
         \block[4][87] , \block[4][86] , \block[4][85] , \block[4][84] ,
         \block[4][83] , \block[4][82] , \block[4][81] , \block[4][80] ,
         \block[4][72] , \block[4][71] , \block[4][70] , \block[4][69] ,
         \block[4][68] , \block[4][67] , \block[4][66] , \block[4][65] ,
         \block[4][64] , \block[4][62] , \block[4][61] , \block[4][59] ,
         \block[4][57] , \block[4][56] , \block[4][55] , \block[4][54] ,
         \block[4][53] , \block[4][52] , \block[4][51] , \block[4][50] ,
         \block[4][49] , \block[4][48] , \block[4][46] , \block[4][40] ,
         \block[4][39] , \block[4][38] , \block[4][37] , \block[4][35] ,
         \block[4][34] , \block[4][33] , \block[4][32] , \block[4][31] ,
         \block[4][30] , \block[4][29] , \block[4][27] , \block[4][25] ,
         \block[4][24] , \block[4][23] , \block[4][22] , \block[4][21] ,
         \block[4][20] , \block[4][19] , \block[4][18] , \block[4][17] ,
         \block[4][16] , \block[4][15] , \block[4][14] , \block[4][8] ,
         \block[4][7] , \block[4][6] , \block[4][4] , \block[4][3] ,
         \block[4][2] , \block[4][1] , \block[4][0] , \block[3][127] ,
         \block[3][125] , \block[3][123] , \block[3][122] , \block[3][121] ,
         \block[3][120] , \block[3][119] , \block[3][118] , \block[3][117] ,
         \block[3][116] , \block[3][115] , \block[3][114] , \block[3][113] ,
         \block[3][112] , \block[3][111] , \block[3][104] , \block[3][103] ,
         \block[3][102] , \block[3][101] , \block[3][100] , \block[3][99] ,
         \block[3][98] , \block[3][97] , \block[3][96] , \block[3][95] ,
         \block[3][93] , \block[3][91] , \block[3][89] , \block[3][88] ,
         \block[3][87] , \block[3][86] , \block[3][85] , \block[3][84] ,
         \block[3][83] , \block[3][82] , \block[3][81] , \block[3][80] ,
         \block[3][72] , \block[3][71] , \block[3][70] , \block[3][69] ,
         \block[3][68] , \block[3][67] , \block[3][66] , \block[3][65] ,
         \block[3][64] , \block[3][63] , \block[3][61] , \block[3][59] ,
         \block[3][57] , \block[3][56] , \block[3][55] , \block[3][54] ,
         \block[3][53] , \block[3][52] , \block[3][51] , \block[3][50] ,
         \block[3][49] , \block[3][48] , \block[3][46] , \block[3][40] ,
         \block[3][39] , \block[3][38] , \block[3][37] , \block[3][35] ,
         \block[3][34] , \block[3][33] , \block[3][32] , \block[3][30] ,
         \block[3][29] , \block[3][27] , \block[3][25] , \block[3][24] ,
         \block[3][23] , \block[3][22] , \block[3][21] , \block[3][20] ,
         \block[3][19] , \block[3][18] , \block[3][17] , \block[3][16] ,
         \block[3][15] , \block[3][14] , \block[3][8] , \block[3][7] ,
         \block[3][6] , \block[3][4] , \block[3][3] , \block[3][2] ,
         \block[3][1] , \block[3][0] , \block[2][127] , \block[2][125] ,
         \block[2][123] , \block[2][122] , \block[2][121] , \block[2][120] ,
         \block[2][119] , \block[2][118] , \block[2][117] , \block[2][116] ,
         \block[2][115] , \block[2][114] , \block[2][113] , \block[2][112] ,
         \block[2][111] , \block[2][104] , \block[2][103] , \block[2][102] ,
         \block[2][101] , \block[2][100] , \block[2][99] , \block[2][98] ,
         \block[2][97] , \block[2][96] , \block[2][95] , \block[2][93] ,
         \block[2][91] , \block[2][89] , \block[2][88] , \block[2][87] ,
         \block[2][86] , \block[2][85] , \block[2][84] , \block[2][83] ,
         \block[2][82] , \block[2][81] , \block[2][80] , \block[2][72] ,
         \block[2][71] , \block[2][70] , \block[2][69] , \block[2][68] ,
         \block[2][67] , \block[2][66] , \block[2][65] , \block[2][64] ,
         \block[2][63] , \block[2][61] , \block[2][59] , \block[2][57] ,
         \block[2][56] , \block[2][55] , \block[2][54] , \block[2][53] ,
         \block[2][52] , \block[2][51] , \block[2][50] , \block[2][49] ,
         \block[2][48] , \block[2][46] , \block[2][40] , \block[2][39] ,
         \block[2][38] , \block[2][37] , \block[2][35] , \block[2][34] ,
         \block[2][33] , \block[2][32] , \block[2][30] , \block[2][29] ,
         \block[2][27] , \block[2][25] , \block[2][24] , \block[2][23] ,
         \block[2][22] , \block[2][21] , \block[2][20] , \block[2][19] ,
         \block[2][18] , \block[2][17] , \block[2][16] , \block[2][15] ,
         \block[2][14] , \block[2][8] , \block[2][7] , \block[2][6] ,
         \block[2][4] , \block[2][3] , \block[2][2] , \block[2][1] ,
         \block[2][0] , \block[1][127] , \block[1][125] , \block[1][123] ,
         \block[1][122] , \block[1][121] , \block[1][120] , \block[1][119] ,
         \block[1][118] , \block[1][117] , \block[1][116] , \block[1][115] ,
         \block[1][114] , \block[1][113] , \block[1][112] , \block[1][111] ,
         \block[1][104] , \block[1][103] , \block[1][102] , \block[1][101] ,
         \block[1][100] , \block[1][99] , \block[1][98] , \block[1][97] ,
         \block[1][96] , \block[1][95] , \block[1][93] , \block[1][91] ,
         \block[1][89] , \block[1][88] , \block[1][87] , \block[1][86] ,
         \block[1][85] , \block[1][84] , \block[1][83] , \block[1][82] ,
         \block[1][81] , \block[1][80] , \block[1][72] , \block[1][71] ,
         \block[1][70] , \block[1][69] , \block[1][68] , \block[1][67] ,
         \block[1][66] , \block[1][65] , \block[1][64] , \block[1][63] ,
         \block[1][61] , \block[1][59] , \block[1][57] , \block[1][56] ,
         \block[1][55] , \block[1][54] , \block[1][53] , \block[1][52] ,
         \block[1][51] , \block[1][50] , \block[1][49] , \block[1][48] ,
         \block[1][46] , \block[1][40] , \block[1][39] , \block[1][38] ,
         \block[1][37] , \block[1][35] , \block[1][34] , \block[1][33] ,
         \block[1][32] , \block[1][30] , \block[1][29] , \block[1][27] ,
         \block[1][25] , \block[1][24] , \block[1][23] , \block[1][22] ,
         \block[1][21] , \block[1][20] , \block[1][19] , \block[1][18] ,
         \block[1][17] , \block[1][16] , \block[1][15] , \block[1][14] ,
         \block[1][8] , \block[1][7] , \block[1][6] , \block[1][4] ,
         \block[1][3] , \block[1][2] , \block[1][1] , \block[1][0] ,
         \block[0][127] , \block[0][125] , \block[0][123] , \block[0][122] ,
         \block[0][121] , \block[0][120] , \block[0][119] , \block[0][118] ,
         \block[0][117] , \block[0][116] , \block[0][115] , \block[0][114] ,
         \block[0][113] , \block[0][112] , \block[0][111] , \block[0][104] ,
         \block[0][103] , \block[0][102] , \block[0][101] , \block[0][100] ,
         \block[0][99] , \block[0][98] , \block[0][97] , \block[0][96] ,
         \block[0][95] , \block[0][93] , \block[0][91] , \block[0][89] ,
         \block[0][88] , \block[0][87] , \block[0][86] , \block[0][85] ,
         \block[0][84] , \block[0][83] , \block[0][82] , \block[0][81] ,
         \block[0][80] , \block[0][72] , \block[0][71] , \block[0][70] ,
         \block[0][69] , \block[0][68] , \block[0][67] , \block[0][66] ,
         \block[0][65] , \block[0][64] , \block[0][63] , \block[0][61] ,
         \block[0][59] , \block[0][57] , \block[0][56] , \block[0][55] ,
         \block[0][54] , \block[0][53] , \block[0][52] , \block[0][51] ,
         \block[0][50] , \block[0][49] , \block[0][48] , \block[0][46] ,
         \block[0][40] , \block[0][39] , \block[0][38] , \block[0][37] ,
         \block[0][35] , \block[0][34] , \block[0][33] , \block[0][32] ,
         \block[0][30] , \block[0][29] , \block[0][27] , \block[0][25] ,
         \block[0][24] , \block[0][23] , \block[0][22] , \block[0][21] ,
         \block[0][20] , \block[0][19] , \block[0][18] , \block[0][17] ,
         \block[0][16] , \block[0][15] , \block[0][14] , \block[0][8] ,
         \block[0][7] , \block[0][6] , \block[0][4] , \block[0][3] ,
         \block[0][2] , \block[0][1] , \block[0][0] , n1, n2, n3, n4, n5, n7,
         n9, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n33, n35,
         n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63,
         n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91,
         n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, n113, n115,
         n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, n137,
         n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159,
         n161, n163, n165, n167, n169, n171, n173, n175, n177, n179, n181,
         n183, n185, n187, n189, n191, n193, n195, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n502, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1253, n1254,
         n1255, n1256, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751;
  wire   [24:0] tag;
  wire   [7:0] blockvalid;
  wire   [7:0] blockdirty;
  wire   [127:0] blockdata;
  wire   [127:0] block_next;
  wire   [24:0] blocktag_next;
  assign N31 = proc_addr[2];
  assign N32 = proc_addr[3];
  assign N33 = proc_addr[4];

  EDFFX4 \blocktag_reg[2][21]  ( .D(blocktag_next[21]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][21] ) );
  EDFFX4 \blocktag_reg[1][21]  ( .D(blocktag_next[21]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][21] ) );
  EDFFX4 \blocktag_reg[0][21]  ( .D(blocktag_next[21]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][21] ) );
  DFFRX4 \blockvalid_reg[6]  ( .D(n1717), .CK(clk), .RN(n1259), .QN(n1733) );
  DFFRX4 \blockvalid_reg[0]  ( .D(n1723), .CK(clk), .RN(n1258), .Q(
        blockvalid[0]), .QN(n1739) );
  EDFFXL \block_reg[7][116]  ( .D(block_next[116]), .E(n1110), .CK(clk), .Q(
        \block[7][116] ) );
  EDFFXL \block_reg[7][112]  ( .D(block_next[112]), .E(n1110), .CK(clk), .Q(
        \block[7][112] ) );
  EDFFXL \block_reg[7][89]  ( .D(block_next[89]), .E(n1108), .CK(clk), .Q(
        \block[7][89] ) );
  EDFFXL \block_reg[7][88]  ( .D(block_next[88]), .E(n1108), .CK(clk), .Q(
        \block[7][88] ) );
  EDFFXL \block_reg[7][87]  ( .D(block_next[87]), .E(n1108), .CK(clk), .Q(
        \block[7][87] ) );
  EDFFXL \block_reg[7][86]  ( .D(block_next[86]), .E(n1108), .CK(clk), .Q(
        \block[7][86] ) );
  EDFFXL \block_reg[7][85]  ( .D(block_next[85]), .E(n1108), .CK(clk), .Q(
        \block[7][85] ) );
  EDFFXL \block_reg[7][84]  ( .D(block_next[84]), .E(n1108), .CK(clk), .Q(
        \block[7][84] ) );
  EDFFXL \block_reg[7][83]  ( .D(block_next[83]), .E(n1108), .CK(clk), .Q(
        \block[7][83] ) );
  EDFFXL \block_reg[7][82]  ( .D(block_next[82]), .E(n1108), .CK(clk), .Q(
        \block[7][82] ) );
  EDFFXL \block_reg[7][81]  ( .D(block_next[81]), .E(n1108), .CK(clk), .Q(
        \block[7][81] ) );
  EDFFXL \block_reg[7][80]  ( .D(block_next[80]), .E(n1108), .CK(clk), .Q(
        \block[7][80] ) );
  EDFFXL \block_reg[7][57]  ( .D(block_next[57]), .E(n1106), .CK(clk), .Q(
        \block[7][57] ) );
  EDFFXL \block_reg[7][25]  ( .D(block_next[25]), .E(n1103), .CK(clk), .Q(
        \block[7][25] ) );
  EDFFXL \block_reg[7][24]  ( .D(block_next[24]), .E(n1103), .CK(clk), .Q(
        \block[7][24] ) );
  EDFFXL \block_reg[7][23]  ( .D(block_next[23]), .E(n1103), .CK(clk), .Q(
        \block[7][23] ) );
  EDFFXL \block_reg[7][22]  ( .D(block_next[22]), .E(n1103), .CK(clk), .Q(
        \block[7][22] ) );
  EDFFXL \block_reg[7][21]  ( .D(block_next[21]), .E(n1103), .CK(clk), .Q(
        \block[7][21] ) );
  EDFFXL \block_reg[7][18]  ( .D(block_next[18]), .E(n1103), .CK(clk), .Q(
        \block[7][18] ) );
  EDFFXL \block_reg[7][16]  ( .D(block_next[16]), .E(n1103), .CK(clk), .Q(
        \block[7][16] ) );
  EDFFXL \block_reg[7][121]  ( .D(block_next[121]), .E(n1111), .CK(clk), .Q(
        \block[7][121] ) );
  EDFFXL \block_reg[7][120]  ( .D(block_next[120]), .E(n1111), .CK(clk), .Q(
        \block[7][120] ) );
  EDFFXL \block_reg[7][119]  ( .D(block_next[119]), .E(n1111), .CK(clk), .Q(
        \block[7][119] ) );
  EDFFXL \block_reg[7][118]  ( .D(block_next[118]), .E(n1111), .CK(clk), .Q(
        \block[7][118] ) );
  EDFFXL \block_reg[7][117]  ( .D(block_next[117]), .E(n1110), .CK(clk), .Q(
        \block[7][117] ) );
  EDFFXL \block_reg[7][48]  ( .D(block_next[48]), .E(n1105), .CK(clk), .Q(
        \block[7][48] ) );
  EDFFXL \block_reg[7][115]  ( .D(block_next[115]), .E(n1110), .CK(clk), .Q(
        \block[7][115] ) );
  EDFFXL \block_reg[7][114]  ( .D(block_next[114]), .E(n1110), .CK(clk), .Q(
        \block[7][114] ) );
  EDFFXL \block_reg[7][113]  ( .D(block_next[113]), .E(n1110), .CK(clk), .Q(
        \block[7][113] ) );
  EDFFXL \block_reg[7][17]  ( .D(block_next[17]), .E(n1103), .CK(clk), .Q(
        \block[7][17] ) );
  EDFFXL \block_reg[7][20]  ( .D(block_next[20]), .E(n1103), .CK(clk), .Q(
        \block[7][20] ) );
  EDFFXL \block_reg[7][19]  ( .D(block_next[19]), .E(n1103), .CK(clk), .Q(
        \block[7][19] ) );
  EDFFXL \block_reg[7][50]  ( .D(block_next[50]), .E(n1105), .CK(clk), .Q(
        \block[7][50] ) );
  EDFFXL \block_reg[7][49]  ( .D(block_next[49]), .E(n1105), .CK(clk), .Q(
        \block[7][49] ) );
  EDFFXL \block_reg[3][116]  ( .D(block_next[116]), .E(n1183), .CK(clk), .Q(
        \block[3][116] ) );
  EDFFXL \block_reg[3][112]  ( .D(block_next[112]), .E(n1183), .CK(clk), .Q(
        \block[3][112] ) );
  EDFFXL \block_reg[3][89]  ( .D(block_next[89]), .E(n1181), .CK(clk), .Q(
        \block[3][89] ) );
  EDFFXL \block_reg[3][88]  ( .D(block_next[88]), .E(n1181), .CK(clk), .Q(
        \block[3][88] ) );
  EDFFXL \block_reg[3][87]  ( .D(block_next[87]), .E(n1181), .CK(clk), .Q(
        \block[3][87] ) );
  EDFFXL \block_reg[3][86]  ( .D(block_next[86]), .E(n1181), .CK(clk), .Q(
        \block[3][86] ) );
  EDFFXL \block_reg[3][85]  ( .D(block_next[85]), .E(n1181), .CK(clk), .Q(
        \block[3][85] ) );
  EDFFXL \block_reg[3][84]  ( .D(block_next[84]), .E(n1181), .CK(clk), .Q(
        \block[3][84] ) );
  EDFFXL \block_reg[3][83]  ( .D(block_next[83]), .E(n1181), .CK(clk), .Q(
        \block[3][83] ) );
  EDFFXL \block_reg[3][82]  ( .D(block_next[82]), .E(n1181), .CK(clk), .Q(
        \block[3][82] ) );
  EDFFXL \block_reg[3][81]  ( .D(block_next[81]), .E(n1181), .CK(clk), .Q(
        \block[3][81] ) );
  EDFFXL \block_reg[3][80]  ( .D(block_next[80]), .E(n1181), .CK(clk), .Q(
        \block[3][80] ) );
  EDFFXL \block_reg[3][57]  ( .D(block_next[57]), .E(n1179), .CK(clk), .Q(
        \block[3][57] ) );
  EDFFXL \block_reg[3][25]  ( .D(block_next[25]), .E(n1176), .CK(clk), .Q(
        \block[3][25] ) );
  EDFFXL \block_reg[3][24]  ( .D(block_next[24]), .E(n1176), .CK(clk), .Q(
        \block[3][24] ) );
  EDFFXL \block_reg[3][23]  ( .D(block_next[23]), .E(n1176), .CK(clk), .Q(
        \block[3][23] ) );
  EDFFXL \block_reg[3][22]  ( .D(block_next[22]), .E(n1176), .CK(clk), .Q(
        \block[3][22] ) );
  EDFFXL \block_reg[3][21]  ( .D(block_next[21]), .E(n1176), .CK(clk), .Q(
        \block[3][21] ) );
  EDFFXL \block_reg[3][18]  ( .D(block_next[18]), .E(n1176), .CK(clk), .Q(
        \block[3][18] ) );
  EDFFXL \block_reg[3][16]  ( .D(block_next[16]), .E(n1176), .CK(clk), .Q(
        \block[3][16] ) );
  EDFFXL \block_reg[3][121]  ( .D(block_next[121]), .E(n1184), .CK(clk), .Q(
        \block[3][121] ) );
  EDFFXL \block_reg[3][120]  ( .D(block_next[120]), .E(n1184), .CK(clk), .Q(
        \block[3][120] ) );
  EDFFXL \block_reg[3][119]  ( .D(block_next[119]), .E(n1184), .CK(clk), .Q(
        \block[3][119] ) );
  EDFFXL \block_reg[3][118]  ( .D(block_next[118]), .E(n1184), .CK(clk), .Q(
        \block[3][118] ) );
  EDFFXL \block_reg[3][117]  ( .D(block_next[117]), .E(n1183), .CK(clk), .Q(
        \block[3][117] ) );
  EDFFXL \block_reg[7][56]  ( .D(block_next[56]), .E(n1106), .CK(clk), .Q(
        \block[7][56] ) );
  EDFFXL \block_reg[7][55]  ( .D(block_next[55]), .E(n1106), .CK(clk), .Q(
        \block[7][55] ) );
  EDFFXL \block_reg[7][54]  ( .D(block_next[54]), .E(n1106), .CK(clk), .Q(
        \block[7][54] ) );
  EDFFXL \block_reg[7][53]  ( .D(block_next[53]), .E(n1106), .CK(clk), .Q(
        \block[7][53] ) );
  EDFFXL \block_reg[7][52]  ( .D(block_next[52]), .E(n1105), .CK(clk), .Q(
        \block[7][52] ) );
  EDFFXL \block_reg[7][51]  ( .D(block_next[51]), .E(n1105), .CK(clk), .Q(
        \block[7][51] ) );
  EDFFXL \block_reg[3][48]  ( .D(block_next[48]), .E(n1178), .CK(clk), .Q(
        \block[3][48] ) );
  EDFFXL \block_reg[3][115]  ( .D(block_next[115]), .E(n1183), .CK(clk), .Q(
        \block[3][115] ) );
  EDFFXL \block_reg[3][114]  ( .D(block_next[114]), .E(n1183), .CK(clk), .Q(
        \block[3][114] ) );
  EDFFXL \block_reg[3][113]  ( .D(block_next[113]), .E(n1183), .CK(clk), .Q(
        \block[3][113] ) );
  EDFFXL \block_reg[3][17]  ( .D(block_next[17]), .E(n1176), .CK(clk), .Q(
        \block[3][17] ) );
  EDFFXL \block_reg[3][20]  ( .D(block_next[20]), .E(n1176), .CK(clk), .Q(
        \block[3][20] ) );
  EDFFXL \block_reg[3][19]  ( .D(block_next[19]), .E(n1176), .CK(clk), .Q(
        \block[3][19] ) );
  EDFFXL \block_reg[3][50]  ( .D(block_next[50]), .E(n1178), .CK(clk), .Q(
        \block[3][50] ) );
  EDFFXL \block_reg[3][49]  ( .D(block_next[49]), .E(n1178), .CK(clk), .Q(
        \block[3][49] ) );
  EDFFXL \block_reg[3][56]  ( .D(block_next[56]), .E(n1179), .CK(clk), .Q(
        \block[3][56] ) );
  EDFFXL \block_reg[3][55]  ( .D(block_next[55]), .E(n1179), .CK(clk), .Q(
        \block[3][55] ) );
  EDFFXL \block_reg[3][54]  ( .D(block_next[54]), .E(n1179), .CK(clk), .Q(
        \block[3][54] ) );
  EDFFXL \block_reg[3][53]  ( .D(block_next[53]), .E(n1179), .CK(clk), .Q(
        \block[3][53] ) );
  EDFFXL \block_reg[3][52]  ( .D(block_next[52]), .E(n1178), .CK(clk), .Q(
        \block[3][52] ) );
  EDFFXL \block_reg[3][51]  ( .D(block_next[51]), .E(n1178), .CK(clk), .Q(
        \block[3][51] ) );
  EDFFXL \block_reg[3][15]  ( .D(block_next[15]), .E(n1176), .CK(clk), .Q(
        \block[3][15] ) );
  EDFFXL \block_reg[7][15]  ( .D(block_next[15]), .E(n1103), .CK(clk), .Q(
        \block[7][15] ) );
  EDFFXL \block_reg[3][11]  ( .D(block_next[11]), .E(n1175), .CK(clk), .QN(
        n516) );
  EDFFXL \block_reg[7][11]  ( .D(block_next[11]), .E(n1102), .CK(clk), .QN(
        n520) );
  EDFFXL \block_reg[3][14]  ( .D(block_next[14]), .E(n1176), .CK(clk), .Q(
        \block[3][14] ) );
  EDFFXL \block_reg[7][14]  ( .D(block_next[14]), .E(n1103), .CK(clk), .Q(
        \block[7][14] ) );
  EDFFXL \block_reg[3][111]  ( .D(block_next[111]), .E(n1183), .CK(clk), .Q(
        \block[3][111] ) );
  EDFFXL \block_reg[7][111]  ( .D(block_next[111]), .E(n1110), .CK(clk), .Q(
        \block[7][111] ) );
  EDFFXL \block_reg[3][79]  ( .D(block_next[79]), .E(n1181), .CK(clk), .QN(
        n456) );
  EDFFXL \block_reg[3][107]  ( .D(block_next[107]), .E(n1183), .CK(clk), .QN(
        n384) );
  EDFFXL \block_reg[7][79]  ( .D(block_next[79]), .E(n1108), .CK(clk), .QN(
        n460) );
  EDFFXL \block_reg[7][107]  ( .D(block_next[107]), .E(n1110), .CK(clk), .QN(
        n388) );
  EDFFXL \block_reg[3][110]  ( .D(block_next[110]), .E(n1183), .CK(clk), .QN(
        n432) );
  EDFFXL \block_reg[3][109]  ( .D(block_next[109]), .E(n1183), .CK(clk), .QN(
        n464) );
  EDFFXL \block_reg[7][110]  ( .D(block_next[110]), .E(n1110), .CK(clk), .QN(
        n436) );
  EDFFXL \block_reg[7][109]  ( .D(block_next[109]), .E(n1110), .CK(clk), .QN(
        n504) );
  EDFFXL \block_reg[3][75]  ( .D(block_next[75]), .E(n1180), .CK(clk), .QN(
        n336) );
  EDFFXL \block_reg[3][13]  ( .D(block_next[13]), .E(n1175), .CK(clk), .QN(
        n540) );
  EDFFXL \block_reg[7][75]  ( .D(block_next[75]), .E(n1107), .CK(clk), .QN(
        n340) );
  EDFFXL \block_reg[7][13]  ( .D(block_next[13]), .E(n1102), .CK(clk), .QN(
        n544) );
  EDFFXL \block_reg[3][12]  ( .D(block_next[12]), .E(n1175), .CK(clk), .QN(
        n532) );
  EDFFXL \block_reg[3][78]  ( .D(block_next[78]), .E(n1180), .CK(clk), .QN(
        n416) );
  EDFFXL \block_reg[7][12]  ( .D(block_next[12]), .E(n1102), .CK(clk), .QN(
        n536) );
  EDFFXL \block_reg[7][78]  ( .D(block_next[78]), .E(n1107), .CK(clk), .QN(
        n420) );
  EDFFXL \block_reg[3][10]  ( .D(block_next[10]), .E(n1175), .CK(clk), .QN(
        n508) );
  EDFFXL \block_reg[3][47]  ( .D(block_next[47]), .E(n1178), .CK(clk), .QN(
        n548) );
  EDFFXL \block_reg[3][8]  ( .D(block_next[8]), .E(n1175), .CK(clk), .Q(
        \block[3][8] ) );
  EDFFXL \block_reg[7][10]  ( .D(block_next[10]), .E(n1102), .CK(clk), .QN(
        n512) );
  EDFFXL \block_reg[7][47]  ( .D(block_next[47]), .E(n1105), .CK(clk), .QN(
        n552) );
  EDFFXL \block_reg[7][8]  ( .D(block_next[8]), .E(n1102), .CK(clk), .Q(
        \block[7][8] ) );
  EDFFXL \block_reg[3][43]  ( .D(block_next[43]), .E(n1178), .CK(clk), .QN(
        n352) );
  EDFFXL \block_reg[3][108]  ( .D(block_next[108]), .E(n1183), .CK(clk), .QN(
        n400) );
  EDFFXL \block_reg[7][108]  ( .D(block_next[108]), .E(n1110), .CK(clk), .QN(
        n404) );
  EDFFXL \block_reg[7][43]  ( .D(block_next[43]), .E(n1105), .CK(clk), .QN(
        n356) );
  EDFFXL \block_reg[3][44]  ( .D(block_next[44]), .E(n1178), .CK(clk), .QN(
        n368) );
  EDFFXL \block_reg[7][44]  ( .D(block_next[44]), .E(n1105), .CK(clk), .QN(
        n372) );
  EDFFXL \block_reg[3][106]  ( .D(block_next[106]), .E(n1183), .CK(clk), .QN(
        n376) );
  EDFFXL \block_reg[7][106]  ( .D(block_next[106]), .E(n1110), .CK(clk), .QN(
        n380) );
  EDFFXL \block_reg[3][46]  ( .D(block_next[46]), .E(n1178), .CK(clk), .Q(
        \block[3][46] ) );
  EDFFXL \block_reg[3][77]  ( .D(block_next[77]), .E(n1180), .CK(clk), .QN(
        n424) );
  EDFFXL \block_reg[3][76]  ( .D(block_next[76]), .E(n1180), .CK(clk), .QN(
        n448) );
  EDFFXL \block_reg[7][46]  ( .D(block_next[46]), .E(n1105), .CK(clk), .Q(
        \block[7][46] ) );
  EDFFXL \block_reg[7][77]  ( .D(block_next[77]), .E(n1107), .CK(clk), .QN(
        n428) );
  EDFFXL \block_reg[7][76]  ( .D(block_next[76]), .E(n1107), .CK(clk), .QN(
        n452) );
  EDFFXL \block_reg[3][104]  ( .D(block_next[104]), .E(n1182), .CK(clk), .Q(
        \block[3][104] ) );
  EDFFXL \block_reg[3][74]  ( .D(block_next[74]), .E(n1180), .CK(clk), .QN(
        n328) );
  EDFFXL \block_reg[7][104]  ( .D(block_next[104]), .E(n1109), .CK(clk), .Q(
        \block[7][104] ) );
  EDFFXL \block_reg[7][74]  ( .D(block_next[74]), .E(n1107), .CK(clk), .QN(
        n332) );
  EDFFXL \block_reg[3][9]  ( .D(block_next[9]), .E(n1175), .CK(clk), .QN(n524)
         );
  EDFFXL \block_reg[7][9]  ( .D(block_next[9]), .E(n1102), .CK(clk), .QN(n528)
         );
  EDFFXL \block_reg[3][45]  ( .D(block_next[45]), .E(n1178), .CK(clk), .QN(
        n408) );
  EDFFXL \block_reg[7][45]  ( .D(block_next[45]), .E(n1105), .CK(clk), .QN(
        n412) );
  EDFFXL \block_reg[3][42]  ( .D(block_next[42]), .E(n1178), .CK(clk), .QN(
        n440) );
  EDFFXL \block_reg[3][105]  ( .D(block_next[105]), .E(n1183), .CK(clk), .QN(
        n392) );
  EDFFXL \block_reg[7][42]  ( .D(block_next[42]), .E(n1105), .CK(clk), .QN(
        n444) );
  EDFFXL \block_reg[7][105]  ( .D(block_next[105]), .E(n1110), .CK(clk), .QN(
        n396) );
  EDFFXL \block_reg[3][73]  ( .D(block_next[73]), .E(n1180), .CK(clk), .QN(
        n344) );
  EDFFXL \block_reg[7][73]  ( .D(block_next[73]), .E(n1107), .CK(clk), .QN(
        n348) );
  EDFFXL \block_reg[3][72]  ( .D(block_next[72]), .E(n1180), .CK(clk), .Q(
        \block[3][72] ) );
  EDFFXL \block_reg[7][72]  ( .D(block_next[72]), .E(n1107), .CK(clk), .Q(
        \block[7][72] ) );
  EDFFXL \block_reg[3][41]  ( .D(block_next[41]), .E(n1178), .CK(clk), .QN(
        n360) );
  EDFFXL \block_reg[7][41]  ( .D(block_next[41]), .E(n1105), .CK(clk), .QN(
        n364) );
  EDFFXL \block_reg[3][40]  ( .D(block_next[40]), .E(n1178), .CK(clk), .Q(
        \block[3][40] ) );
  EDFFXL \block_reg[7][40]  ( .D(block_next[40]), .E(n1105), .CK(clk), .Q(
        \block[7][40] ) );
  EDFFXL \block_reg[3][6]  ( .D(block_next[6]), .E(n1175), .CK(clk), .Q(
        \block[3][6] ) );
  EDFFXL \block_reg[7][6]  ( .D(block_next[6]), .E(n1102), .CK(clk), .Q(
        \block[7][6] ) );
  EDFFXL \block_reg[3][102]  ( .D(block_next[102]), .E(n1182), .CK(clk), .Q(
        \block[3][102] ) );
  EDFFXL \block_reg[7][102]  ( .D(block_next[102]), .E(n1109), .CK(clk), .Q(
        \block[7][102] ) );
  EDFFXL \block_reg[3][70]  ( .D(block_next[70]), .E(n1180), .CK(clk), .Q(
        \block[3][70] ) );
  EDFFXL \block_reg[7][70]  ( .D(block_next[70]), .E(n1107), .CK(clk), .Q(
        \block[7][70] ) );
  EDFFXL \block_reg[3][38]  ( .D(block_next[38]), .E(n1177), .CK(clk), .Q(
        \block[3][38] ) );
  EDFFXL \block_reg[7][38]  ( .D(block_next[38]), .E(n1104), .CK(clk), .Q(
        \block[7][38] ) );
  EDFFXL \block_reg[3][0]  ( .D(block_next[0]), .E(n1174), .CK(clk), .Q(
        \block[3][0] ) );
  EDFFXL \block_reg[7][0]  ( .D(block_next[0]), .E(n1101), .CK(clk), .Q(
        \block[7][0] ) );
  EDFFXL \block_reg[3][96]  ( .D(block_next[96]), .E(n1182), .CK(clk), .Q(
        \block[3][96] ) );
  EDFFXL \block_reg[7][96]  ( .D(block_next[96]), .E(n1109), .CK(clk), .Q(
        \block[7][96] ) );
  EDFFXL \block_reg[3][64]  ( .D(block_next[64]), .E(n1179), .CK(clk), .Q(
        \block[3][64] ) );
  EDFFXL \block_reg[7][64]  ( .D(block_next[64]), .E(n1106), .CK(clk), .Q(
        \block[7][64] ) );
  EDFFXL \block_reg[3][32]  ( .D(block_next[32]), .E(n1177), .CK(clk), .Q(
        \block[3][32] ) );
  EDFFXL \block_reg[7][32]  ( .D(block_next[32]), .E(n1104), .CK(clk), .Q(
        \block[7][32] ) );
  EDFFXL \block_reg[3][5]  ( .D(block_next[5]), .E(n1175), .CK(clk), .QN(n312)
         );
  EDFFXL \block_reg[7][5]  ( .D(block_next[5]), .E(n1102), .CK(clk), .QN(n316)
         );
  EDFFXL \block_reg[3][7]  ( .D(block_next[7]), .E(n1175), .CK(clk), .Q(
        \block[3][7] ) );
  EDFFXL \block_reg[7][7]  ( .D(block_next[7]), .E(n1102), .CK(clk), .Q(
        \block[7][7] ) );
  EDFFXL \block_reg[3][3]  ( .D(block_next[3]), .E(n1175), .CK(clk), .Q(
        \block[3][3] ) );
  EDFFXL \block_reg[7][3]  ( .D(block_next[3]), .E(n1102), .CK(clk), .Q(
        \block[7][3] ) );
  EDFFXL \block_reg[3][4]  ( .D(block_next[4]), .E(n1175), .CK(clk), .Q(
        \block[3][4] ) );
  EDFFXL \block_reg[3][1]  ( .D(block_next[1]), .E(n1175), .CK(clk), .Q(
        \block[3][1] ) );
  EDFFXL \block_reg[7][4]  ( .D(block_next[4]), .E(n1102), .CK(clk), .Q(
        \block[7][4] ) );
  EDFFXL \block_reg[7][1]  ( .D(block_next[1]), .E(n1102), .CK(clk), .Q(
        \block[7][1] ) );
  EDFFXL \block_reg[3][2]  ( .D(block_next[2]), .E(n1175), .CK(clk), .Q(
        \block[3][2] ) );
  EDFFXL \block_reg[7][2]  ( .D(block_next[2]), .E(n1102), .CK(clk), .Q(
        \block[7][2] ) );
  EDFFXL \block_reg[3][103]  ( .D(block_next[103]), .E(n1182), .CK(clk), .Q(
        \block[3][103] ) );
  EDFFXL \block_reg[7][103]  ( .D(block_next[103]), .E(n1109), .CK(clk), .Q(
        \block[7][103] ) );
  EDFFXL \block_reg[3][101]  ( .D(block_next[101]), .E(n1182), .CK(clk), .Q(
        \block[3][101] ) );
  EDFFXL \block_reg[7][101]  ( .D(block_next[101]), .E(n1109), .CK(clk), .Q(
        \block[7][101] ) );
  EDFFXL \block_reg[3][71]  ( .D(block_next[71]), .E(n1180), .CK(clk), .Q(
        \block[3][71] ) );
  EDFFXL \block_reg[7][71]  ( .D(block_next[71]), .E(n1107), .CK(clk), .Q(
        \block[7][71] ) );
  EDFFXL \block_reg[3][68]  ( .D(block_next[68]), .E(n1180), .CK(clk), .Q(
        \block[3][68] ) );
  EDFFXL \block_reg[7][68]  ( .D(block_next[68]), .E(n1107), .CK(clk), .Q(
        \block[7][68] ) );
  EDFFXL \block_reg[3][67]  ( .D(block_next[67]), .E(n1180), .CK(clk), .Q(
        \block[3][67] ) );
  EDFFXL \block_reg[7][67]  ( .D(block_next[67]), .E(n1107), .CK(clk), .Q(
        \block[7][67] ) );
  EDFFXL \block_reg[3][37]  ( .D(block_next[37]), .E(n1177), .CK(clk), .Q(
        \block[3][37] ) );
  EDFFXL \block_reg[3][39]  ( .D(block_next[39]), .E(n1177), .CK(clk), .Q(
        \block[3][39] ) );
  EDFFXL \block_reg[7][37]  ( .D(block_next[37]), .E(n1104), .CK(clk), .Q(
        \block[7][37] ) );
  EDFFXL \block_reg[7][39]  ( .D(block_next[39]), .E(n1104), .CK(clk), .Q(
        \block[7][39] ) );
  EDFFXL \block_reg[3][69]  ( .D(block_next[69]), .E(n1180), .CK(clk), .Q(
        \block[3][69] ) );
  EDFFXL \block_reg[3][100]  ( .D(block_next[100]), .E(n1182), .CK(clk), .Q(
        \block[3][100] ) );
  EDFFXL \block_reg[7][69]  ( .D(block_next[69]), .E(n1107), .CK(clk), .Q(
        \block[7][69] ) );
  EDFFXL \block_reg[7][100]  ( .D(block_next[100]), .E(n1109), .CK(clk), .Q(
        \block[7][100] ) );
  EDFFXL \block_reg[3][99]  ( .D(block_next[99]), .E(n1182), .CK(clk), .Q(
        \block[3][99] ) );
  EDFFXL \block_reg[7][99]  ( .D(block_next[99]), .E(n1109), .CK(clk), .Q(
        \block[7][99] ) );
  EDFFXL \block_reg[3][97]  ( .D(block_next[97]), .E(n1182), .CK(clk), .Q(
        \block[3][97] ) );
  EDFFXL \block_reg[7][97]  ( .D(block_next[97]), .E(n1109), .CK(clk), .Q(
        \block[7][97] ) );
  EDFFXL \block_reg[3][65]  ( .D(block_next[65]), .E(n1179), .CK(clk), .Q(
        \block[3][65] ) );
  EDFFXL \block_reg[7][65]  ( .D(block_next[65]), .E(n1106), .CK(clk), .Q(
        \block[7][65] ) );
  EDFFXL \block_reg[3][98]  ( .D(block_next[98]), .E(n1182), .CK(clk), .Q(
        \block[3][98] ) );
  EDFFXL \block_reg[3][36]  ( .D(block_next[36]), .E(n1177), .CK(clk), .QN(
        n320) );
  EDFFXL \block_reg[7][36]  ( .D(block_next[36]), .E(n1104), .CK(clk), .QN(
        n324) );
  EDFFXL \block_reg[7][98]  ( .D(block_next[98]), .E(n1109), .CK(clk), .Q(
        \block[7][98] ) );
  EDFFXL \block_reg[3][66]  ( .D(block_next[66]), .E(n1180), .CK(clk), .Q(
        \block[3][66] ) );
  EDFFXL \block_reg[7][66]  ( .D(block_next[66]), .E(n1107), .CK(clk), .Q(
        \block[7][66] ) );
  EDFFXL \block_reg[3][35]  ( .D(block_next[35]), .E(n1177), .CK(clk), .Q(
        \block[3][35] ) );
  EDFFXL \block_reg[7][35]  ( .D(block_next[35]), .E(n1104), .CK(clk), .Q(
        \block[7][35] ) );
  EDFFXL \block_reg[3][33]  ( .D(block_next[33]), .E(n1177), .CK(clk), .Q(
        \block[3][33] ) );
  EDFFXL \block_reg[7][33]  ( .D(block_next[33]), .E(n1104), .CK(clk), .Q(
        \block[7][33] ) );
  EDFFXL \block_reg[3][34]  ( .D(block_next[34]), .E(n1177), .CK(clk), .Q(
        \block[3][34] ) );
  EDFFXL \block_reg[7][34]  ( .D(block_next[34]), .E(n1104), .CK(clk), .Q(
        \block[7][34] ) );
  EDFFXL \block_reg[3][122]  ( .D(block_next[122]), .E(n1184), .CK(clk), .Q(
        \block[3][122] ) );
  EDFFXL \block_reg[7][122]  ( .D(block_next[122]), .E(n1111), .CK(clk), .Q(
        \block[7][122] ) );
  EDFFXL \block_reg[3][26]  ( .D(block_next[26]), .E(n1176), .CK(clk), .QN(
        n294) );
  EDFFXL \block_reg[7][26]  ( .D(block_next[26]), .E(n1103), .CK(clk), .QN(
        n298) );
  EDFFXL \block_reg[5][116]  ( .D(block_next[116]), .E(n1145), .CK(clk), .Q(
        \block[5][116] ) );
  EDFFXL \block_reg[5][112]  ( .D(block_next[112]), .E(n1145), .CK(clk), .Q(
        \block[5][112] ) );
  EDFFXL \block_reg[5][89]  ( .D(block_next[89]), .E(n1143), .CK(clk), .Q(
        \block[5][89] ) );
  EDFFXL \block_reg[5][88]  ( .D(block_next[88]), .E(n1143), .CK(clk), .Q(
        \block[5][88] ) );
  EDFFXL \block_reg[5][87]  ( .D(block_next[87]), .E(n1143), .CK(clk), .Q(
        \block[5][87] ) );
  EDFFXL \block_reg[5][86]  ( .D(block_next[86]), .E(n1143), .CK(clk), .Q(
        \block[5][86] ) );
  EDFFXL \block_reg[5][85]  ( .D(block_next[85]), .E(n1143), .CK(clk), .Q(
        \block[5][85] ) );
  EDFFXL \block_reg[5][84]  ( .D(block_next[84]), .E(n1143), .CK(clk), .Q(
        \block[5][84] ) );
  EDFFXL \block_reg[5][83]  ( .D(block_next[83]), .E(n1143), .CK(clk), .Q(
        \block[5][83] ) );
  EDFFXL \block_reg[5][82]  ( .D(block_next[82]), .E(n1143), .CK(clk), .Q(
        \block[5][82] ) );
  EDFFXL \block_reg[5][81]  ( .D(block_next[81]), .E(n1143), .CK(clk), .Q(
        \block[5][81] ) );
  EDFFXL \block_reg[5][80]  ( .D(block_next[80]), .E(n1143), .CK(clk), .Q(
        \block[5][80] ) );
  EDFFXL \block_reg[5][57]  ( .D(block_next[57]), .E(n1141), .CK(clk), .Q(
        \block[5][57] ) );
  EDFFXL \block_reg[5][25]  ( .D(block_next[25]), .E(n1138), .CK(clk), .Q(
        \block[5][25] ) );
  EDFFXL \block_reg[5][24]  ( .D(block_next[24]), .E(n1138), .CK(clk), .Q(
        \block[5][24] ) );
  EDFFXL \block_reg[5][23]  ( .D(block_next[23]), .E(n1138), .CK(clk), .Q(
        \block[5][23] ) );
  EDFFXL \block_reg[5][22]  ( .D(block_next[22]), .E(n1138), .CK(clk), .Q(
        \block[5][22] ) );
  EDFFXL \block_reg[5][21]  ( .D(block_next[21]), .E(n1138), .CK(clk), .Q(
        \block[5][21] ) );
  EDFFXL \block_reg[5][18]  ( .D(block_next[18]), .E(n1138), .CK(clk), .Q(
        \block[5][18] ) );
  EDFFXL \block_reg[5][16]  ( .D(block_next[16]), .E(n1138), .CK(clk), .Q(
        \block[5][16] ) );
  EDFFXL \block_reg[5][121]  ( .D(block_next[121]), .E(n1146), .CK(clk), .Q(
        \block[5][121] ) );
  EDFFXL \block_reg[5][120]  ( .D(block_next[120]), .E(n1146), .CK(clk), .Q(
        \block[5][120] ) );
  EDFFXL \block_reg[5][119]  ( .D(block_next[119]), .E(n1146), .CK(clk), .Q(
        \block[5][119] ) );
  EDFFXL \block_reg[5][118]  ( .D(block_next[118]), .E(n1146), .CK(clk), .Q(
        \block[5][118] ) );
  EDFFXL \block_reg[5][117]  ( .D(block_next[117]), .E(n1145), .CK(clk), .Q(
        \block[5][117] ) );
  EDFFXL \block_reg[5][48]  ( .D(block_next[48]), .E(n1140), .CK(clk), .Q(
        \block[5][48] ) );
  EDFFXL \block_reg[5][115]  ( .D(block_next[115]), .E(n1145), .CK(clk), .Q(
        \block[5][115] ) );
  EDFFXL \block_reg[5][114]  ( .D(block_next[114]), .E(n1145), .CK(clk), .Q(
        \block[5][114] ) );
  EDFFXL \block_reg[5][113]  ( .D(block_next[113]), .E(n1145), .CK(clk), .Q(
        \block[5][113] ) );
  EDFFXL \block_reg[1][116]  ( .D(block_next[116]), .E(n1221), .CK(clk), .Q(
        \block[1][116] ) );
  EDFFXL \block_reg[1][112]  ( .D(block_next[112]), .E(n1221), .CK(clk), .Q(
        \block[1][112] ) );
  EDFFXL \block_reg[1][89]  ( .D(block_next[89]), .E(n1219), .CK(clk), .Q(
        \block[1][89] ) );
  EDFFXL \block_reg[1][88]  ( .D(block_next[88]), .E(n1219), .CK(clk), .Q(
        \block[1][88] ) );
  EDFFXL \block_reg[1][87]  ( .D(block_next[87]), .E(n1219), .CK(clk), .Q(
        \block[1][87] ) );
  EDFFXL \block_reg[1][86]  ( .D(block_next[86]), .E(n1219), .CK(clk), .Q(
        \block[1][86] ) );
  EDFFXL \block_reg[1][85]  ( .D(block_next[85]), .E(n1219), .CK(clk), .Q(
        \block[1][85] ) );
  EDFFXL \block_reg[1][84]  ( .D(block_next[84]), .E(n1219), .CK(clk), .Q(
        \block[1][84] ) );
  EDFFXL \block_reg[1][83]  ( .D(block_next[83]), .E(n1219), .CK(clk), .Q(
        \block[1][83] ) );
  EDFFXL \block_reg[1][82]  ( .D(block_next[82]), .E(n1219), .CK(clk), .Q(
        \block[1][82] ) );
  EDFFXL \block_reg[1][81]  ( .D(block_next[81]), .E(n1219), .CK(clk), .Q(
        \block[1][81] ) );
  EDFFXL \block_reg[1][80]  ( .D(block_next[80]), .E(n1219), .CK(clk), .Q(
        \block[1][80] ) );
  EDFFXL \block_reg[1][57]  ( .D(block_next[57]), .E(n1217), .CK(clk), .Q(
        \block[1][57] ) );
  EDFFXL \block_reg[1][25]  ( .D(block_next[25]), .E(n1214), .CK(clk), .Q(
        \block[1][25] ) );
  EDFFXL \block_reg[1][24]  ( .D(block_next[24]), .E(n1214), .CK(clk), .Q(
        \block[1][24] ) );
  EDFFXL \block_reg[1][23]  ( .D(block_next[23]), .E(n1214), .CK(clk), .Q(
        \block[1][23] ) );
  EDFFXL \block_reg[1][22]  ( .D(block_next[22]), .E(n1214), .CK(clk), .Q(
        \block[1][22] ) );
  EDFFXL \block_reg[1][21]  ( .D(block_next[21]), .E(n1214), .CK(clk), .Q(
        \block[1][21] ) );
  EDFFXL \block_reg[1][18]  ( .D(block_next[18]), .E(n1214), .CK(clk), .Q(
        \block[1][18] ) );
  EDFFXL \block_reg[1][16]  ( .D(block_next[16]), .E(n1214), .CK(clk), .Q(
        \block[1][16] ) );
  EDFFXL \block_reg[5][17]  ( .D(block_next[17]), .E(n1138), .CK(clk), .Q(
        \block[5][17] ) );
  EDFFXL \block_reg[1][121]  ( .D(block_next[121]), .E(n1222), .CK(clk), .Q(
        \block[1][121] ) );
  EDFFXL \block_reg[1][120]  ( .D(block_next[120]), .E(n1222), .CK(clk), .Q(
        \block[1][120] ) );
  EDFFXL \block_reg[1][119]  ( .D(block_next[119]), .E(n1222), .CK(clk), .Q(
        \block[1][119] ) );
  EDFFXL \block_reg[1][118]  ( .D(block_next[118]), .E(n1222), .CK(clk), .Q(
        \block[1][118] ) );
  EDFFXL \block_reg[1][117]  ( .D(block_next[117]), .E(n1221), .CK(clk), .Q(
        \block[1][117] ) );
  EDFFXL \block_reg[1][48]  ( .D(block_next[48]), .E(n1216), .CK(clk), .Q(
        \block[1][48] ) );
  EDFFXL \block_reg[5][20]  ( .D(block_next[20]), .E(n1138), .CK(clk), .Q(
        \block[5][20] ) );
  EDFFXL \block_reg[5][19]  ( .D(block_next[19]), .E(n1138), .CK(clk), .Q(
        \block[5][19] ) );
  EDFFXL \block_reg[5][50]  ( .D(block_next[50]), .E(n1140), .CK(clk), .Q(
        \block[5][50] ) );
  EDFFXL \block_reg[5][49]  ( .D(block_next[49]), .E(n1140), .CK(clk), .Q(
        \block[5][49] ) );
  EDFFXL \block_reg[5][56]  ( .D(block_next[56]), .E(n1141), .CK(clk), .Q(
        \block[5][56] ) );
  EDFFXL \block_reg[5][55]  ( .D(block_next[55]), .E(n1141), .CK(clk), .Q(
        \block[5][55] ) );
  EDFFXL \block_reg[5][54]  ( .D(block_next[54]), .E(n1141), .CK(clk), .Q(
        \block[5][54] ) );
  EDFFXL \block_reg[5][53]  ( .D(block_next[53]), .E(n1141), .CK(clk), .Q(
        \block[5][53] ) );
  EDFFXL \block_reg[5][52]  ( .D(block_next[52]), .E(n1140), .CK(clk), .Q(
        \block[5][52] ) );
  EDFFXL \block_reg[5][51]  ( .D(block_next[51]), .E(n1140), .CK(clk), .Q(
        \block[5][51] ) );
  EDFFXL \block_reg[1][115]  ( .D(block_next[115]), .E(n1221), .CK(clk), .Q(
        \block[1][115] ) );
  EDFFXL \block_reg[1][114]  ( .D(block_next[114]), .E(n1221), .CK(clk), .Q(
        \block[1][114] ) );
  EDFFXL \block_reg[1][113]  ( .D(block_next[113]), .E(n1221), .CK(clk), .Q(
        \block[1][113] ) );
  EDFFXL \block_reg[1][17]  ( .D(block_next[17]), .E(n1214), .CK(clk), .Q(
        \block[1][17] ) );
  EDFFXL \block_reg[1][20]  ( .D(block_next[20]), .E(n1214), .CK(clk), .Q(
        \block[1][20] ) );
  EDFFXL \block_reg[1][19]  ( .D(block_next[19]), .E(n1214), .CK(clk), .Q(
        \block[1][19] ) );
  EDFFXL \block_reg[1][50]  ( .D(block_next[50]), .E(n1216), .CK(clk), .Q(
        \block[1][50] ) );
  EDFFXL \block_reg[1][49]  ( .D(block_next[49]), .E(n1216), .CK(clk), .Q(
        \block[1][49] ) );
  EDFFXL \block_reg[1][56]  ( .D(block_next[56]), .E(n1217), .CK(clk), .Q(
        \block[1][56] ) );
  EDFFXL \block_reg[1][55]  ( .D(block_next[55]), .E(n1217), .CK(clk), .Q(
        \block[1][55] ) );
  EDFFXL \block_reg[1][54]  ( .D(block_next[54]), .E(n1217), .CK(clk), .Q(
        \block[1][54] ) );
  EDFFXL \block_reg[1][53]  ( .D(block_next[53]), .E(n1217), .CK(clk), .Q(
        \block[1][53] ) );
  EDFFXL \block_reg[1][52]  ( .D(block_next[52]), .E(n1216), .CK(clk), .Q(
        \block[1][52] ) );
  EDFFXL \block_reg[1][51]  ( .D(block_next[51]), .E(n1216), .CK(clk), .Q(
        \block[1][51] ) );
  EDFFXL \block_reg[5][15]  ( .D(block_next[15]), .E(n1138), .CK(clk), .Q(
        \block[5][15] ) );
  EDFFXL \block_reg[1][15]  ( .D(block_next[15]), .E(n1214), .CK(clk), .Q(
        \block[1][15] ) );
  EDFFXL \block_reg[1][11]  ( .D(block_next[11]), .E(n1213), .CK(clk), .QN(
        n514) );
  EDFFXL \block_reg[5][11]  ( .D(block_next[11]), .E(n1137), .CK(clk), .QN(
        n518) );
  EDFFXL \block_reg[1][14]  ( .D(block_next[14]), .E(n1214), .CK(clk), .Q(
        \block[1][14] ) );
  EDFFXL \block_reg[5][14]  ( .D(block_next[14]), .E(n1138), .CK(clk), .Q(
        \block[5][14] ) );
  EDFFXL \block_reg[1][111]  ( .D(block_next[111]), .E(n1221), .CK(clk), .Q(
        \block[1][111] ) );
  EDFFXL \block_reg[5][111]  ( .D(block_next[111]), .E(n1145), .CK(clk), .Q(
        \block[5][111] ) );
  EDFFXL \block_reg[1][79]  ( .D(block_next[79]), .E(n1219), .CK(clk), .QN(
        n454) );
  EDFFXL \block_reg[1][107]  ( .D(block_next[107]), .E(n1221), .CK(clk), .QN(
        n382) );
  EDFFXL \block_reg[5][79]  ( .D(block_next[79]), .E(n1143), .CK(clk), .QN(
        n458) );
  EDFFXL \block_reg[5][107]  ( .D(block_next[107]), .E(n1145), .CK(clk), .QN(
        n386) );
  EDFFXL \block_reg[1][110]  ( .D(block_next[110]), .E(n1221), .CK(clk), .QN(
        n430) );
  EDFFXL \block_reg[1][109]  ( .D(block_next[109]), .E(n1221), .CK(clk), .QN(
        n462) );
  EDFFXL \block_reg[5][109]  ( .D(block_next[109]), .E(n1145), .CK(clk), .QN(
        n466) );
  EDFFXL \block_reg[5][110]  ( .D(block_next[110]), .E(n1145), .CK(clk), .QN(
        n434) );
  EDFFXL \block_reg[1][75]  ( .D(block_next[75]), .E(n1218), .CK(clk), .QN(
        n334) );
  EDFFXL \block_reg[1][13]  ( .D(block_next[13]), .E(n1213), .CK(clk), .QN(
        n538) );
  EDFFXL \block_reg[5][75]  ( .D(block_next[75]), .E(n1142), .CK(clk), .QN(
        n338) );
  EDFFXL \block_reg[5][13]  ( .D(block_next[13]), .E(n1137), .CK(clk), .QN(
        n542) );
  EDFFXL \block_reg[1][12]  ( .D(block_next[12]), .E(n1213), .CK(clk), .QN(
        n530) );
  EDFFXL \block_reg[1][78]  ( .D(block_next[78]), .E(n1218), .CK(clk), .QN(
        n414) );
  EDFFXL \block_reg[5][78]  ( .D(block_next[78]), .E(n1142), .CK(clk), .QN(
        n418) );
  EDFFXL \block_reg[5][12]  ( .D(block_next[12]), .E(n1137), .CK(clk), .QN(
        n534) );
  EDFFXL \block_reg[1][8]  ( .D(block_next[8]), .E(n1213), .CK(clk), .Q(
        \block[1][8] ) );
  EDFFXL \block_reg[1][10]  ( .D(block_next[10]), .E(n1213), .CK(clk), .QN(
        n506) );
  EDFFXL \block_reg[1][47]  ( .D(block_next[47]), .E(n1216), .CK(clk), .QN(
        n546) );
  EDFFXL \block_reg[5][8]  ( .D(block_next[8]), .E(n1137), .CK(clk), .Q(
        \block[5][8] ) );
  EDFFXL \block_reg[5][10]  ( .D(block_next[10]), .E(n1137), .CK(clk), .QN(
        n510) );
  EDFFXL \block_reg[5][47]  ( .D(block_next[47]), .E(n1140), .CK(clk), .QN(
        n550) );
  EDFFXL \block_reg[1][108]  ( .D(block_next[108]), .E(n1221), .CK(clk), .QN(
        n398) );
  EDFFXL \block_reg[1][43]  ( .D(block_next[43]), .E(n1216), .CK(clk), .QN(
        n350) );
  EDFFXL \block_reg[1][44]  ( .D(block_next[44]), .E(n1216), .CK(clk), .QN(
        n366) );
  EDFFXL \block_reg[5][108]  ( .D(block_next[108]), .E(n1145), .CK(clk), .QN(
        n402) );
  EDFFXL \block_reg[5][43]  ( .D(block_next[43]), .E(n1140), .CK(clk), .QN(
        n354) );
  EDFFXL \block_reg[5][44]  ( .D(block_next[44]), .E(n1140), .CK(clk), .QN(
        n370) );
  EDFFXL \block_reg[1][106]  ( .D(block_next[106]), .E(n1221), .CK(clk), .QN(
        n374) );
  EDFFXL \block_reg[5][106]  ( .D(block_next[106]), .E(n1145), .CK(clk), .QN(
        n378) );
  EDFFXL \block_reg[1][46]  ( .D(block_next[46]), .E(n1216), .CK(clk), .Q(
        \block[1][46] ) );
  EDFFXL \block_reg[1][77]  ( .D(block_next[77]), .E(n1218), .CK(clk), .QN(
        n422) );
  EDFFXL \block_reg[1][76]  ( .D(block_next[76]), .E(n1218), .CK(clk), .QN(
        n446) );
  EDFFXL \block_reg[5][77]  ( .D(block_next[77]), .E(n1142), .CK(clk), .QN(
        n426) );
  EDFFXL \block_reg[5][46]  ( .D(block_next[46]), .E(n1140), .CK(clk), .Q(
        \block[5][46] ) );
  EDFFXL \block_reg[5][76]  ( .D(block_next[76]), .E(n1142), .CK(clk), .QN(
        n450) );
  EDFFXL \block_reg[1][104]  ( .D(block_next[104]), .E(n1220), .CK(clk), .Q(
        \block[1][104] ) );
  EDFFXL \block_reg[5][104]  ( .D(block_next[104]), .E(n1144), .CK(clk), .Q(
        \block[5][104] ) );
  EDFFXL \block_reg[1][74]  ( .D(block_next[74]), .E(n1218), .CK(clk), .QN(
        n326) );
  EDFFXL \block_reg[5][74]  ( .D(block_next[74]), .E(n1142), .CK(clk), .QN(
        n330) );
  EDFFXL \block_reg[1][9]  ( .D(block_next[9]), .E(n1213), .CK(clk), .QN(n522)
         );
  EDFFXL \block_reg[5][9]  ( .D(block_next[9]), .E(n1137), .CK(clk), .QN(n526)
         );
  EDFFXL \block_reg[1][45]  ( .D(block_next[45]), .E(n1216), .CK(clk), .QN(
        n406) );
  EDFFXL \block_reg[5][45]  ( .D(block_next[45]), .E(n1140), .CK(clk), .QN(
        n410) );
  EDFFXL \block_reg[1][42]  ( .D(block_next[42]), .E(n1216), .CK(clk), .QN(
        n438) );
  EDFFXL \block_reg[1][105]  ( .D(block_next[105]), .E(n1221), .CK(clk), .QN(
        n390) );
  EDFFXL \block_reg[5][42]  ( .D(block_next[42]), .E(n1140), .CK(clk), .QN(
        n442) );
  EDFFXL \block_reg[5][105]  ( .D(block_next[105]), .E(n1145), .CK(clk), .QN(
        n394) );
  EDFFXL \block_reg[1][73]  ( .D(block_next[73]), .E(n1218), .CK(clk), .QN(
        n342) );
  EDFFXL \block_reg[5][73]  ( .D(block_next[73]), .E(n1142), .CK(clk), .QN(
        n346) );
  EDFFXL \block_reg[1][72]  ( .D(block_next[72]), .E(n1218), .CK(clk), .Q(
        \block[1][72] ) );
  EDFFXL \block_reg[5][72]  ( .D(block_next[72]), .E(n1142), .CK(clk), .Q(
        \block[5][72] ) );
  EDFFXL \block_reg[1][41]  ( .D(block_next[41]), .E(n1216), .CK(clk), .QN(
        n358) );
  EDFFXL \block_reg[5][41]  ( .D(block_next[41]), .E(n1140), .CK(clk), .QN(
        n362) );
  EDFFXL \block_reg[1][40]  ( .D(block_next[40]), .E(n1216), .CK(clk), .Q(
        \block[1][40] ) );
  EDFFXL \block_reg[5][40]  ( .D(block_next[40]), .E(n1140), .CK(clk), .Q(
        \block[5][40] ) );
  EDFFXL \block_reg[1][6]  ( .D(block_next[6]), .E(n1213), .CK(clk), .Q(
        \block[1][6] ) );
  EDFFXL \block_reg[5][6]  ( .D(block_next[6]), .E(n1137), .CK(clk), .Q(
        \block[5][6] ) );
  EDFFXL \block_reg[1][102]  ( .D(block_next[102]), .E(n1220), .CK(clk), .Q(
        \block[1][102] ) );
  EDFFXL \block_reg[5][102]  ( .D(block_next[102]), .E(n1144), .CK(clk), .Q(
        \block[5][102] ) );
  EDFFXL \block_reg[1][70]  ( .D(block_next[70]), .E(n1218), .CK(clk), .Q(
        \block[1][70] ) );
  EDFFXL \block_reg[5][70]  ( .D(block_next[70]), .E(n1142), .CK(clk), .Q(
        \block[5][70] ) );
  EDFFXL \block_reg[1][38]  ( .D(block_next[38]), .E(n1215), .CK(clk), .Q(
        \block[1][38] ) );
  EDFFXL \block_reg[5][38]  ( .D(block_next[38]), .E(n1139), .CK(clk), .Q(
        \block[5][38] ) );
  EDFFXL \block_reg[1][0]  ( .D(block_next[0]), .E(n1212), .CK(clk), .Q(
        \block[1][0] ) );
  EDFFXL \block_reg[5][0]  ( .D(block_next[0]), .E(n1136), .CK(clk), .Q(
        \block[5][0] ) );
  EDFFXL \block_reg[1][96]  ( .D(block_next[96]), .E(n1220), .CK(clk), .Q(
        \block[1][96] ) );
  EDFFXL \block_reg[5][96]  ( .D(block_next[96]), .E(n1144), .CK(clk), .Q(
        \block[5][96] ) );
  EDFFXL \block_reg[1][64]  ( .D(block_next[64]), .E(n1217), .CK(clk), .Q(
        \block[1][64] ) );
  EDFFXL \block_reg[5][64]  ( .D(block_next[64]), .E(n1141), .CK(clk), .Q(
        \block[5][64] ) );
  EDFFXL \block_reg[1][32]  ( .D(block_next[32]), .E(n1215), .CK(clk), .Q(
        \block[1][32] ) );
  EDFFXL \block_reg[5][32]  ( .D(block_next[32]), .E(n1139), .CK(clk), .Q(
        \block[5][32] ) );
  EDFFXL \block_reg[1][5]  ( .D(block_next[5]), .E(n1213), .CK(clk), .QN(n310)
         );
  EDFFXL \block_reg[5][5]  ( .D(block_next[5]), .E(n1137), .CK(clk), .QN(n314)
         );
  EDFFXL \block_reg[1][7]  ( .D(block_next[7]), .E(n1213), .CK(clk), .Q(
        \block[1][7] ) );
  EDFFXL \block_reg[5][7]  ( .D(block_next[7]), .E(n1137), .CK(clk), .Q(
        \block[5][7] ) );
  EDFFXL \block_reg[1][3]  ( .D(block_next[3]), .E(n1213), .CK(clk), .Q(
        \block[1][3] ) );
  EDFFXL \block_reg[5][3]  ( .D(block_next[3]), .E(n1137), .CK(clk), .Q(
        \block[5][3] ) );
  EDFFXL \block_reg[1][4]  ( .D(block_next[4]), .E(n1213), .CK(clk), .Q(
        \block[1][4] ) );
  EDFFXL \block_reg[1][1]  ( .D(block_next[1]), .E(n1213), .CK(clk), .Q(
        \block[1][1] ) );
  EDFFXL \block_reg[5][4]  ( .D(block_next[4]), .E(n1137), .CK(clk), .Q(
        \block[5][4] ) );
  EDFFXL \block_reg[5][1]  ( .D(block_next[1]), .E(n1137), .CK(clk), .Q(
        \block[5][1] ) );
  EDFFXL \block_reg[1][2]  ( .D(block_next[2]), .E(n1213), .CK(clk), .Q(
        \block[1][2] ) );
  EDFFXL \block_reg[5][2]  ( .D(block_next[2]), .E(n1137), .CK(clk), .Q(
        \block[5][2] ) );
  EDFFXL \block_reg[1][103]  ( .D(block_next[103]), .E(n1220), .CK(clk), .Q(
        \block[1][103] ) );
  EDFFXL \block_reg[5][103]  ( .D(block_next[103]), .E(n1144), .CK(clk), .Q(
        \block[5][103] ) );
  EDFFXL \block_reg[1][101]  ( .D(block_next[101]), .E(n1220), .CK(clk), .Q(
        \block[1][101] ) );
  EDFFXL \block_reg[5][101]  ( .D(block_next[101]), .E(n1144), .CK(clk), .Q(
        \block[5][101] ) );
  EDFFXL \block_reg[1][71]  ( .D(block_next[71]), .E(n1218), .CK(clk), .Q(
        \block[1][71] ) );
  EDFFXL \block_reg[5][71]  ( .D(block_next[71]), .E(n1142), .CK(clk), .Q(
        \block[5][71] ) );
  EDFFXL \block_reg[1][68]  ( .D(block_next[68]), .E(n1218), .CK(clk), .Q(
        \block[1][68] ) );
  EDFFXL \block_reg[5][68]  ( .D(block_next[68]), .E(n1142), .CK(clk), .Q(
        \block[5][68] ) );
  EDFFXL \block_reg[1][67]  ( .D(block_next[67]), .E(n1218), .CK(clk), .Q(
        \block[1][67] ) );
  EDFFXL \block_reg[1][37]  ( .D(block_next[37]), .E(n1215), .CK(clk), .Q(
        \block[1][37] ) );
  EDFFXL \block_reg[5][67]  ( .D(block_next[67]), .E(n1142), .CK(clk), .Q(
        \block[5][67] ) );
  EDFFXL \block_reg[5][37]  ( .D(block_next[37]), .E(n1139), .CK(clk), .Q(
        \block[5][37] ) );
  EDFFXL \block_reg[1][39]  ( .D(block_next[39]), .E(n1215), .CK(clk), .Q(
        \block[1][39] ) );
  EDFFXL \block_reg[5][39]  ( .D(block_next[39]), .E(n1139), .CK(clk), .Q(
        \block[5][39] ) );
  EDFFXL \block_reg[1][69]  ( .D(block_next[69]), .E(n1218), .CK(clk), .Q(
        \block[1][69] ) );
  EDFFXL \block_reg[1][100]  ( .D(block_next[100]), .E(n1220), .CK(clk), .Q(
        \block[1][100] ) );
  EDFFXL \block_reg[5][69]  ( .D(block_next[69]), .E(n1142), .CK(clk), .Q(
        \block[5][69] ) );
  EDFFXL \block_reg[5][100]  ( .D(block_next[100]), .E(n1144), .CK(clk), .Q(
        \block[5][100] ) );
  EDFFXL \block_reg[1][99]  ( .D(block_next[99]), .E(n1220), .CK(clk), .Q(
        \block[1][99] ) );
  EDFFXL \block_reg[1][97]  ( .D(block_next[97]), .E(n1220), .CK(clk), .Q(
        \block[1][97] ) );
  EDFFXL \block_reg[5][99]  ( .D(block_next[99]), .E(n1144), .CK(clk), .Q(
        \block[5][99] ) );
  EDFFXL \block_reg[5][97]  ( .D(block_next[97]), .E(n1144), .CK(clk), .Q(
        \block[5][97] ) );
  EDFFXL \block_reg[1][65]  ( .D(block_next[65]), .E(n1217), .CK(clk), .Q(
        \block[1][65] ) );
  EDFFXL \block_reg[5][65]  ( .D(block_next[65]), .E(n1141), .CK(clk), .Q(
        \block[5][65] ) );
  EDFFXL \block_reg[1][36]  ( .D(block_next[36]), .E(n1215), .CK(clk), .QN(
        n318) );
  EDFFXL \block_reg[1][98]  ( .D(block_next[98]), .E(n1220), .CK(clk), .Q(
        \block[1][98] ) );
  EDFFXL \block_reg[5][36]  ( .D(block_next[36]), .E(n1139), .CK(clk), .QN(
        n322) );
  EDFFXL \block_reg[5][98]  ( .D(block_next[98]), .E(n1144), .CK(clk), .Q(
        \block[5][98] ) );
  EDFFXL \block_reg[1][66]  ( .D(block_next[66]), .E(n1218), .CK(clk), .Q(
        \block[1][66] ) );
  EDFFXL \block_reg[5][66]  ( .D(block_next[66]), .E(n1142), .CK(clk), .Q(
        \block[5][66] ) );
  EDFFXL \block_reg[1][35]  ( .D(block_next[35]), .E(n1215), .CK(clk), .Q(
        \block[1][35] ) );
  EDFFXL \block_reg[5][35]  ( .D(block_next[35]), .E(n1139), .CK(clk), .Q(
        \block[5][35] ) );
  EDFFXL \block_reg[1][33]  ( .D(block_next[33]), .E(n1215), .CK(clk), .Q(
        \block[1][33] ) );
  EDFFXL \block_reg[5][33]  ( .D(block_next[33]), .E(n1139), .CK(clk), .Q(
        \block[5][33] ) );
  EDFFXL \block_reg[1][34]  ( .D(block_next[34]), .E(n1215), .CK(clk), .Q(
        \block[1][34] ) );
  EDFFXL \block_reg[5][34]  ( .D(block_next[34]), .E(n1139), .CK(clk), .Q(
        \block[5][34] ) );
  EDFFXL \block_reg[1][122]  ( .D(block_next[122]), .E(n1222), .CK(clk), .Q(
        \block[1][122] ) );
  EDFFXL \block_reg[5][122]  ( .D(block_next[122]), .E(n1146), .CK(clk), .Q(
        \block[5][122] ) );
  EDFFXL \block_reg[1][26]  ( .D(block_next[26]), .E(n1214), .CK(clk), .QN(
        n292) );
  EDFFXL \block_reg[5][26]  ( .D(block_next[26]), .E(n1138), .CK(clk), .QN(
        n296) );
  EDFFXL \block_reg[4][116]  ( .D(block_next[116]), .E(n1164), .CK(clk), .Q(
        \block[4][116] ) );
  EDFFXL \block_reg[4][112]  ( .D(block_next[112]), .E(n1164), .CK(clk), .Q(
        \block[4][112] ) );
  EDFFXL \block_reg[4][89]  ( .D(block_next[89]), .E(n1162), .CK(clk), .Q(
        \block[4][89] ) );
  EDFFXL \block_reg[4][88]  ( .D(block_next[88]), .E(n1162), .CK(clk), .Q(
        \block[4][88] ) );
  EDFFXL \block_reg[4][87]  ( .D(block_next[87]), .E(n1162), .CK(clk), .Q(
        \block[4][87] ) );
  EDFFXL \block_reg[4][86]  ( .D(block_next[86]), .E(n1162), .CK(clk), .Q(
        \block[4][86] ) );
  EDFFXL \block_reg[4][85]  ( .D(block_next[85]), .E(n1162), .CK(clk), .Q(
        \block[4][85] ) );
  EDFFXL \block_reg[4][84]  ( .D(block_next[84]), .E(n1162), .CK(clk), .Q(
        \block[4][84] ) );
  EDFFXL \block_reg[4][83]  ( .D(block_next[83]), .E(n1162), .CK(clk), .Q(
        \block[4][83] ) );
  EDFFXL \block_reg[4][82]  ( .D(block_next[82]), .E(n1162), .CK(clk), .Q(
        \block[4][82] ) );
  EDFFXL \block_reg[4][81]  ( .D(block_next[81]), .E(n1162), .CK(clk), .Q(
        \block[4][81] ) );
  EDFFXL \block_reg[4][80]  ( .D(block_next[80]), .E(n1162), .CK(clk), .Q(
        \block[4][80] ) );
  EDFFXL \block_reg[4][57]  ( .D(block_next[57]), .E(n1160), .CK(clk), .Q(
        \block[4][57] ) );
  EDFFXL \block_reg[4][25]  ( .D(block_next[25]), .E(n1157), .CK(clk), .Q(
        \block[4][25] ) );
  EDFFXL \block_reg[4][24]  ( .D(block_next[24]), .E(n1157), .CK(clk), .Q(
        \block[4][24] ) );
  EDFFXL \block_reg[4][23]  ( .D(block_next[23]), .E(n1157), .CK(clk), .Q(
        \block[4][23] ) );
  EDFFXL \block_reg[4][22]  ( .D(block_next[22]), .E(n1157), .CK(clk), .Q(
        \block[4][22] ) );
  EDFFXL \block_reg[4][21]  ( .D(block_next[21]), .E(n1157), .CK(clk), .Q(
        \block[4][21] ) );
  EDFFXL \block_reg[4][18]  ( .D(block_next[18]), .E(n1157), .CK(clk), .Q(
        \block[4][18] ) );
  EDFFXL \block_reg[4][16]  ( .D(block_next[16]), .E(n1157), .CK(clk), .Q(
        \block[4][16] ) );
  EDFFXL \block_reg[4][121]  ( .D(block_next[121]), .E(n1165), .CK(clk), .Q(
        \block[4][121] ) );
  EDFFXL \block_reg[4][120]  ( .D(block_next[120]), .E(n1165), .CK(clk), .Q(
        \block[4][120] ) );
  EDFFXL \block_reg[4][119]  ( .D(block_next[119]), .E(n1165), .CK(clk), .Q(
        \block[4][119] ) );
  EDFFXL \block_reg[4][118]  ( .D(block_next[118]), .E(n1165), .CK(clk), .Q(
        \block[4][118] ) );
  EDFFXL \block_reg[4][117]  ( .D(block_next[117]), .E(n1164), .CK(clk), .Q(
        \block[4][117] ) );
  EDFFXL \block_reg[4][48]  ( .D(block_next[48]), .E(n1159), .CK(clk), .Q(
        \block[4][48] ) );
  EDFFXL \block_reg[4][115]  ( .D(block_next[115]), .E(n1164), .CK(clk), .Q(
        \block[4][115] ) );
  EDFFXL \block_reg[4][114]  ( .D(block_next[114]), .E(n1164), .CK(clk), .Q(
        \block[4][114] ) );
  EDFFXL \block_reg[4][113]  ( .D(block_next[113]), .E(n1164), .CK(clk), .Q(
        \block[4][113] ) );
  EDFFXL \block_reg[4][17]  ( .D(block_next[17]), .E(n1157), .CK(clk), .Q(
        \block[4][17] ) );
  EDFFXL \block_reg[0][116]  ( .D(block_next[116]), .E(n1240), .CK(clk), .Q(
        \block[0][116] ) );
  EDFFXL \block_reg[0][112]  ( .D(block_next[112]), .E(n1240), .CK(clk), .Q(
        \block[0][112] ) );
  EDFFXL \block_reg[0][89]  ( .D(block_next[89]), .E(n1238), .CK(clk), .Q(
        \block[0][89] ) );
  EDFFXL \block_reg[0][88]  ( .D(block_next[88]), .E(n1238), .CK(clk), .Q(
        \block[0][88] ) );
  EDFFXL \block_reg[0][87]  ( .D(block_next[87]), .E(n1238), .CK(clk), .Q(
        \block[0][87] ) );
  EDFFXL \block_reg[0][86]  ( .D(block_next[86]), .E(n1238), .CK(clk), .Q(
        \block[0][86] ) );
  EDFFXL \block_reg[0][85]  ( .D(block_next[85]), .E(n1238), .CK(clk), .Q(
        \block[0][85] ) );
  EDFFXL \block_reg[0][84]  ( .D(block_next[84]), .E(n1238), .CK(clk), .Q(
        \block[0][84] ) );
  EDFFXL \block_reg[0][83]  ( .D(block_next[83]), .E(n1238), .CK(clk), .Q(
        \block[0][83] ) );
  EDFFXL \block_reg[0][82]  ( .D(block_next[82]), .E(n1238), .CK(clk), .Q(
        \block[0][82] ) );
  EDFFXL \block_reg[0][81]  ( .D(block_next[81]), .E(n1238), .CK(clk), .Q(
        \block[0][81] ) );
  EDFFXL \block_reg[0][80]  ( .D(block_next[80]), .E(n1238), .CK(clk), .Q(
        \block[0][80] ) );
  EDFFXL \block_reg[0][57]  ( .D(block_next[57]), .E(n1236), .CK(clk), .Q(
        \block[0][57] ) );
  EDFFXL \block_reg[0][25]  ( .D(block_next[25]), .E(n1233), .CK(clk), .Q(
        \block[0][25] ) );
  EDFFXL \block_reg[0][24]  ( .D(block_next[24]), .E(n1233), .CK(clk), .Q(
        \block[0][24] ) );
  EDFFXL \block_reg[0][23]  ( .D(block_next[23]), .E(n1233), .CK(clk), .Q(
        \block[0][23] ) );
  EDFFXL \block_reg[0][22]  ( .D(block_next[22]), .E(n1233), .CK(clk), .Q(
        \block[0][22] ) );
  EDFFXL \block_reg[0][21]  ( .D(block_next[21]), .E(n1233), .CK(clk), .Q(
        \block[0][21] ) );
  EDFFXL \block_reg[0][18]  ( .D(block_next[18]), .E(n1233), .CK(clk), .Q(
        \block[0][18] ) );
  EDFFXL \block_reg[0][16]  ( .D(block_next[16]), .E(n1233), .CK(clk), .Q(
        \block[0][16] ) );
  EDFFXL \block_reg[0][121]  ( .D(block_next[121]), .E(n1241), .CK(clk), .Q(
        \block[0][121] ) );
  EDFFXL \block_reg[0][120]  ( .D(block_next[120]), .E(n1241), .CK(clk), .Q(
        \block[0][120] ) );
  EDFFXL \block_reg[0][119]  ( .D(block_next[119]), .E(n1241), .CK(clk), .Q(
        \block[0][119] ) );
  EDFFXL \block_reg[0][118]  ( .D(block_next[118]), .E(n1241), .CK(clk), .Q(
        \block[0][118] ) );
  EDFFXL \block_reg[0][117]  ( .D(block_next[117]), .E(n1240), .CK(clk), .Q(
        \block[0][117] ) );
  EDFFXL \block_reg[0][48]  ( .D(block_next[48]), .E(n1235), .CK(clk), .Q(
        \block[0][48] ) );
  EDFFXL \block_reg[4][20]  ( .D(block_next[20]), .E(n1157), .CK(clk), .Q(
        \block[4][20] ) );
  EDFFXL \block_reg[4][19]  ( .D(block_next[19]), .E(n1157), .CK(clk), .Q(
        \block[4][19] ) );
  EDFFXL \block_reg[4][50]  ( .D(block_next[50]), .E(n1159), .CK(clk), .Q(
        \block[4][50] ) );
  EDFFXL \block_reg[4][49]  ( .D(block_next[49]), .E(n1159), .CK(clk), .Q(
        \block[4][49] ) );
  EDFFXL \block_reg[4][56]  ( .D(block_next[56]), .E(n1160), .CK(clk), .Q(
        \block[4][56] ) );
  EDFFXL \block_reg[4][55]  ( .D(block_next[55]), .E(n1160), .CK(clk), .Q(
        \block[4][55] ) );
  EDFFXL \block_reg[4][54]  ( .D(block_next[54]), .E(n1160), .CK(clk), .Q(
        \block[4][54] ) );
  EDFFXL \block_reg[4][53]  ( .D(block_next[53]), .E(n1160), .CK(clk), .Q(
        \block[4][53] ) );
  EDFFXL \block_reg[4][52]  ( .D(block_next[52]), .E(n1159), .CK(clk), .Q(
        \block[4][52] ) );
  EDFFXL \block_reg[4][51]  ( .D(block_next[51]), .E(n1159), .CK(clk), .Q(
        \block[4][51] ) );
  EDFFXL \block_reg[0][115]  ( .D(block_next[115]), .E(n1240), .CK(clk), .Q(
        \block[0][115] ) );
  EDFFXL \block_reg[0][114]  ( .D(block_next[114]), .E(n1240), .CK(clk), .Q(
        \block[0][114] ) );
  EDFFXL \block_reg[0][113]  ( .D(block_next[113]), .E(n1240), .CK(clk), .Q(
        \block[0][113] ) );
  EDFFXL \block_reg[0][17]  ( .D(block_next[17]), .E(n1233), .CK(clk), .Q(
        \block[0][17] ) );
  EDFFXL \block_reg[0][20]  ( .D(block_next[20]), .E(n1233), .CK(clk), .Q(
        \block[0][20] ) );
  EDFFXL \block_reg[0][19]  ( .D(block_next[19]), .E(n1233), .CK(clk), .Q(
        \block[0][19] ) );
  EDFFXL \block_reg[0][50]  ( .D(block_next[50]), .E(n1235), .CK(clk), .Q(
        \block[0][50] ) );
  EDFFXL \block_reg[0][49]  ( .D(block_next[49]), .E(n1235), .CK(clk), .Q(
        \block[0][49] ) );
  EDFFXL \block_reg[0][56]  ( .D(block_next[56]), .E(n1236), .CK(clk), .Q(
        \block[0][56] ) );
  EDFFXL \block_reg[0][55]  ( .D(block_next[55]), .E(n1236), .CK(clk), .Q(
        \block[0][55] ) );
  EDFFXL \block_reg[0][54]  ( .D(block_next[54]), .E(n1236), .CK(clk), .Q(
        \block[0][54] ) );
  EDFFXL \block_reg[0][53]  ( .D(block_next[53]), .E(n1236), .CK(clk), .Q(
        \block[0][53] ) );
  EDFFXL \block_reg[0][52]  ( .D(block_next[52]), .E(n1235), .CK(clk), .Q(
        \block[0][52] ) );
  EDFFXL \block_reg[0][51]  ( .D(block_next[51]), .E(n1235), .CK(clk), .Q(
        \block[0][51] ) );
  EDFFXL \block_reg[0][15]  ( .D(block_next[15]), .E(n1233), .CK(clk), .Q(
        \block[0][15] ) );
  EDFFXL \block_reg[4][15]  ( .D(block_next[15]), .E(n1157), .CK(clk), .Q(
        \block[4][15] ) );
  EDFFXL \block_reg[0][11]  ( .D(block_next[11]), .E(n1232), .CK(clk), .QN(
        n513) );
  EDFFXL \block_reg[4][11]  ( .D(block_next[11]), .E(n1156), .CK(clk), .QN(
        n517) );
  EDFFXL \block_reg[0][14]  ( .D(block_next[14]), .E(n1233), .CK(clk), .Q(
        \block[0][14] ) );
  EDFFXL \block_reg[4][14]  ( .D(block_next[14]), .E(n1157), .CK(clk), .Q(
        \block[4][14] ) );
  EDFFXL \block_reg[0][111]  ( .D(block_next[111]), .E(n1240), .CK(clk), .Q(
        \block[0][111] ) );
  EDFFXL \block_reg[4][111]  ( .D(block_next[111]), .E(n1164), .CK(clk), .Q(
        \block[4][111] ) );
  EDFFXL \block_reg[0][79]  ( .D(block_next[79]), .E(n1238), .CK(clk), .QN(
        n453) );
  EDFFXL \block_reg[0][107]  ( .D(block_next[107]), .E(n1240), .CK(clk), .QN(
        n381) );
  EDFFXL \block_reg[4][79]  ( .D(block_next[79]), .E(n1162), .CK(clk), .QN(
        n457) );
  EDFFXL \block_reg[4][107]  ( .D(block_next[107]), .E(n1164), .CK(clk), .QN(
        n385) );
  EDFFXL \block_reg[0][109]  ( .D(block_next[109]), .E(n1240), .CK(clk), .QN(
        n461) );
  EDFFXL \block_reg[0][110]  ( .D(block_next[110]), .E(n1240), .CK(clk), .QN(
        n429) );
  EDFFXL \block_reg[4][109]  ( .D(block_next[109]), .E(n1164), .CK(clk), .QN(
        n465) );
  EDFFXL \block_reg[4][110]  ( .D(block_next[110]), .E(n1164), .CK(clk), .QN(
        n433) );
  EDFFXL \block_reg[0][75]  ( .D(block_next[75]), .E(n1237), .CK(clk), .QN(
        n333) );
  EDFFXL \block_reg[0][13]  ( .D(block_next[13]), .E(n1232), .CK(clk), .QN(
        n537) );
  EDFFXL \block_reg[4][75]  ( .D(block_next[75]), .E(n1161), .CK(clk), .QN(
        n337) );
  EDFFXL \block_reg[4][13]  ( .D(block_next[13]), .E(n1156), .CK(clk), .QN(
        n541) );
  EDFFXL \block_reg[0][78]  ( .D(block_next[78]), .E(n1237), .CK(clk), .QN(
        n413) );
  EDFFXL \block_reg[0][12]  ( .D(block_next[12]), .E(n1232), .CK(clk), .QN(
        n529) );
  EDFFXL \block_reg[4][78]  ( .D(block_next[78]), .E(n1161), .CK(clk), .QN(
        n417) );
  EDFFXL \block_reg[4][12]  ( .D(block_next[12]), .E(n1156), .CK(clk), .QN(
        n533) );
  EDFFXL \block_reg[0][8]  ( .D(block_next[8]), .E(n1232), .CK(clk), .Q(
        \block[0][8] ) );
  EDFFXL \block_reg[0][10]  ( .D(block_next[10]), .E(n1232), .CK(clk), .QN(
        n505) );
  EDFFXL \block_reg[4][8]  ( .D(block_next[8]), .E(n1156), .CK(clk), .Q(
        \block[4][8] ) );
  EDFFXL \block_reg[0][47]  ( .D(block_next[47]), .E(n1235), .CK(clk), .QN(
        n545) );
  EDFFXL \block_reg[4][10]  ( .D(block_next[10]), .E(n1156), .CK(clk), .QN(
        n509) );
  EDFFXL \block_reg[4][47]  ( .D(block_next[47]), .E(n1159), .CK(clk), .QN(
        n549) );
  EDFFXL \block_reg[0][108]  ( .D(block_next[108]), .E(n1240), .CK(clk), .QN(
        n397) );
  EDFFXL \block_reg[0][43]  ( .D(block_next[43]), .E(n1235), .CK(clk), .QN(
        n349) );
  EDFFXL \block_reg[0][44]  ( .D(block_next[44]), .E(n1235), .CK(clk), .QN(
        n365) );
  EDFFXL \block_reg[4][44]  ( .D(block_next[44]), .E(n1159), .CK(clk), .QN(
        n369) );
  EDFFXL \block_reg[4][108]  ( .D(block_next[108]), .E(n1164), .CK(clk), .QN(
        n401) );
  EDFFXL \block_reg[4][43]  ( .D(block_next[43]), .E(n1159), .CK(clk), .QN(
        n353) );
  EDFFXL \block_reg[0][106]  ( .D(block_next[106]), .E(n1240), .CK(clk), .QN(
        n373) );
  EDFFXL \block_reg[4][106]  ( .D(block_next[106]), .E(n1164), .CK(clk), .QN(
        n377) );
  EDFFXL \block_reg[0][46]  ( .D(block_next[46]), .E(n1235), .CK(clk), .Q(
        \block[0][46] ) );
  EDFFXL \block_reg[0][77]  ( .D(block_next[77]), .E(n1237), .CK(clk), .QN(
        n421) );
  EDFFXL \block_reg[0][76]  ( .D(block_next[76]), .E(n1237), .CK(clk), .QN(
        n445) );
  EDFFXL \block_reg[4][77]  ( .D(block_next[77]), .E(n1161), .CK(clk), .QN(
        n425) );
  EDFFXL \block_reg[4][46]  ( .D(block_next[46]), .E(n1159), .CK(clk), .Q(
        \block[4][46] ) );
  EDFFXL \block_reg[0][104]  ( .D(block_next[104]), .E(n1239), .CK(clk), .Q(
        \block[0][104] ) );
  EDFFXL \block_reg[4][76]  ( .D(block_next[76]), .E(n1161), .CK(clk), .QN(
        n449) );
  EDFFXL \block_reg[4][104]  ( .D(block_next[104]), .E(n1163), .CK(clk), .Q(
        \block[4][104] ) );
  EDFFXL \block_reg[0][74]  ( .D(block_next[74]), .E(n1237), .CK(clk), .QN(
        n325) );
  EDFFXL \block_reg[4][74]  ( .D(block_next[74]), .E(n1161), .CK(clk), .QN(
        n329) );
  EDFFXL \block_reg[0][9]  ( .D(block_next[9]), .E(n1232), .CK(clk), .QN(n521)
         );
  EDFFXL \block_reg[4][9]  ( .D(block_next[9]), .E(n1156), .CK(clk), .QN(n525)
         );
  EDFFXL \block_reg[0][45]  ( .D(block_next[45]), .E(n1235), .CK(clk), .QN(
        n405) );
  EDFFXL \block_reg[4][45]  ( .D(block_next[45]), .E(n1159), .CK(clk), .QN(
        n409) );
  EDFFXL \block_reg[0][42]  ( .D(block_next[42]), .E(n1235), .CK(clk), .QN(
        n437) );
  EDFFXL \block_reg[0][105]  ( .D(block_next[105]), .E(n1240), .CK(clk), .QN(
        n389) );
  EDFFXL \block_reg[4][42]  ( .D(block_next[42]), .E(n1159), .CK(clk), .QN(
        n441) );
  EDFFXL \block_reg[4][105]  ( .D(block_next[105]), .E(n1164), .CK(clk), .QN(
        n393) );
  EDFFXL \block_reg[0][73]  ( .D(block_next[73]), .E(n1237), .CK(clk), .QN(
        n341) );
  EDFFXL \block_reg[4][73]  ( .D(block_next[73]), .E(n1161), .CK(clk), .QN(
        n345) );
  EDFFXL \block_reg[0][72]  ( .D(block_next[72]), .E(n1237), .CK(clk), .Q(
        \block[0][72] ) );
  EDFFXL \block_reg[4][72]  ( .D(block_next[72]), .E(n1161), .CK(clk), .Q(
        \block[4][72] ) );
  EDFFXL \block_reg[0][41]  ( .D(block_next[41]), .E(n1235), .CK(clk), .QN(
        n357) );
  EDFFXL \block_reg[4][41]  ( .D(block_next[41]), .E(n1159), .CK(clk), .QN(
        n361) );
  EDFFXL \block_reg[0][40]  ( .D(block_next[40]), .E(n1235), .CK(clk), .Q(
        \block[0][40] ) );
  EDFFXL \block_reg[4][40]  ( .D(block_next[40]), .E(n1159), .CK(clk), .Q(
        \block[4][40] ) );
  EDFFXL \block_reg[0][6]  ( .D(block_next[6]), .E(n1232), .CK(clk), .Q(
        \block[0][6] ) );
  EDFFXL \block_reg[4][6]  ( .D(block_next[6]), .E(n1156), .CK(clk), .Q(
        \block[4][6] ) );
  EDFFXL \block_reg[0][102]  ( .D(block_next[102]), .E(n1239), .CK(clk), .Q(
        \block[0][102] ) );
  EDFFXL \block_reg[4][102]  ( .D(block_next[102]), .E(n1163), .CK(clk), .Q(
        \block[4][102] ) );
  EDFFXL \block_reg[0][70]  ( .D(block_next[70]), .E(n1237), .CK(clk), .Q(
        \block[0][70] ) );
  EDFFXL \block_reg[4][70]  ( .D(block_next[70]), .E(n1161), .CK(clk), .Q(
        \block[4][70] ) );
  EDFFXL \block_reg[0][38]  ( .D(block_next[38]), .E(n1234), .CK(clk), .Q(
        \block[0][38] ) );
  EDFFXL \block_reg[4][38]  ( .D(block_next[38]), .E(n1158), .CK(clk), .Q(
        \block[4][38] ) );
  EDFFXL \block_reg[0][0]  ( .D(block_next[0]), .E(n1231), .CK(clk), .Q(
        \block[0][0] ) );
  EDFFXL \block_reg[4][0]  ( .D(block_next[0]), .E(n1155), .CK(clk), .Q(
        \block[4][0] ) );
  EDFFXL \block_reg[0][96]  ( .D(block_next[96]), .E(n1239), .CK(clk), .Q(
        \block[0][96] ) );
  EDFFXL \block_reg[4][96]  ( .D(block_next[96]), .E(n1163), .CK(clk), .Q(
        \block[4][96] ) );
  EDFFXL \block_reg[0][64]  ( .D(block_next[64]), .E(n1236), .CK(clk), .Q(
        \block[0][64] ) );
  EDFFXL \block_reg[4][64]  ( .D(block_next[64]), .E(n1160), .CK(clk), .Q(
        \block[4][64] ) );
  EDFFXL \block_reg[0][32]  ( .D(block_next[32]), .E(n1234), .CK(clk), .Q(
        \block[0][32] ) );
  EDFFXL \block_reg[4][32]  ( .D(block_next[32]), .E(n1158), .CK(clk), .Q(
        \block[4][32] ) );
  EDFFXL \block_reg[0][5]  ( .D(block_next[5]), .E(n1232), .CK(clk), .QN(n309)
         );
  EDFFXL \block_reg[4][5]  ( .D(block_next[5]), .E(n1156), .CK(clk), .QN(n313)
         );
  EDFFXL \block_reg[0][7]  ( .D(block_next[7]), .E(n1232), .CK(clk), .Q(
        \block[0][7] ) );
  EDFFXL \block_reg[4][7]  ( .D(block_next[7]), .E(n1156), .CK(clk), .Q(
        \block[4][7] ) );
  EDFFXL \block_reg[0][3]  ( .D(block_next[3]), .E(n1232), .CK(clk), .Q(
        \block[0][3] ) );
  EDFFXL \block_reg[0][4]  ( .D(block_next[4]), .E(n1232), .CK(clk), .Q(
        \block[0][4] ) );
  EDFFXL \block_reg[4][3]  ( .D(block_next[3]), .E(n1156), .CK(clk), .Q(
        \block[4][3] ) );
  EDFFXL \block_reg[0][1]  ( .D(block_next[1]), .E(n1232), .CK(clk), .Q(
        \block[0][1] ) );
  EDFFXL \block_reg[4][4]  ( .D(block_next[4]), .E(n1156), .CK(clk), .Q(
        \block[4][4] ) );
  EDFFXL \block_reg[4][1]  ( .D(block_next[1]), .E(n1156), .CK(clk), .Q(
        \block[4][1] ) );
  EDFFXL \block_reg[0][2]  ( .D(block_next[2]), .E(n1232), .CK(clk), .Q(
        \block[0][2] ) );
  EDFFXL \block_reg[4][2]  ( .D(block_next[2]), .E(n1156), .CK(clk), .Q(
        \block[4][2] ) );
  EDFFXL \block_reg[0][103]  ( .D(block_next[103]), .E(n1239), .CK(clk), .Q(
        \block[0][103] ) );
  EDFFXL \block_reg[4][103]  ( .D(block_next[103]), .E(n1163), .CK(clk), .Q(
        \block[4][103] ) );
  EDFFXL \block_reg[0][101]  ( .D(block_next[101]), .E(n1239), .CK(clk), .Q(
        \block[0][101] ) );
  EDFFXL \block_reg[4][101]  ( .D(block_next[101]), .E(n1163), .CK(clk), .Q(
        \block[4][101] ) );
  EDFFXL \block_reg[0][71]  ( .D(block_next[71]), .E(n1237), .CK(clk), .Q(
        \block[0][71] ) );
  EDFFXL \block_reg[4][71]  ( .D(block_next[71]), .E(n1161), .CK(clk), .Q(
        \block[4][71] ) );
  EDFFXL \block_reg[0][68]  ( .D(block_next[68]), .E(n1237), .CK(clk), .Q(
        \block[0][68] ) );
  EDFFXL \block_reg[4][68]  ( .D(block_next[68]), .E(n1161), .CK(clk), .Q(
        \block[4][68] ) );
  EDFFXL \block_reg[0][67]  ( .D(block_next[67]), .E(n1237), .CK(clk), .Q(
        \block[0][67] ) );
  EDFFXL \block_reg[0][37]  ( .D(block_next[37]), .E(n1234), .CK(clk), .Q(
        \block[0][37] ) );
  EDFFXL \block_reg[4][37]  ( .D(block_next[37]), .E(n1158), .CK(clk), .Q(
        \block[4][37] ) );
  EDFFXL \block_reg[4][67]  ( .D(block_next[67]), .E(n1161), .CK(clk), .Q(
        \block[4][67] ) );
  EDFFXL \block_reg[0][39]  ( .D(block_next[39]), .E(n1234), .CK(clk), .Q(
        \block[0][39] ) );
  EDFFXL \block_reg[4][39]  ( .D(block_next[39]), .E(n1158), .CK(clk), .Q(
        \block[4][39] ) );
  EDFFXL \block_reg[0][69]  ( .D(block_next[69]), .E(n1237), .CK(clk), .Q(
        \block[0][69] ) );
  EDFFXL \block_reg[0][100]  ( .D(block_next[100]), .E(n1239), .CK(clk), .Q(
        \block[0][100] ) );
  EDFFXL \block_reg[4][69]  ( .D(block_next[69]), .E(n1161), .CK(clk), .Q(
        \block[4][69] ) );
  EDFFXL \block_reg[4][100]  ( .D(block_next[100]), .E(n1163), .CK(clk), .Q(
        \block[4][100] ) );
  EDFFXL \block_reg[0][99]  ( .D(block_next[99]), .E(n1239), .CK(clk), .Q(
        \block[0][99] ) );
  EDFFXL \block_reg[0][97]  ( .D(block_next[97]), .E(n1239), .CK(clk), .Q(
        \block[0][97] ) );
  EDFFXL \block_reg[4][99]  ( .D(block_next[99]), .E(n1163), .CK(clk), .Q(
        \block[4][99] ) );
  EDFFXL \block_reg[4][97]  ( .D(block_next[97]), .E(n1163), .CK(clk), .Q(
        \block[4][97] ) );
  EDFFXL \block_reg[0][65]  ( .D(block_next[65]), .E(n1236), .CK(clk), .Q(
        \block[0][65] ) );
  EDFFXL \block_reg[4][65]  ( .D(block_next[65]), .E(n1160), .CK(clk), .Q(
        \block[4][65] ) );
  EDFFXL \block_reg[0][36]  ( .D(block_next[36]), .E(n1234), .CK(clk), .QN(
        n317) );
  EDFFXL \block_reg[0][98]  ( .D(block_next[98]), .E(n1239), .CK(clk), .Q(
        \block[0][98] ) );
  EDFFXL \block_reg[4][36]  ( .D(block_next[36]), .E(n1158), .CK(clk), .QN(
        n321) );
  EDFFXL \block_reg[4][98]  ( .D(block_next[98]), .E(n1163), .CK(clk), .Q(
        \block[4][98] ) );
  EDFFXL \block_reg[0][66]  ( .D(block_next[66]), .E(n1237), .CK(clk), .Q(
        \block[0][66] ) );
  EDFFXL \block_reg[4][66]  ( .D(block_next[66]), .E(n1161), .CK(clk), .Q(
        \block[4][66] ) );
  EDFFXL \block_reg[0][35]  ( .D(block_next[35]), .E(n1234), .CK(clk), .Q(
        \block[0][35] ) );
  EDFFXL \block_reg[4][35]  ( .D(block_next[35]), .E(n1158), .CK(clk), .Q(
        \block[4][35] ) );
  EDFFXL \block_reg[0][33]  ( .D(block_next[33]), .E(n1234), .CK(clk), .Q(
        \block[0][33] ) );
  EDFFXL \block_reg[4][33]  ( .D(block_next[33]), .E(n1158), .CK(clk), .Q(
        \block[4][33] ) );
  EDFFXL \block_reg[0][34]  ( .D(block_next[34]), .E(n1234), .CK(clk), .Q(
        \block[0][34] ) );
  EDFFXL \block_reg[4][34]  ( .D(block_next[34]), .E(n1158), .CK(clk), .Q(
        \block[4][34] ) );
  EDFFXL \block_reg[0][122]  ( .D(block_next[122]), .E(n1241), .CK(clk), .Q(
        \block[0][122] ) );
  EDFFXL \block_reg[4][122]  ( .D(block_next[122]), .E(n1165), .CK(clk), .Q(
        \block[4][122] ) );
  EDFFXL \block_reg[0][26]  ( .D(block_next[26]), .E(n1233), .CK(clk), .QN(
        n291) );
  EDFFXL \block_reg[4][26]  ( .D(block_next[26]), .E(n1157), .CK(clk), .QN(
        n295) );
  EDFFXL \block_reg[6][116]  ( .D(block_next[116]), .E(n1125), .CK(clk), .Q(
        \block[6][116] ) );
  EDFFXL \block_reg[6][112]  ( .D(block_next[112]), .E(n1125), .CK(clk), .Q(
        \block[6][112] ) );
  EDFFXL \block_reg[6][89]  ( .D(block_next[89]), .E(n1123), .CK(clk), .Q(
        \block[6][89] ) );
  EDFFXL \block_reg[6][88]  ( .D(block_next[88]), .E(n1123), .CK(clk), .Q(
        \block[6][88] ) );
  EDFFXL \block_reg[6][87]  ( .D(block_next[87]), .E(n1123), .CK(clk), .Q(
        \block[6][87] ) );
  EDFFXL \block_reg[6][86]  ( .D(block_next[86]), .E(n1123), .CK(clk), .Q(
        \block[6][86] ) );
  EDFFXL \block_reg[6][85]  ( .D(block_next[85]), .E(n1123), .CK(clk), .Q(
        \block[6][85] ) );
  EDFFXL \block_reg[6][84]  ( .D(block_next[84]), .E(n1123), .CK(clk), .Q(
        \block[6][84] ) );
  EDFFXL \block_reg[6][83]  ( .D(block_next[83]), .E(n1123), .CK(clk), .Q(
        \block[6][83] ) );
  EDFFXL \block_reg[6][82]  ( .D(block_next[82]), .E(n1123), .CK(clk), .Q(
        \block[6][82] ) );
  EDFFXL \block_reg[6][81]  ( .D(block_next[81]), .E(n1123), .CK(clk), .Q(
        \block[6][81] ) );
  EDFFXL \block_reg[6][80]  ( .D(block_next[80]), .E(n1123), .CK(clk), .Q(
        \block[6][80] ) );
  EDFFXL \block_reg[6][57]  ( .D(block_next[57]), .E(n1121), .CK(clk), .Q(
        \block[6][57] ) );
  EDFFXL \block_reg[6][25]  ( .D(block_next[25]), .E(n1118), .CK(clk), .Q(
        \block[6][25] ) );
  EDFFXL \block_reg[6][24]  ( .D(block_next[24]), .E(n1118), .CK(clk), .Q(
        \block[6][24] ) );
  EDFFXL \block_reg[6][23]  ( .D(block_next[23]), .E(n1118), .CK(clk), .Q(
        \block[6][23] ) );
  EDFFXL \block_reg[6][22]  ( .D(block_next[22]), .E(n1118), .CK(clk), .Q(
        \block[6][22] ) );
  EDFFXL \block_reg[6][21]  ( .D(block_next[21]), .E(n1118), .CK(clk), .Q(
        \block[6][21] ) );
  EDFFXL \block_reg[6][18]  ( .D(block_next[18]), .E(n1118), .CK(clk), .Q(
        \block[6][18] ) );
  EDFFXL \block_reg[6][16]  ( .D(block_next[16]), .E(n1118), .CK(clk), .Q(
        \block[6][16] ) );
  EDFFXL \block_reg[6][121]  ( .D(block_next[121]), .E(n1126), .CK(clk), .Q(
        \block[6][121] ) );
  EDFFXL \block_reg[6][120]  ( .D(block_next[120]), .E(n1126), .CK(clk), .Q(
        \block[6][120] ) );
  EDFFXL \block_reg[6][119]  ( .D(block_next[119]), .E(n1126), .CK(clk), .Q(
        \block[6][119] ) );
  EDFFXL \block_reg[6][118]  ( .D(block_next[118]), .E(n1126), .CK(clk), .Q(
        \block[6][118] ) );
  EDFFXL \block_reg[6][117]  ( .D(block_next[117]), .E(n1125), .CK(clk), .Q(
        \block[6][117] ) );
  EDFFXL \block_reg[6][48]  ( .D(block_next[48]), .E(n1120), .CK(clk), .Q(
        \block[6][48] ) );
  EDFFXL \block_reg[6][115]  ( .D(block_next[115]), .E(n1125), .CK(clk), .Q(
        \block[6][115] ) );
  EDFFXL \block_reg[6][114]  ( .D(block_next[114]), .E(n1125), .CK(clk), .Q(
        \block[6][114] ) );
  EDFFXL \block_reg[6][113]  ( .D(block_next[113]), .E(n1125), .CK(clk), .Q(
        \block[6][113] ) );
  EDFFXL \block_reg[6][17]  ( .D(block_next[17]), .E(n1118), .CK(clk), .Q(
        \block[6][17] ) );
  EDFFXL \block_reg[6][20]  ( .D(block_next[20]), .E(n1118), .CK(clk), .Q(
        \block[6][20] ) );
  EDFFXL \block_reg[6][19]  ( .D(block_next[19]), .E(n1118), .CK(clk), .Q(
        \block[6][19] ) );
  EDFFXL \block_reg[6][50]  ( .D(block_next[50]), .E(n1120), .CK(clk), .Q(
        \block[6][50] ) );
  EDFFXL \block_reg[6][49]  ( .D(block_next[49]), .E(n1120), .CK(clk), .Q(
        \block[6][49] ) );
  EDFFXL \block_reg[2][116]  ( .D(block_next[116]), .E(n1202), .CK(clk), .Q(
        \block[2][116] ) );
  EDFFXL \block_reg[2][112]  ( .D(block_next[112]), .E(n1202), .CK(clk), .Q(
        \block[2][112] ) );
  EDFFXL \block_reg[2][89]  ( .D(block_next[89]), .E(n1200), .CK(clk), .Q(
        \block[2][89] ) );
  EDFFXL \block_reg[2][88]  ( .D(block_next[88]), .E(n1200), .CK(clk), .Q(
        \block[2][88] ) );
  EDFFXL \block_reg[2][87]  ( .D(block_next[87]), .E(n1200), .CK(clk), .Q(
        \block[2][87] ) );
  EDFFXL \block_reg[2][86]  ( .D(block_next[86]), .E(n1200), .CK(clk), .Q(
        \block[2][86] ) );
  EDFFXL \block_reg[2][85]  ( .D(block_next[85]), .E(n1200), .CK(clk), .Q(
        \block[2][85] ) );
  EDFFXL \block_reg[2][84]  ( .D(block_next[84]), .E(n1200), .CK(clk), .Q(
        \block[2][84] ) );
  EDFFXL \block_reg[2][83]  ( .D(block_next[83]), .E(n1200), .CK(clk), .Q(
        \block[2][83] ) );
  EDFFXL \block_reg[2][82]  ( .D(block_next[82]), .E(n1200), .CK(clk), .Q(
        \block[2][82] ) );
  EDFFXL \block_reg[2][81]  ( .D(block_next[81]), .E(n1200), .CK(clk), .Q(
        \block[2][81] ) );
  EDFFXL \block_reg[2][80]  ( .D(block_next[80]), .E(n1200), .CK(clk), .Q(
        \block[2][80] ) );
  EDFFXL \block_reg[2][57]  ( .D(block_next[57]), .E(n1198), .CK(clk), .Q(
        \block[2][57] ) );
  EDFFXL \block_reg[2][25]  ( .D(block_next[25]), .E(n1195), .CK(clk), .Q(
        \block[2][25] ) );
  EDFFXL \block_reg[2][24]  ( .D(block_next[24]), .E(n1195), .CK(clk), .Q(
        \block[2][24] ) );
  EDFFXL \block_reg[2][23]  ( .D(block_next[23]), .E(n1195), .CK(clk), .Q(
        \block[2][23] ) );
  EDFFXL \block_reg[2][22]  ( .D(block_next[22]), .E(n1195), .CK(clk), .Q(
        \block[2][22] ) );
  EDFFXL \block_reg[2][21]  ( .D(block_next[21]), .E(n1195), .CK(clk), .Q(
        \block[2][21] ) );
  EDFFXL \block_reg[2][18]  ( .D(block_next[18]), .E(n1195), .CK(clk), .Q(
        \block[2][18] ) );
  EDFFXL \block_reg[2][16]  ( .D(block_next[16]), .E(n1195), .CK(clk), .Q(
        \block[2][16] ) );
  EDFFXL \block_reg[2][121]  ( .D(block_next[121]), .E(n1203), .CK(clk), .Q(
        \block[2][121] ) );
  EDFFXL \block_reg[2][120]  ( .D(block_next[120]), .E(n1203), .CK(clk), .Q(
        \block[2][120] ) );
  EDFFXL \block_reg[2][119]  ( .D(block_next[119]), .E(n1203), .CK(clk), .Q(
        \block[2][119] ) );
  EDFFXL \block_reg[2][118]  ( .D(block_next[118]), .E(n1203), .CK(clk), .Q(
        \block[2][118] ) );
  EDFFXL \block_reg[2][117]  ( .D(block_next[117]), .E(n1202), .CK(clk), .Q(
        \block[2][117] ) );
  EDFFXL \block_reg[6][56]  ( .D(block_next[56]), .E(n1121), .CK(clk), .Q(
        \block[6][56] ) );
  EDFFXL \block_reg[6][55]  ( .D(block_next[55]), .E(n1121), .CK(clk), .Q(
        \block[6][55] ) );
  EDFFXL \block_reg[6][54]  ( .D(block_next[54]), .E(n1121), .CK(clk), .Q(
        \block[6][54] ) );
  EDFFXL \block_reg[6][53]  ( .D(block_next[53]), .E(n1121), .CK(clk), .Q(
        \block[6][53] ) );
  EDFFXL \block_reg[6][52]  ( .D(block_next[52]), .E(n1120), .CK(clk), .Q(
        \block[6][52] ) );
  EDFFXL \block_reg[6][51]  ( .D(block_next[51]), .E(n1120), .CK(clk), .Q(
        \block[6][51] ) );
  EDFFXL \block_reg[2][48]  ( .D(block_next[48]), .E(n1197), .CK(clk), .Q(
        \block[2][48] ) );
  EDFFXL \block_reg[2][115]  ( .D(block_next[115]), .E(n1202), .CK(clk), .Q(
        \block[2][115] ) );
  EDFFXL \block_reg[2][114]  ( .D(block_next[114]), .E(n1202), .CK(clk), .Q(
        \block[2][114] ) );
  EDFFXL \block_reg[2][113]  ( .D(block_next[113]), .E(n1202), .CK(clk), .Q(
        \block[2][113] ) );
  EDFFXL \block_reg[2][17]  ( .D(block_next[17]), .E(n1195), .CK(clk), .Q(
        \block[2][17] ) );
  EDFFXL \block_reg[2][20]  ( .D(block_next[20]), .E(n1195), .CK(clk), .Q(
        \block[2][20] ) );
  EDFFXL \block_reg[2][19]  ( .D(block_next[19]), .E(n1195), .CK(clk), .Q(
        \block[2][19] ) );
  EDFFXL \block_reg[2][50]  ( .D(block_next[50]), .E(n1197), .CK(clk), .Q(
        \block[2][50] ) );
  EDFFXL \block_reg[2][49]  ( .D(block_next[49]), .E(n1197), .CK(clk), .Q(
        \block[2][49] ) );
  EDFFXL \block_reg[2][56]  ( .D(block_next[56]), .E(n1198), .CK(clk), .Q(
        \block[2][56] ) );
  EDFFXL \block_reg[2][55]  ( .D(block_next[55]), .E(n1198), .CK(clk), .Q(
        \block[2][55] ) );
  EDFFXL \block_reg[2][54]  ( .D(block_next[54]), .E(n1198), .CK(clk), .Q(
        \block[2][54] ) );
  EDFFXL \block_reg[2][53]  ( .D(block_next[53]), .E(n1198), .CK(clk), .Q(
        \block[2][53] ) );
  EDFFXL \block_reg[2][52]  ( .D(block_next[52]), .E(n1197), .CK(clk), .Q(
        \block[2][52] ) );
  EDFFXL \block_reg[2][51]  ( .D(block_next[51]), .E(n1197), .CK(clk), .Q(
        \block[2][51] ) );
  EDFFXL \block_reg[2][15]  ( .D(block_next[15]), .E(n1195), .CK(clk), .Q(
        \block[2][15] ) );
  EDFFXL \block_reg[6][15]  ( .D(block_next[15]), .E(n1118), .CK(clk), .Q(
        \block[6][15] ) );
  EDFFXL \block_reg[2][11]  ( .D(block_next[11]), .E(n1194), .CK(clk), .QN(
        n515) );
  EDFFXL \block_reg[6][11]  ( .D(block_next[11]), .E(n1117), .CK(clk), .QN(
        n519) );
  EDFFXL \block_reg[2][14]  ( .D(block_next[14]), .E(n1195), .CK(clk), .Q(
        \block[2][14] ) );
  EDFFXL \block_reg[6][14]  ( .D(block_next[14]), .E(n1118), .CK(clk), .Q(
        \block[6][14] ) );
  EDFFXL \block_reg[2][111]  ( .D(block_next[111]), .E(n1202), .CK(clk), .Q(
        \block[2][111] ) );
  EDFFXL \block_reg[6][111]  ( .D(block_next[111]), .E(n1125), .CK(clk), .Q(
        \block[6][111] ) );
  EDFFXL \block_reg[2][79]  ( .D(block_next[79]), .E(n1200), .CK(clk), .QN(
        n455) );
  EDFFXL \block_reg[2][107]  ( .D(block_next[107]), .E(n1202), .CK(clk), .QN(
        n383) );
  EDFFXL \block_reg[6][79]  ( .D(block_next[79]), .E(n1123), .CK(clk), .QN(
        n459) );
  EDFFXL \block_reg[6][107]  ( .D(block_next[107]), .E(n1125), .CK(clk), .QN(
        n387) );
  EDFFXL \block_reg[2][110]  ( .D(block_next[110]), .E(n1202), .CK(clk), .QN(
        n431) );
  EDFFXL \block_reg[2][109]  ( .D(block_next[109]), .E(n1202), .CK(clk), .QN(
        n463) );
  EDFFXL \block_reg[6][110]  ( .D(block_next[110]), .E(n1125), .CK(clk), .QN(
        n435) );
  EDFFXL \block_reg[6][109]  ( .D(block_next[109]), .E(n1125), .CK(clk), .QN(
        n502) );
  EDFFXL \block_reg[2][75]  ( .D(block_next[75]), .E(n1199), .CK(clk), .QN(
        n335) );
  EDFFXL \block_reg[2][13]  ( .D(block_next[13]), .E(n1194), .CK(clk), .QN(
        n539) );
  EDFFXL \block_reg[6][75]  ( .D(block_next[75]), .E(n1122), .CK(clk), .QN(
        n339) );
  EDFFXL \block_reg[6][13]  ( .D(block_next[13]), .E(n1117), .CK(clk), .QN(
        n543) );
  EDFFXL \block_reg[2][12]  ( .D(block_next[12]), .E(n1194), .CK(clk), .QN(
        n531) );
  EDFFXL \block_reg[2][78]  ( .D(block_next[78]), .E(n1199), .CK(clk), .QN(
        n415) );
  EDFFXL \block_reg[6][12]  ( .D(block_next[12]), .E(n1117), .CK(clk), .QN(
        n535) );
  EDFFXL \block_reg[6][78]  ( .D(block_next[78]), .E(n1122), .CK(clk), .QN(
        n419) );
  EDFFXL \block_reg[2][10]  ( .D(block_next[10]), .E(n1194), .CK(clk), .QN(
        n507) );
  EDFFXL \block_reg[2][47]  ( .D(block_next[47]), .E(n1197), .CK(clk), .QN(
        n547) );
  EDFFXL \block_reg[2][8]  ( .D(block_next[8]), .E(n1194), .CK(clk), .Q(
        \block[2][8] ) );
  EDFFXL \block_reg[6][8]  ( .D(block_next[8]), .E(n1117), .CK(clk), .Q(
        \block[6][8] ) );
  EDFFXL \block_reg[6][10]  ( .D(block_next[10]), .E(n1117), .CK(clk), .QN(
        n511) );
  EDFFXL \block_reg[6][47]  ( .D(block_next[47]), .E(n1120), .CK(clk), .QN(
        n551) );
  EDFFXL \block_reg[2][108]  ( .D(block_next[108]), .E(n1202), .CK(clk), .QN(
        n399) );
  EDFFXL \block_reg[2][43]  ( .D(block_next[43]), .E(n1197), .CK(clk), .QN(
        n351) );
  EDFFXL \block_reg[2][44]  ( .D(block_next[44]), .E(n1197), .CK(clk), .QN(
        n367) );
  EDFFXL \block_reg[6][108]  ( .D(block_next[108]), .E(n1125), .CK(clk), .QN(
        n403) );
  EDFFXL \block_reg[6][43]  ( .D(block_next[43]), .E(n1120), .CK(clk), .QN(
        n355) );
  EDFFXL \block_reg[6][44]  ( .D(block_next[44]), .E(n1120), .CK(clk), .QN(
        n371) );
  EDFFXL \block_reg[2][106]  ( .D(block_next[106]), .E(n1202), .CK(clk), .QN(
        n375) );
  EDFFXL \block_reg[6][106]  ( .D(block_next[106]), .E(n1125), .CK(clk), .QN(
        n379) );
  EDFFXL \block_reg[2][46]  ( .D(block_next[46]), .E(n1197), .CK(clk), .Q(
        \block[2][46] ) );
  EDFFXL \block_reg[2][77]  ( .D(block_next[77]), .E(n1199), .CK(clk), .QN(
        n423) );
  EDFFXL \block_reg[2][76]  ( .D(block_next[76]), .E(n1199), .CK(clk), .QN(
        n447) );
  EDFFXL \block_reg[6][46]  ( .D(block_next[46]), .E(n1120), .CK(clk), .Q(
        \block[6][46] ) );
  EDFFXL \block_reg[6][77]  ( .D(block_next[77]), .E(n1122), .CK(clk), .QN(
        n427) );
  EDFFXL \block_reg[6][76]  ( .D(block_next[76]), .E(n1122), .CK(clk), .QN(
        n451) );
  EDFFXL \block_reg[2][104]  ( .D(block_next[104]), .E(n1201), .CK(clk), .Q(
        \block[2][104] ) );
  EDFFXL \block_reg[2][74]  ( .D(block_next[74]), .E(n1199), .CK(clk), .QN(
        n327) );
  EDFFXL \block_reg[6][104]  ( .D(block_next[104]), .E(n1124), .CK(clk), .Q(
        \block[6][104] ) );
  EDFFXL \block_reg[6][74]  ( .D(block_next[74]), .E(n1122), .CK(clk), .QN(
        n331) );
  EDFFXL \block_reg[2][9]  ( .D(block_next[9]), .E(n1194), .CK(clk), .QN(n523)
         );
  EDFFXL \block_reg[6][9]  ( .D(block_next[9]), .E(n1117), .CK(clk), .QN(n527)
         );
  EDFFXL \block_reg[2][45]  ( .D(block_next[45]), .E(n1197), .CK(clk), .QN(
        n407) );
  EDFFXL \block_reg[6][45]  ( .D(block_next[45]), .E(n1120), .CK(clk), .QN(
        n411) );
  EDFFXL \block_reg[2][42]  ( .D(block_next[42]), .E(n1197), .CK(clk), .QN(
        n439) );
  EDFFXL \block_reg[2][105]  ( .D(block_next[105]), .E(n1202), .CK(clk), .QN(
        n391) );
  EDFFXL \block_reg[6][42]  ( .D(block_next[42]), .E(n1120), .CK(clk), .QN(
        n443) );
  EDFFXL \block_reg[6][105]  ( .D(block_next[105]), .E(n1125), .CK(clk), .QN(
        n395) );
  EDFFXL \block_reg[2][73]  ( .D(block_next[73]), .E(n1199), .CK(clk), .QN(
        n343) );
  EDFFXL \block_reg[6][73]  ( .D(block_next[73]), .E(n1122), .CK(clk), .QN(
        n347) );
  EDFFXL \block_reg[2][72]  ( .D(block_next[72]), .E(n1199), .CK(clk), .Q(
        \block[2][72] ) );
  EDFFXL \block_reg[6][72]  ( .D(block_next[72]), .E(n1122), .CK(clk), .Q(
        \block[6][72] ) );
  EDFFXL \block_reg[2][41]  ( .D(block_next[41]), .E(n1197), .CK(clk), .QN(
        n359) );
  EDFFXL \block_reg[6][41]  ( .D(block_next[41]), .E(n1120), .CK(clk), .QN(
        n363) );
  EDFFXL \block_reg[2][40]  ( .D(block_next[40]), .E(n1197), .CK(clk), .Q(
        \block[2][40] ) );
  EDFFXL \block_reg[6][40]  ( .D(block_next[40]), .E(n1120), .CK(clk), .Q(
        \block[6][40] ) );
  EDFFXL \block_reg[2][6]  ( .D(block_next[6]), .E(n1194), .CK(clk), .Q(
        \block[2][6] ) );
  EDFFXL \block_reg[6][6]  ( .D(block_next[6]), .E(n1117), .CK(clk), .Q(
        \block[6][6] ) );
  EDFFXL \block_reg[2][102]  ( .D(block_next[102]), .E(n1201), .CK(clk), .Q(
        \block[2][102] ) );
  EDFFXL \block_reg[6][102]  ( .D(block_next[102]), .E(n1124), .CK(clk), .Q(
        \block[6][102] ) );
  EDFFXL \block_reg[2][70]  ( .D(block_next[70]), .E(n1199), .CK(clk), .Q(
        \block[2][70] ) );
  EDFFXL \block_reg[6][70]  ( .D(block_next[70]), .E(n1122), .CK(clk), .Q(
        \block[6][70] ) );
  EDFFXL \block_reg[2][38]  ( .D(block_next[38]), .E(n1196), .CK(clk), .Q(
        \block[2][38] ) );
  EDFFXL \block_reg[6][38]  ( .D(block_next[38]), .E(n1119), .CK(clk), .Q(
        \block[6][38] ) );
  EDFFXL \block_reg[2][0]  ( .D(block_next[0]), .E(n1193), .CK(clk), .Q(
        \block[2][0] ) );
  EDFFXL \block_reg[6][0]  ( .D(block_next[0]), .E(n1116), .CK(clk), .Q(
        \block[6][0] ) );
  EDFFXL \block_reg[2][96]  ( .D(block_next[96]), .E(n1201), .CK(clk), .Q(
        \block[2][96] ) );
  EDFFXL \block_reg[6][96]  ( .D(block_next[96]), .E(n1124), .CK(clk), .Q(
        \block[6][96] ) );
  EDFFXL \block_reg[2][64]  ( .D(block_next[64]), .E(n1198), .CK(clk), .Q(
        \block[2][64] ) );
  EDFFXL \block_reg[6][64]  ( .D(block_next[64]), .E(n1121), .CK(clk), .Q(
        \block[6][64] ) );
  EDFFXL \block_reg[2][32]  ( .D(block_next[32]), .E(n1196), .CK(clk), .Q(
        \block[2][32] ) );
  EDFFXL \block_reg[6][32]  ( .D(block_next[32]), .E(n1119), .CK(clk), .Q(
        \block[6][32] ) );
  EDFFXL \block_reg[2][5]  ( .D(block_next[5]), .E(n1194), .CK(clk), .QN(n311)
         );
  EDFFXL \block_reg[6][5]  ( .D(block_next[5]), .E(n1117), .CK(clk), .QN(n315)
         );
  EDFFXL \block_reg[2][7]  ( .D(block_next[7]), .E(n1194), .CK(clk), .Q(
        \block[2][7] ) );
  EDFFXL \block_reg[6][7]  ( .D(block_next[7]), .E(n1117), .CK(clk), .Q(
        \block[6][7] ) );
  EDFFXL \block_reg[2][3]  ( .D(block_next[3]), .E(n1194), .CK(clk), .Q(
        \block[2][3] ) );
  EDFFXL \block_reg[6][3]  ( .D(block_next[3]), .E(n1117), .CK(clk), .Q(
        \block[6][3] ) );
  EDFFXL \block_reg[2][4]  ( .D(block_next[4]), .E(n1194), .CK(clk), .Q(
        \block[2][4] ) );
  EDFFXL \block_reg[2][1]  ( .D(block_next[1]), .E(n1194), .CK(clk), .Q(
        \block[2][1] ) );
  EDFFXL \block_reg[6][4]  ( .D(block_next[4]), .E(n1117), .CK(clk), .Q(
        \block[6][4] ) );
  EDFFXL \block_reg[6][1]  ( .D(block_next[1]), .E(n1117), .CK(clk), .Q(
        \block[6][1] ) );
  EDFFXL \block_reg[2][2]  ( .D(block_next[2]), .E(n1194), .CK(clk), .Q(
        \block[2][2] ) );
  EDFFXL \block_reg[6][2]  ( .D(block_next[2]), .E(n1117), .CK(clk), .Q(
        \block[6][2] ) );
  EDFFXL \block_reg[2][103]  ( .D(block_next[103]), .E(n1201), .CK(clk), .Q(
        \block[2][103] ) );
  EDFFXL \block_reg[6][103]  ( .D(block_next[103]), .E(n1124), .CK(clk), .Q(
        \block[6][103] ) );
  EDFFXL \block_reg[2][101]  ( .D(block_next[101]), .E(n1201), .CK(clk), .Q(
        \block[2][101] ) );
  EDFFXL \block_reg[6][101]  ( .D(block_next[101]), .E(n1124), .CK(clk), .Q(
        \block[6][101] ) );
  EDFFXL \block_reg[2][71]  ( .D(block_next[71]), .E(n1199), .CK(clk), .Q(
        \block[2][71] ) );
  EDFFXL \block_reg[6][71]  ( .D(block_next[71]), .E(n1122), .CK(clk), .Q(
        \block[6][71] ) );
  EDFFXL \block_reg[2][68]  ( .D(block_next[68]), .E(n1199), .CK(clk), .Q(
        \block[2][68] ) );
  EDFFXL \block_reg[6][68]  ( .D(block_next[68]), .E(n1122), .CK(clk), .Q(
        \block[6][68] ) );
  EDFFXL \block_reg[2][67]  ( .D(block_next[67]), .E(n1199), .CK(clk), .Q(
        \block[2][67] ) );
  EDFFXL \block_reg[2][37]  ( .D(block_next[37]), .E(n1196), .CK(clk), .Q(
        \block[2][37] ) );
  EDFFXL \block_reg[6][67]  ( .D(block_next[67]), .E(n1122), .CK(clk), .Q(
        \block[6][67] ) );
  EDFFXL \block_reg[2][39]  ( .D(block_next[39]), .E(n1196), .CK(clk), .Q(
        \block[2][39] ) );
  EDFFXL \block_reg[6][37]  ( .D(block_next[37]), .E(n1119), .CK(clk), .Q(
        \block[6][37] ) );
  EDFFXL \block_reg[6][39]  ( .D(block_next[39]), .E(n1119), .CK(clk), .Q(
        \block[6][39] ) );
  EDFFXL \block_reg[2][69]  ( .D(block_next[69]), .E(n1199), .CK(clk), .Q(
        \block[2][69] ) );
  EDFFXL \block_reg[2][100]  ( .D(block_next[100]), .E(n1201), .CK(clk), .Q(
        \block[2][100] ) );
  EDFFXL \block_reg[6][69]  ( .D(block_next[69]), .E(n1122), .CK(clk), .Q(
        \block[6][69] ) );
  EDFFXL \block_reg[6][100]  ( .D(block_next[100]), .E(n1124), .CK(clk), .Q(
        \block[6][100] ) );
  EDFFXL \block_reg[2][99]  ( .D(block_next[99]), .E(n1201), .CK(clk), .Q(
        \block[2][99] ) );
  EDFFXL \block_reg[6][99]  ( .D(block_next[99]), .E(n1124), .CK(clk), .Q(
        \block[6][99] ) );
  EDFFXL \block_reg[2][97]  ( .D(block_next[97]), .E(n1201), .CK(clk), .Q(
        \block[2][97] ) );
  EDFFXL \block_reg[6][97]  ( .D(block_next[97]), .E(n1124), .CK(clk), .Q(
        \block[6][97] ) );
  EDFFXL \block_reg[2][65]  ( .D(block_next[65]), .E(n1198), .CK(clk), .Q(
        \block[2][65] ) );
  EDFFXL \block_reg[6][65]  ( .D(block_next[65]), .E(n1121), .CK(clk), .Q(
        \block[6][65] ) );
  EDFFXL \block_reg[2][36]  ( .D(block_next[36]), .E(n1196), .CK(clk), .QN(
        n319) );
  EDFFXL \block_reg[2][98]  ( .D(block_next[98]), .E(n1201), .CK(clk), .Q(
        \block[2][98] ) );
  EDFFXL \block_reg[6][36]  ( .D(block_next[36]), .E(n1119), .CK(clk), .QN(
        n323) );
  EDFFXL \block_reg[6][98]  ( .D(block_next[98]), .E(n1124), .CK(clk), .Q(
        \block[6][98] ) );
  EDFFXL \block_reg[2][66]  ( .D(block_next[66]), .E(n1199), .CK(clk), .Q(
        \block[2][66] ) );
  EDFFXL \block_reg[6][66]  ( .D(block_next[66]), .E(n1122), .CK(clk), .Q(
        \block[6][66] ) );
  EDFFXL \block_reg[2][35]  ( .D(block_next[35]), .E(n1196), .CK(clk), .Q(
        \block[2][35] ) );
  EDFFXL \block_reg[6][35]  ( .D(block_next[35]), .E(n1119), .CK(clk), .Q(
        \block[6][35] ) );
  EDFFXL \block_reg[2][33]  ( .D(block_next[33]), .E(n1196), .CK(clk), .Q(
        \block[2][33] ) );
  EDFFXL \block_reg[6][33]  ( .D(block_next[33]), .E(n1119), .CK(clk), .Q(
        \block[6][33] ) );
  EDFFXL \block_reg[2][34]  ( .D(block_next[34]), .E(n1196), .CK(clk), .Q(
        \block[2][34] ) );
  EDFFXL \block_reg[6][34]  ( .D(block_next[34]), .E(n1119), .CK(clk), .Q(
        \block[6][34] ) );
  EDFFXL \block_reg[2][122]  ( .D(block_next[122]), .E(n1203), .CK(clk), .Q(
        \block[2][122] ) );
  EDFFXL \block_reg[6][122]  ( .D(block_next[122]), .E(n1126), .CK(clk), .Q(
        \block[6][122] ) );
  EDFFXL \block_reg[2][26]  ( .D(block_next[26]), .E(n1195), .CK(clk), .QN(
        n293) );
  EDFFXL \block_reg[6][26]  ( .D(block_next[26]), .E(n1118), .CK(clk), .QN(
        n297) );
  DFFRX1 \blockdirty_reg[7]  ( .D(n1724), .CK(clk), .RN(n1259), .Q(
        blockdirty[7]), .QN(n1740) );
  DFFRX1 \blockdirty_reg[6]  ( .D(n1725), .CK(clk), .RN(n1259), .Q(
        blockdirty[6]), .QN(n1741) );
  EDFFXL \block_reg[3][30]  ( .D(block_next[30]), .E(n1177), .CK(clk), .Q(
        \block[3][30] ) );
  EDFFXL \block_reg[7][30]  ( .D(block_next[30]), .E(n1104), .CK(clk), .Q(
        \block[7][30] ) );
  EDFFXL \block_reg[3][29]  ( .D(block_next[29]), .E(n1177), .CK(clk), .Q(
        \block[3][29] ) );
  EDFFXL \block_reg[7][29]  ( .D(block_next[29]), .E(n1104), .CK(clk), .Q(
        \block[7][29] ) );
  EDFFXL \block_reg[3][126]  ( .D(block_next[126]), .E(n1184), .CK(clk), .QN(
        n274) );
  EDFFXL \block_reg[7][126]  ( .D(block_next[126]), .E(n1111), .CK(clk), .QN(
        n278) );
  EDFFXL \block_reg[3][125]  ( .D(block_next[125]), .E(n1184), .CK(clk), .Q(
        \block[3][125] ) );
  EDFFXL \block_reg[7][125]  ( .D(block_next[125]), .E(n1111), .CK(clk), .Q(
        \block[7][125] ) );
  EDFFXL \block_reg[3][94]  ( .D(block_next[94]), .E(n1182), .CK(clk), .QN(
        n282) );
  EDFFXL \block_reg[7][94]  ( .D(block_next[94]), .E(n1109), .CK(clk), .Q(
        \block[7][94] ) );
  EDFFXL \block_reg[3][93]  ( .D(block_next[93]), .E(n1182), .CK(clk), .Q(
        \block[3][93] ) );
  EDFFXL \block_reg[7][93]  ( .D(block_next[93]), .E(n1109), .CK(clk), .Q(
        \block[7][93] ) );
  EDFFXL \block_reg[3][62]  ( .D(block_next[62]), .E(n1179), .CK(clk), .QN(
        n270) );
  EDFFXL \block_reg[7][62]  ( .D(block_next[62]), .E(n1106), .CK(clk), .Q(
        \block[7][62] ) );
  EDFFXL \block_reg[3][61]  ( .D(block_next[61]), .E(n1179), .CK(clk), .Q(
        \block[3][61] ) );
  EDFFXL \block_reg[7][61]  ( .D(block_next[61]), .E(n1106), .CK(clk), .Q(
        \block[7][61] ) );
  EDFFXL \block_reg[3][90]  ( .D(block_next[90]), .E(n1181), .CK(clk), .QN(
        n304) );
  EDFFXL \block_reg[7][90]  ( .D(block_next[90]), .E(n1108), .CK(clk), .QN(
        n308) );
  EDFFXL \block_reg[3][58]  ( .D(block_next[58]), .E(n1179), .CK(clk), .QN(
        n286) );
  EDFFXL \block_reg[7][58]  ( .D(block_next[58]), .E(n1106), .CK(clk), .QN(
        n290) );
  EDFFXL \block_reg[3][27]  ( .D(block_next[27]), .E(n1177), .CK(clk), .Q(
        \block[3][27] ) );
  EDFFXL \block_reg[7][27]  ( .D(block_next[27]), .E(n1104), .CK(clk), .Q(
        \block[7][27] ) );
  EDFFXL \block_reg[3][123]  ( .D(block_next[123]), .E(n1184), .CK(clk), .Q(
        \block[3][123] ) );
  EDFFXL \block_reg[7][123]  ( .D(block_next[123]), .E(n1111), .CK(clk), .Q(
        \block[7][123] ) );
  EDFFXL \block_reg[3][91]  ( .D(block_next[91]), .E(n1181), .CK(clk), .Q(
        \block[3][91] ) );
  EDFFXL \block_reg[7][91]  ( .D(block_next[91]), .E(n1108), .CK(clk), .Q(
        \block[7][91] ) );
  EDFFXL \block_reg[3][59]  ( .D(block_next[59]), .E(n1179), .CK(clk), .Q(
        \block[3][59] ) );
  EDFFXL \block_reg[7][59]  ( .D(block_next[59]), .E(n1106), .CK(clk), .Q(
        \block[7][59] ) );
  EDFFXL \block_reg[3][28]  ( .D(block_next[28]), .E(n1177), .CK(clk), .QN(
        n663) );
  EDFFXL \block_reg[7][28]  ( .D(block_next[28]), .E(n1104), .CK(clk), .QN(
        n667) );
  EDFFXL \block_reg[3][124]  ( .D(block_next[124]), .E(n1184), .CK(clk), .QN(
        n655) );
  EDFFXL \block_reg[7][124]  ( .D(block_next[124]), .E(n1111), .CK(clk), .QN(
        n659) );
  EDFFXL \block_reg[3][92]  ( .D(block_next[92]), .E(n1182), .CK(clk), .QN(
        n647) );
  EDFFXL \block_reg[7][92]  ( .D(block_next[92]), .E(n1109), .CK(clk), .QN(
        n651) );
  EDFFXL \block_reg[3][60]  ( .D(block_next[60]), .E(n1179), .CK(clk), .QN(
        n639) );
  EDFFXL \block_reg[7][60]  ( .D(block_next[60]), .E(n1106), .CK(clk), .QN(
        n643) );
  EDFFXL \block_reg[3][31]  ( .D(block_next[31]), .E(n1177), .CK(clk), .QN(
        n635) );
  EDFFXL \block_reg[7][31]  ( .D(block_next[31]), .E(n1104), .CK(clk), .Q(
        \block[7][31] ) );
  EDFFXL \block_reg[3][127]  ( .D(block_next[127]), .E(n1184), .CK(clk), .Q(
        \block[3][127] ) );
  EDFFXL \block_reg[7][127]  ( .D(block_next[127]), .E(n1111), .CK(clk), .QN(
        n631) );
  EDFFXL \block_reg[3][95]  ( .D(block_next[95]), .E(n1182), .CK(clk), .Q(
        \block[3][95] ) );
  EDFFXL \block_reg[7][95]  ( .D(block_next[95]), .E(n1109), .CK(clk), .QN(
        n627) );
  EDFFXL \block_reg[3][63]  ( .D(block_next[63]), .E(n1179), .CK(clk), .Q(
        \block[3][63] ) );
  EDFFXL \block_reg[7][63]  ( .D(block_next[63]), .E(n1106), .CK(clk), .QN(
        n623) );
  EDFFXL \block_reg[1][30]  ( .D(block_next[30]), .E(n1215), .CK(clk), .Q(
        \block[1][30] ) );
  EDFFXL \block_reg[5][30]  ( .D(block_next[30]), .E(n1139), .CK(clk), .Q(
        \block[5][30] ) );
  EDFFXL \block_reg[1][29]  ( .D(block_next[29]), .E(n1215), .CK(clk), .Q(
        \block[1][29] ) );
  EDFFXL \block_reg[5][29]  ( .D(block_next[29]), .E(n1139), .CK(clk), .Q(
        \block[5][29] ) );
  EDFFXL \block_reg[1][126]  ( .D(block_next[126]), .E(n1222), .CK(clk), .QN(
        n272) );
  EDFFXL \block_reg[5][126]  ( .D(block_next[126]), .E(n1146), .CK(clk), .QN(
        n276) );
  EDFFXL \block_reg[1][125]  ( .D(block_next[125]), .E(n1222), .CK(clk), .Q(
        \block[1][125] ) );
  EDFFXL \block_reg[5][125]  ( .D(block_next[125]), .E(n1146), .CK(clk), .Q(
        \block[5][125] ) );
  EDFFXL \block_reg[1][94]  ( .D(block_next[94]), .E(n1220), .CK(clk), .QN(
        n280) );
  EDFFXL \block_reg[5][94]  ( .D(block_next[94]), .E(n1144), .CK(clk), .Q(
        \block[5][94] ) );
  EDFFXL \block_reg[1][93]  ( .D(block_next[93]), .E(n1220), .CK(clk), .Q(
        \block[1][93] ) );
  EDFFXL \block_reg[5][93]  ( .D(block_next[93]), .E(n1144), .CK(clk), .Q(
        \block[5][93] ) );
  EDFFXL \block_reg[1][62]  ( .D(block_next[62]), .E(n1217), .CK(clk), .QN(
        n268) );
  EDFFXL \block_reg[5][62]  ( .D(block_next[62]), .E(n1141), .CK(clk), .Q(
        \block[5][62] ) );
  EDFFXL \block_reg[1][61]  ( .D(block_next[61]), .E(n1217), .CK(clk), .Q(
        \block[1][61] ) );
  EDFFXL \block_reg[5][61]  ( .D(block_next[61]), .E(n1141), .CK(clk), .Q(
        \block[5][61] ) );
  EDFFXL \block_reg[1][90]  ( .D(block_next[90]), .E(n1219), .CK(clk), .QN(
        n302) );
  EDFFXL \block_reg[5][90]  ( .D(block_next[90]), .E(n1143), .CK(clk), .QN(
        n306) );
  EDFFXL \block_reg[1][58]  ( .D(block_next[58]), .E(n1217), .CK(clk), .QN(
        n284) );
  EDFFXL \block_reg[5][58]  ( .D(block_next[58]), .E(n1141), .CK(clk), .QN(
        n288) );
  EDFFXL \block_reg[1][27]  ( .D(block_next[27]), .E(n1215), .CK(clk), .Q(
        \block[1][27] ) );
  EDFFXL \block_reg[5][27]  ( .D(block_next[27]), .E(n1139), .CK(clk), .Q(
        \block[5][27] ) );
  EDFFXL \block_reg[1][123]  ( .D(block_next[123]), .E(n1222), .CK(clk), .Q(
        \block[1][123] ) );
  EDFFXL \block_reg[5][123]  ( .D(block_next[123]), .E(n1146), .CK(clk), .Q(
        \block[5][123] ) );
  EDFFXL \block_reg[1][91]  ( .D(block_next[91]), .E(n1219), .CK(clk), .Q(
        \block[1][91] ) );
  EDFFXL \block_reg[5][91]  ( .D(block_next[91]), .E(n1143), .CK(clk), .Q(
        \block[5][91] ) );
  EDFFXL \block_reg[1][59]  ( .D(block_next[59]), .E(n1217), .CK(clk), .Q(
        \block[1][59] ) );
  EDFFXL \block_reg[5][59]  ( .D(block_next[59]), .E(n1141), .CK(clk), .Q(
        \block[5][59] ) );
  EDFFXL \block_reg[1][28]  ( .D(block_next[28]), .E(n1215), .CK(clk), .QN(
        n661) );
  EDFFXL \block_reg[5][28]  ( .D(block_next[28]), .E(n1139), .CK(clk), .QN(
        n665) );
  EDFFXL \block_reg[1][124]  ( .D(block_next[124]), .E(n1222), .CK(clk), .QN(
        n653) );
  EDFFXL \block_reg[5][124]  ( .D(block_next[124]), .E(n1146), .CK(clk), .QN(
        n657) );
  EDFFXL \block_reg[1][92]  ( .D(block_next[92]), .E(n1220), .CK(clk), .QN(
        n645) );
  EDFFXL \block_reg[5][92]  ( .D(block_next[92]), .E(n1144), .CK(clk), .QN(
        n649) );
  EDFFXL \block_reg[1][60]  ( .D(block_next[60]), .E(n1217), .CK(clk), .QN(
        n637) );
  EDFFXL \block_reg[5][60]  ( .D(block_next[60]), .E(n1141), .CK(clk), .QN(
        n641) );
  EDFFXL \block_reg[1][31]  ( .D(block_next[31]), .E(n1215), .CK(clk), .QN(
        n633) );
  EDFFXL \block_reg[5][31]  ( .D(block_next[31]), .E(n1139), .CK(clk), .Q(
        \block[5][31] ) );
  EDFFXL \block_reg[1][127]  ( .D(block_next[127]), .E(n1222), .CK(clk), .Q(
        \block[1][127] ) );
  EDFFXL \block_reg[5][127]  ( .D(block_next[127]), .E(n1146), .CK(clk), .QN(
        n629) );
  EDFFXL \block_reg[1][95]  ( .D(block_next[95]), .E(n1220), .CK(clk), .Q(
        \block[1][95] ) );
  EDFFXL \block_reg[5][95]  ( .D(block_next[95]), .E(n1144), .CK(clk), .QN(
        n625) );
  EDFFXL \block_reg[1][63]  ( .D(block_next[63]), .E(n1217), .CK(clk), .Q(
        \block[1][63] ) );
  EDFFXL \block_reg[5][63]  ( .D(block_next[63]), .E(n1141), .CK(clk), .QN(
        n621) );
  EDFFXL \block_reg[0][30]  ( .D(block_next[30]), .E(n1234), .CK(clk), .Q(
        \block[0][30] ) );
  EDFFXL \block_reg[4][30]  ( .D(block_next[30]), .E(n1158), .CK(clk), .Q(
        \block[4][30] ) );
  EDFFXL \block_reg[0][29]  ( .D(block_next[29]), .E(n1234), .CK(clk), .Q(
        \block[0][29] ) );
  EDFFXL \block_reg[4][29]  ( .D(block_next[29]), .E(n1158), .CK(clk), .Q(
        \block[4][29] ) );
  EDFFXL \block_reg[0][126]  ( .D(block_next[126]), .E(n1241), .CK(clk), .QN(
        n271) );
  EDFFXL \block_reg[4][126]  ( .D(block_next[126]), .E(n1165), .CK(clk), .QN(
        n275) );
  EDFFXL \block_reg[0][125]  ( .D(block_next[125]), .E(n1241), .CK(clk), .Q(
        \block[0][125] ) );
  EDFFXL \block_reg[4][125]  ( .D(block_next[125]), .E(n1165), .CK(clk), .Q(
        \block[4][125] ) );
  EDFFXL \block_reg[0][94]  ( .D(block_next[94]), .E(n1239), .CK(clk), .QN(
        n279) );
  EDFFXL \block_reg[4][94]  ( .D(block_next[94]), .E(n1163), .CK(clk), .Q(
        \block[4][94] ) );
  EDFFXL \block_reg[0][93]  ( .D(block_next[93]), .E(n1239), .CK(clk), .Q(
        \block[0][93] ) );
  EDFFXL \block_reg[4][93]  ( .D(block_next[93]), .E(n1163), .CK(clk), .Q(
        \block[4][93] ) );
  EDFFXL \block_reg[0][62]  ( .D(block_next[62]), .E(n1236), .CK(clk), .QN(
        n267) );
  EDFFXL \block_reg[4][62]  ( .D(block_next[62]), .E(n1160), .CK(clk), .Q(
        \block[4][62] ) );
  EDFFXL \block_reg[0][61]  ( .D(block_next[61]), .E(n1236), .CK(clk), .Q(
        \block[0][61] ) );
  EDFFXL \block_reg[4][61]  ( .D(block_next[61]), .E(n1160), .CK(clk), .Q(
        \block[4][61] ) );
  EDFFXL \block_reg[0][90]  ( .D(block_next[90]), .E(n1238), .CK(clk), .QN(
        n301) );
  EDFFXL \block_reg[4][90]  ( .D(block_next[90]), .E(n1162), .CK(clk), .QN(
        n305) );
  EDFFXL \block_reg[0][58]  ( .D(block_next[58]), .E(n1236), .CK(clk), .QN(
        n283) );
  EDFFXL \block_reg[4][58]  ( .D(block_next[58]), .E(n1160), .CK(clk), .QN(
        n287) );
  EDFFXL \block_reg[0][27]  ( .D(block_next[27]), .E(n1234), .CK(clk), .Q(
        \block[0][27] ) );
  EDFFXL \block_reg[4][27]  ( .D(block_next[27]), .E(n1158), .CK(clk), .Q(
        \block[4][27] ) );
  EDFFXL \block_reg[0][123]  ( .D(block_next[123]), .E(n1241), .CK(clk), .Q(
        \block[0][123] ) );
  EDFFXL \block_reg[4][123]  ( .D(block_next[123]), .E(n1165), .CK(clk), .Q(
        \block[4][123] ) );
  EDFFXL \block_reg[0][91]  ( .D(block_next[91]), .E(n1238), .CK(clk), .Q(
        \block[0][91] ) );
  EDFFXL \block_reg[4][91]  ( .D(block_next[91]), .E(n1162), .CK(clk), .Q(
        \block[4][91] ) );
  EDFFXL \block_reg[0][59]  ( .D(block_next[59]), .E(n1236), .CK(clk), .Q(
        \block[0][59] ) );
  EDFFXL \block_reg[4][59]  ( .D(block_next[59]), .E(n1160), .CK(clk), .Q(
        \block[4][59] ) );
  EDFFXL \block_reg[0][28]  ( .D(block_next[28]), .E(n1234), .CK(clk), .QN(
        n660) );
  EDFFXL \block_reg[4][28]  ( .D(block_next[28]), .E(n1158), .CK(clk), .QN(
        n664) );
  EDFFXL \block_reg[0][124]  ( .D(block_next[124]), .E(n1241), .CK(clk), .QN(
        n652) );
  EDFFXL \block_reg[4][124]  ( .D(block_next[124]), .E(n1165), .CK(clk), .QN(
        n656) );
  EDFFXL \block_reg[0][92]  ( .D(block_next[92]), .E(n1239), .CK(clk), .QN(
        n644) );
  EDFFXL \block_reg[4][92]  ( .D(block_next[92]), .E(n1163), .CK(clk), .QN(
        n648) );
  EDFFXL \block_reg[0][60]  ( .D(block_next[60]), .E(n1236), .CK(clk), .QN(
        n636) );
  EDFFXL \block_reg[4][60]  ( .D(block_next[60]), .E(n1160), .CK(clk), .QN(
        n640) );
  EDFFXL \block_reg[0][31]  ( .D(block_next[31]), .E(n1234), .CK(clk), .QN(
        n632) );
  EDFFXL \block_reg[4][31]  ( .D(block_next[31]), .E(n1158), .CK(clk), .Q(
        \block[4][31] ) );
  EDFFXL \block_reg[0][127]  ( .D(block_next[127]), .E(n1241), .CK(clk), .Q(
        \block[0][127] ) );
  EDFFXL \block_reg[4][127]  ( .D(block_next[127]), .E(n1165), .CK(clk), .QN(
        n628) );
  EDFFXL \block_reg[0][95]  ( .D(block_next[95]), .E(n1239), .CK(clk), .Q(
        \block[0][95] ) );
  EDFFXL \block_reg[4][95]  ( .D(block_next[95]), .E(n1163), .CK(clk), .QN(
        n624) );
  EDFFXL \block_reg[0][63]  ( .D(block_next[63]), .E(n1236), .CK(clk), .Q(
        \block[0][63] ) );
  EDFFXL \block_reg[4][63]  ( .D(block_next[63]), .E(n1160), .CK(clk), .QN(
        n620) );
  EDFFXL \block_reg[2][30]  ( .D(block_next[30]), .E(n1196), .CK(clk), .Q(
        \block[2][30] ) );
  EDFFXL \block_reg[6][30]  ( .D(block_next[30]), .E(n1119), .CK(clk), .Q(
        \block[6][30] ) );
  EDFFXL \block_reg[2][29]  ( .D(block_next[29]), .E(n1196), .CK(clk), .Q(
        \block[2][29] ) );
  EDFFXL \block_reg[6][29]  ( .D(block_next[29]), .E(n1119), .CK(clk), .Q(
        \block[6][29] ) );
  EDFFXL \block_reg[2][126]  ( .D(block_next[126]), .E(n1203), .CK(clk), .QN(
        n273) );
  EDFFXL \block_reg[6][126]  ( .D(block_next[126]), .E(n1126), .CK(clk), .QN(
        n277) );
  EDFFXL \block_reg[2][125]  ( .D(block_next[125]), .E(n1203), .CK(clk), .Q(
        \block[2][125] ) );
  EDFFXL \block_reg[6][125]  ( .D(block_next[125]), .E(n1126), .CK(clk), .Q(
        \block[6][125] ) );
  EDFFXL \block_reg[2][94]  ( .D(block_next[94]), .E(n1201), .CK(clk), .QN(
        n281) );
  EDFFXL \block_reg[6][94]  ( .D(block_next[94]), .E(n1124), .CK(clk), .Q(
        \block[6][94] ) );
  EDFFXL \block_reg[2][93]  ( .D(block_next[93]), .E(n1201), .CK(clk), .Q(
        \block[2][93] ) );
  EDFFXL \block_reg[6][93]  ( .D(block_next[93]), .E(n1124), .CK(clk), .Q(
        \block[6][93] ) );
  EDFFXL \block_reg[2][62]  ( .D(block_next[62]), .E(n1198), .CK(clk), .QN(
        n269) );
  EDFFXL \block_reg[6][62]  ( .D(block_next[62]), .E(n1121), .CK(clk), .Q(
        \block[6][62] ) );
  EDFFXL \block_reg[2][61]  ( .D(block_next[61]), .E(n1198), .CK(clk), .Q(
        \block[2][61] ) );
  EDFFXL \block_reg[6][61]  ( .D(block_next[61]), .E(n1121), .CK(clk), .Q(
        \block[6][61] ) );
  EDFFXL \block_reg[2][90]  ( .D(block_next[90]), .E(n1200), .CK(clk), .QN(
        n303) );
  EDFFXL \block_reg[6][90]  ( .D(block_next[90]), .E(n1123), .CK(clk), .QN(
        n307) );
  EDFFXL \block_reg[2][58]  ( .D(block_next[58]), .E(n1198), .CK(clk), .QN(
        n285) );
  EDFFXL \block_reg[6][58]  ( .D(block_next[58]), .E(n1121), .CK(clk), .QN(
        n289) );
  EDFFXL \block_reg[2][27]  ( .D(block_next[27]), .E(n1196), .CK(clk), .Q(
        \block[2][27] ) );
  EDFFXL \block_reg[6][27]  ( .D(block_next[27]), .E(n1119), .CK(clk), .Q(
        \block[6][27] ) );
  EDFFXL \block_reg[2][123]  ( .D(block_next[123]), .E(n1203), .CK(clk), .Q(
        \block[2][123] ) );
  EDFFXL \block_reg[6][123]  ( .D(block_next[123]), .E(n1126), .CK(clk), .Q(
        \block[6][123] ) );
  EDFFXL \block_reg[2][91]  ( .D(block_next[91]), .E(n1200), .CK(clk), .Q(
        \block[2][91] ) );
  EDFFXL \block_reg[6][91]  ( .D(block_next[91]), .E(n1123), .CK(clk), .Q(
        \block[6][91] ) );
  EDFFXL \block_reg[2][59]  ( .D(block_next[59]), .E(n1198), .CK(clk), .Q(
        \block[2][59] ) );
  EDFFXL \block_reg[6][59]  ( .D(block_next[59]), .E(n1121), .CK(clk), .Q(
        \block[6][59] ) );
  EDFFXL \block_reg[2][28]  ( .D(block_next[28]), .E(n1196), .CK(clk), .QN(
        n662) );
  EDFFXL \block_reg[6][28]  ( .D(block_next[28]), .E(n1119), .CK(clk), .QN(
        n666) );
  EDFFXL \block_reg[2][124]  ( .D(block_next[124]), .E(n1203), .CK(clk), .QN(
        n654) );
  EDFFXL \block_reg[6][124]  ( .D(block_next[124]), .E(n1126), .CK(clk), .QN(
        n658) );
  EDFFXL \block_reg[2][92]  ( .D(block_next[92]), .E(n1201), .CK(clk), .QN(
        n646) );
  EDFFXL \block_reg[6][92]  ( .D(block_next[92]), .E(n1124), .CK(clk), .QN(
        n650) );
  EDFFXL \block_reg[2][60]  ( .D(block_next[60]), .E(n1198), .CK(clk), .QN(
        n638) );
  EDFFXL \block_reg[6][60]  ( .D(block_next[60]), .E(n1121), .CK(clk), .QN(
        n642) );
  EDFFXL \block_reg[2][31]  ( .D(block_next[31]), .E(n1196), .CK(clk), .QN(
        n634) );
  EDFFXL \block_reg[6][31]  ( .D(block_next[31]), .E(n1119), .CK(clk), .Q(
        \block[6][31] ) );
  EDFFXL \block_reg[2][127]  ( .D(block_next[127]), .E(n1203), .CK(clk), .Q(
        \block[2][127] ) );
  EDFFXL \block_reg[6][127]  ( .D(block_next[127]), .E(n1126), .CK(clk), .QN(
        n630) );
  EDFFXL \block_reg[2][95]  ( .D(block_next[95]), .E(n1201), .CK(clk), .Q(
        \block[2][95] ) );
  EDFFXL \block_reg[6][95]  ( .D(block_next[95]), .E(n1124), .CK(clk), .QN(
        n626) );
  EDFFXL \block_reg[2][63]  ( .D(block_next[63]), .E(n1198), .CK(clk), .Q(
        \block[2][63] ) );
  EDFFXL \block_reg[6][63]  ( .D(block_next[63]), .E(n1121), .CK(clk), .QN(
        n622) );
  DFFRX1 \blockdirty_reg[3]  ( .D(n1728), .CK(clk), .RN(n1258), .Q(
        blockdirty[3]), .QN(n1744) );
  DFFRX1 \blockdirty_reg[5]  ( .D(n1726), .CK(clk), .RN(n1258), .Q(
        blockdirty[5]), .QN(n1742) );
  DFFRX1 \blockdirty_reg[1]  ( .D(n1730), .CK(clk), .RN(n1258), .Q(
        blockdirty[1]), .QN(n1746) );
  DFFRX1 \blockdirty_reg[4]  ( .D(n1727), .CK(clk), .RN(n1258), .Q(
        blockdirty[4]), .QN(n1743) );
  DFFRX1 \blockdirty_reg[0]  ( .D(n1731), .CK(clk), .RN(n1258), .Q(
        blockdirty[0]), .QN(n1747) );
  DFFRX1 \blockdirty_reg[2]  ( .D(n1729), .CK(clk), .RN(n1258), .Q(
        blockdirty[2]), .QN(n1745) );
  EDFFX1 \blocktag_reg[3][20]  ( .D(blocktag_next[20]), .E(n1174), .CK(clk), 
        .QN(n205) );
  EDFFX1 \blocktag_reg[7][20]  ( .D(blocktag_next[20]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][20] ) );
  EDFFX1 \blocktag_reg[3][19]  ( .D(blocktag_next[19]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][19] ) );
  EDFFX1 \blocktag_reg[3][0]  ( .D(n4), .E(n1173), .CK(clk), .Q(
        \blocktag[3][0] ) );
  EDFFX1 \blocktag_reg[7][19]  ( .D(blocktag_next[19]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][19] ) );
  EDFFX1 \blocktag_reg[7][0]  ( .D(n4), .E(n1100), .CK(clk), .Q(
        \blocktag[7][0] ) );
  EDFFX1 \blocktag_reg[3][23]  ( .D(blocktag_next[23]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][23] ) );
  EDFFX1 \blocktag_reg[3][24]  ( .D(blocktag_next[24]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][24] ) );
  EDFFX1 \blocktag_reg[7][23]  ( .D(blocktag_next[23]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][23] ) );
  EDFFX1 \blocktag_reg[7][24]  ( .D(blocktag_next[24]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][24] ) );
  EDFFX1 \blocktag_reg[3][2]  ( .D(blocktag_next[2]), .E(n1173), .CK(clk), .Q(
        \blocktag[3][2] ) );
  EDFFX1 \blocktag_reg[7][2]  ( .D(blocktag_next[2]), .E(n1100), .CK(clk), .Q(
        \blocktag[7][2] ) );
  EDFFX1 \blocktag_reg[3][11]  ( .D(blocktag_next[11]), .E(n1173), .CK(clk), 
        .Q(\blocktag[3][11] ) );
  EDFFX1 \blocktag_reg[7][11]  ( .D(blocktag_next[11]), .E(n1100), .CK(clk), 
        .Q(\blocktag[7][11] ) );
  EDFFX1 \blocktag_reg[3][1]  ( .D(blocktag_next[1]), .E(n1173), .CK(clk), .Q(
        \blocktag[3][1] ) );
  EDFFX1 \blocktag_reg[7][1]  ( .D(blocktag_next[1]), .E(n1100), .CK(clk), 
        .QN(n609) );
  EDFFX1 \blocktag_reg[3][18]  ( .D(blocktag_next[18]), .E(n1174), .CK(clk), 
        .QN(n593) );
  EDFFX1 \blocktag_reg[7][18]  ( .D(blocktag_next[18]), .E(n1101), .CK(clk), 
        .QN(n597) );
  EDFFX1 \blocktag_reg[3][12]  ( .D(blocktag_next[12]), .E(n1173), .CK(clk), 
        .Q(n256) );
  EDFFX1 \blocktag_reg[3][3]  ( .D(blocktag_next[3]), .E(n1173), .CK(clk), 
        .QN(n585) );
  EDFFX1 \blocktag_reg[7][12]  ( .D(blocktag_next[12]), .E(n1100), .CK(clk), 
        .Q(n252) );
  EDFFX1 \blocktag_reg[7][3]  ( .D(blocktag_next[3]), .E(n1100), .CK(clk), 
        .QN(n589) );
  EDFFX1 \blocktag_reg[3][17]  ( .D(blocktag_next[17]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][17] ) );
  EDFFX1 \blocktag_reg[7][17]  ( .D(blocktag_next[17]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][17] ) );
  EDFFX1 \blocktag_reg[3][5]  ( .D(blocktag_next[5]), .E(n1173), .CK(clk), 
        .QN(n577) );
  EDFFX1 \blocktag_reg[3][14]  ( .D(blocktag_next[14]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][14] ) );
  EDFFX1 \blocktag_reg[7][5]  ( .D(blocktag_next[5]), .E(n1100), .CK(clk), 
        .QN(n581) );
  EDFFX1 \blocktag_reg[3][22]  ( .D(blocktag_next[22]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][22] ) );
  EDFFX1 \blocktag_reg[7][14]  ( .D(blocktag_next[14]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][14] ) );
  EDFFX1 \blocktag_reg[7][22]  ( .D(blocktag_next[22]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][22] ) );
  EDFFX1 \blocktag_reg[3][16]  ( .D(blocktag_next[16]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][16] ) );
  EDFFX1 \blocktag_reg[7][16]  ( .D(blocktag_next[16]), .E(n1101), .CK(clk), 
        .Q(n248) );
  EDFFX1 \blocktag_reg[3][10]  ( .D(blocktag_next[10]), .E(n1173), .CK(clk), 
        .Q(\blocktag[3][10] ) );
  EDFFX1 \blocktag_reg[7][10]  ( .D(blocktag_next[10]), .E(n1100), .CK(clk), 
        .Q(\blocktag[7][10] ) );
  EDFFX1 \blocktag_reg[3][7]  ( .D(n3), .E(n1173), .CK(clk), .Q(n244) );
  EDFFX1 \blocktag_reg[7][7]  ( .D(n3), .E(n1100), .CK(clk), .Q(n240) );
  EDFFX1 \blocktag_reg[3][15]  ( .D(blocktag_next[15]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][15] ) );
  EDFFX1 \blocktag_reg[3][8]  ( .D(blocktag_next[8]), .E(n1173), .CK(clk), .Q(
        n236) );
  EDFFX1 \blocktag_reg[7][15]  ( .D(blocktag_next[15]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][15] ) );
  EDFFX1 \blocktag_reg[7][8]  ( .D(blocktag_next[8]), .E(n1100), .CK(clk), .Q(
        n232) );
  EDFFX1 \blocktag_reg[3][13]  ( .D(blocktag_next[13]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][13] ) );
  EDFFX1 \blocktag_reg[7][13]  ( .D(blocktag_next[13]), .E(n1101), .CK(clk), 
        .Q(\blocktag[7][13] ) );
  EDFFX1 \blocktag_reg[1][20]  ( .D(blocktag_next[20]), .E(n1212), .CK(clk), 
        .QN(n203) );
  EDFFX1 \blocktag_reg[5][20]  ( .D(blocktag_next[20]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][20] ) );
  EDFFX1 \blocktag_reg[1][19]  ( .D(blocktag_next[19]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][19] ) );
  EDFFX1 \blocktag_reg[1][0]  ( .D(n4), .E(n1211), .CK(clk), .Q(
        \blocktag[1][0] ) );
  EDFFX1 \blocktag_reg[5][19]  ( .D(blocktag_next[19]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][19] ) );
  EDFFX1 \blocktag_reg[5][0]  ( .D(n4), .E(n1135), .CK(clk), .Q(
        \blocktag[5][0] ) );
  EDFFX1 \blocktag_reg[1][23]  ( .D(blocktag_next[23]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][23] ) );
  EDFFX1 \blocktag_reg[1][24]  ( .D(blocktag_next[24]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][24] ) );
  EDFFX1 \blocktag_reg[5][23]  ( .D(blocktag_next[23]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][23] ) );
  EDFFX1 \blocktag_reg[5][24]  ( .D(blocktag_next[24]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][24] ) );
  EDFFX1 \blocktag_reg[1][2]  ( .D(blocktag_next[2]), .E(n1211), .CK(clk), .Q(
        \blocktag[1][2] ) );
  EDFFX1 \blocktag_reg[5][2]  ( .D(blocktag_next[2]), .E(n1135), .CK(clk), .Q(
        \blocktag[5][2] ) );
  EDFFX1 \blocktag_reg[1][11]  ( .D(blocktag_next[11]), .E(n1211), .CK(clk), 
        .Q(\blocktag[1][11] ) );
  EDFFX1 \blocktag_reg[5][11]  ( .D(blocktag_next[11]), .E(n1135), .CK(clk), 
        .Q(\blocktag[5][11] ) );
  EDFFX1 \blocktag_reg[1][1]  ( .D(blocktag_next[1]), .E(n1211), .CK(clk), .Q(
        \blocktag[1][1] ) );
  EDFFX1 \blocktag_reg[5][1]  ( .D(blocktag_next[1]), .E(n1135), .CK(clk), 
        .QN(n607) );
  EDFFX1 \blocktag_reg[1][18]  ( .D(blocktag_next[18]), .E(n1212), .CK(clk), 
        .QN(n591) );
  EDFFX1 \blocktag_reg[5][18]  ( .D(blocktag_next[18]), .E(n1136), .CK(clk), 
        .QN(n595) );
  EDFFX1 \blocktag_reg[1][12]  ( .D(blocktag_next[12]), .E(n1211), .CK(clk), 
        .Q(n254) );
  EDFFX1 \blocktag_reg[1][3]  ( .D(blocktag_next[3]), .E(n1211), .CK(clk), 
        .QN(n583) );
  EDFFX1 \blocktag_reg[5][12]  ( .D(blocktag_next[12]), .E(n1135), .CK(clk), 
        .Q(n250) );
  EDFFX1 \blocktag_reg[5][3]  ( .D(blocktag_next[3]), .E(n1135), .CK(clk), 
        .QN(n587) );
  EDFFX1 \blocktag_reg[1][17]  ( .D(blocktag_next[17]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][17] ) );
  EDFFX1 \blocktag_reg[5][17]  ( .D(blocktag_next[17]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][17] ) );
  EDFFX1 \blocktag_reg[1][5]  ( .D(blocktag_next[5]), .E(n1211), .CK(clk), 
        .QN(n575) );
  EDFFX1 \blocktag_reg[1][14]  ( .D(blocktag_next[14]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][14] ) );
  EDFFX1 \blocktag_reg[5][5]  ( .D(blocktag_next[5]), .E(n1135), .CK(clk), 
        .QN(n579) );
  EDFFX1 \blocktag_reg[1][22]  ( .D(blocktag_next[22]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][22] ) );
  EDFFX1 \blocktag_reg[5][14]  ( .D(blocktag_next[14]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][14] ) );
  EDFFX1 \blocktag_reg[5][22]  ( .D(blocktag_next[22]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][22] ) );
  EDFFX1 \blocktag_reg[1][16]  ( .D(blocktag_next[16]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][16] ) );
  EDFFX1 \blocktag_reg[5][16]  ( .D(blocktag_next[16]), .E(n1136), .CK(clk), 
        .Q(n246) );
  EDFFX1 \blocktag_reg[1][10]  ( .D(blocktag_next[10]), .E(n1211), .CK(clk), 
        .Q(\blocktag[1][10] ) );
  EDFFX1 \blocktag_reg[5][10]  ( .D(blocktag_next[10]), .E(n1135), .CK(clk), 
        .Q(\blocktag[5][10] ) );
  EDFFX1 \blocktag_reg[1][7]  ( .D(n3), .E(n1211), .CK(clk), .Q(n242) );
  EDFFX1 \blocktag_reg[5][7]  ( .D(n3), .E(n1135), .CK(clk), .Q(n238) );
  EDFFX1 \blocktag_reg[1][15]  ( .D(blocktag_next[15]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][15] ) );
  EDFFX1 \blocktag_reg[1][8]  ( .D(blocktag_next[8]), .E(n1211), .CK(clk), .Q(
        n234) );
  EDFFX1 \blocktag_reg[5][15]  ( .D(blocktag_next[15]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][15] ) );
  EDFFX1 \blocktag_reg[5][8]  ( .D(blocktag_next[8]), .E(n1135), .CK(clk), .Q(
        n230) );
  EDFFX1 \blocktag_reg[1][13]  ( .D(blocktag_next[13]), .E(n1212), .CK(clk), 
        .Q(\blocktag[1][13] ) );
  EDFFX1 \blocktag_reg[5][13]  ( .D(blocktag_next[13]), .E(n1136), .CK(clk), 
        .Q(\blocktag[5][13] ) );
  EDFFX1 \blocktag_reg[0][20]  ( .D(blocktag_next[20]), .E(n1231), .CK(clk), 
        .QN(n204) );
  EDFFX1 \blocktag_reg[4][20]  ( .D(blocktag_next[20]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][20] ) );
  EDFFX1 \blocktag_reg[0][19]  ( .D(blocktag_next[19]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][19] ) );
  EDFFX1 \blocktag_reg[0][0]  ( .D(n4), .E(n1230), .CK(clk), .Q(
        \blocktag[0][0] ) );
  EDFFX1 \blocktag_reg[4][19]  ( .D(blocktag_next[19]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][19] ) );
  EDFFX1 \blocktag_reg[4][0]  ( .D(n4), .E(n1154), .CK(clk), .Q(
        \blocktag[4][0] ) );
  EDFFX1 \blocktag_reg[0][23]  ( .D(blocktag_next[23]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][23] ) );
  EDFFX1 \blocktag_reg[0][24]  ( .D(blocktag_next[24]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][24] ) );
  EDFFX1 \blocktag_reg[4][23]  ( .D(blocktag_next[23]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][23] ) );
  EDFFX1 \blocktag_reg[4][24]  ( .D(blocktag_next[24]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][24] ) );
  EDFFX1 \blocktag_reg[0][2]  ( .D(blocktag_next[2]), .E(n1230), .CK(clk), .Q(
        \blocktag[0][2] ) );
  EDFFX1 \blocktag_reg[4][2]  ( .D(blocktag_next[2]), .E(n1154), .CK(clk), .Q(
        \blocktag[4][2] ) );
  EDFFX1 \blocktag_reg[0][11]  ( .D(blocktag_next[11]), .E(n1230), .CK(clk), 
        .Q(\blocktag[0][11] ) );
  EDFFX1 \blocktag_reg[4][11]  ( .D(blocktag_next[11]), .E(n1154), .CK(clk), 
        .Q(\blocktag[4][11] ) );
  EDFFX1 \blocktag_reg[0][1]  ( .D(blocktag_next[1]), .E(n1230), .CK(clk), .Q(
        \blocktag[0][1] ) );
  EDFFX1 \blocktag_reg[4][1]  ( .D(blocktag_next[1]), .E(n1154), .CK(clk), 
        .QN(n606) );
  EDFFX1 \blocktag_reg[0][18]  ( .D(blocktag_next[18]), .E(n1231), .CK(clk), 
        .QN(n590) );
  EDFFX1 \blocktag_reg[4][18]  ( .D(blocktag_next[18]), .E(n1155), .CK(clk), 
        .QN(n594) );
  EDFFX1 \blocktag_reg[0][12]  ( .D(blocktag_next[12]), .E(n1230), .CK(clk), 
        .Q(n253) );
  EDFFX1 \blocktag_reg[0][3]  ( .D(blocktag_next[3]), .E(n1230), .CK(clk), 
        .QN(n582) );
  EDFFX1 \blocktag_reg[4][12]  ( .D(blocktag_next[12]), .E(n1154), .CK(clk), 
        .Q(n249) );
  EDFFX1 \blocktag_reg[4][3]  ( .D(blocktag_next[3]), .E(n1154), .CK(clk), 
        .QN(n586) );
  EDFFX1 \blocktag_reg[0][17]  ( .D(blocktag_next[17]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][17] ) );
  EDFFX1 \blocktag_reg[4][17]  ( .D(blocktag_next[17]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][17] ) );
  EDFFX1 \blocktag_reg[0][5]  ( .D(blocktag_next[5]), .E(n1230), .CK(clk), 
        .QN(n574) );
  EDFFX1 \blocktag_reg[0][14]  ( .D(blocktag_next[14]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][14] ) );
  EDFFX1 \blocktag_reg[4][5]  ( .D(blocktag_next[5]), .E(n1154), .CK(clk), 
        .QN(n578) );
  EDFFX1 \blocktag_reg[0][22]  ( .D(blocktag_next[22]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][22] ) );
  EDFFX1 \blocktag_reg[4][14]  ( .D(blocktag_next[14]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][14] ) );
  EDFFX1 \blocktag_reg[4][22]  ( .D(blocktag_next[22]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][22] ) );
  EDFFX1 \blocktag_reg[0][16]  ( .D(blocktag_next[16]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][16] ) );
  EDFFX1 \blocktag_reg[4][16]  ( .D(blocktag_next[16]), .E(n1155), .CK(clk), 
        .Q(n245) );
  EDFFX1 \blocktag_reg[0][10]  ( .D(blocktag_next[10]), .E(n1230), .CK(clk), 
        .Q(\blocktag[0][10] ) );
  EDFFX1 \blocktag_reg[4][10]  ( .D(blocktag_next[10]), .E(n1154), .CK(clk), 
        .Q(\blocktag[4][10] ) );
  EDFFX1 \blocktag_reg[0][7]  ( .D(n3), .E(n1230), .CK(clk), .Q(n241) );
  EDFFX1 \blocktag_reg[4][7]  ( .D(n3), .E(n1154), .CK(clk), .Q(n237) );
  EDFFX1 \blocktag_reg[0][15]  ( .D(blocktag_next[15]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][15] ) );
  EDFFX1 \blocktag_reg[0][8]  ( .D(blocktag_next[8]), .E(n1230), .CK(clk), .Q(
        n233) );
  EDFFX1 \blocktag_reg[4][15]  ( .D(blocktag_next[15]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][15] ) );
  EDFFX1 \blocktag_reg[4][8]  ( .D(blocktag_next[8]), .E(n1154), .CK(clk), .Q(
        n229) );
  EDFFX1 \blocktag_reg[0][13]  ( .D(blocktag_next[13]), .E(n1231), .CK(clk), 
        .Q(\blocktag[0][13] ) );
  EDFFX1 \blocktag_reg[4][13]  ( .D(blocktag_next[13]), .E(n1155), .CK(clk), 
        .Q(\blocktag[4][13] ) );
  EDFFX1 \blocktag_reg[2][20]  ( .D(blocktag_next[20]), .E(n1193), .CK(clk), 
        .QN(n206) );
  EDFFX1 \blocktag_reg[6][20]  ( .D(blocktag_next[20]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][20] ) );
  EDFFX1 \blocktag_reg[2][19]  ( .D(blocktag_next[19]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][19] ) );
  EDFFX1 \blocktag_reg[2][0]  ( .D(n4), .E(n1192), .CK(clk), .Q(
        \blocktag[2][0] ) );
  EDFFX1 \blocktag_reg[6][19]  ( .D(blocktag_next[19]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][19] ) );
  EDFFX1 \blocktag_reg[6][0]  ( .D(n4), .E(n1115), .CK(clk), .Q(
        \blocktag[6][0] ) );
  EDFFX1 \blocktag_reg[2][23]  ( .D(blocktag_next[23]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][23] ) );
  EDFFX1 \blocktag_reg[2][24]  ( .D(blocktag_next[24]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][24] ) );
  EDFFX1 \blocktag_reg[6][23]  ( .D(blocktag_next[23]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][23] ) );
  EDFFX1 \blocktag_reg[6][24]  ( .D(blocktag_next[24]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][24] ) );
  EDFFX1 \blocktag_reg[2][2]  ( .D(blocktag_next[2]), .E(n1192), .CK(clk), .Q(
        \blocktag[2][2] ) );
  EDFFX1 \blocktag_reg[6][2]  ( .D(blocktag_next[2]), .E(n1115), .CK(clk), .Q(
        \blocktag[6][2] ) );
  EDFFX1 \blocktag_reg[2][11]  ( .D(blocktag_next[11]), .E(n1192), .CK(clk), 
        .Q(\blocktag[2][11] ) );
  EDFFX1 \blocktag_reg[6][11]  ( .D(blocktag_next[11]), .E(n1115), .CK(clk), 
        .Q(\blocktag[6][11] ) );
  EDFFX1 \blocktag_reg[2][1]  ( .D(blocktag_next[1]), .E(n1192), .CK(clk), .Q(
        \blocktag[2][1] ) );
  EDFFX1 \blocktag_reg[6][1]  ( .D(blocktag_next[1]), .E(n1115), .CK(clk), 
        .QN(n608) );
  EDFFX1 \blocktag_reg[2][18]  ( .D(blocktag_next[18]), .E(n1193), .CK(clk), 
        .QN(n592) );
  EDFFX1 \blocktag_reg[6][18]  ( .D(blocktag_next[18]), .E(n1116), .CK(clk), 
        .QN(n596) );
  EDFFX1 \blocktag_reg[2][12]  ( .D(blocktag_next[12]), .E(n1192), .CK(clk), 
        .Q(n255) );
  EDFFX1 \blocktag_reg[2][3]  ( .D(blocktag_next[3]), .E(n1192), .CK(clk), 
        .QN(n584) );
  EDFFX1 \blocktag_reg[6][12]  ( .D(blocktag_next[12]), .E(n1115), .CK(clk), 
        .Q(n251) );
  EDFFX1 \blocktag_reg[6][3]  ( .D(blocktag_next[3]), .E(n1115), .CK(clk), 
        .QN(n588) );
  EDFFX1 \blocktag_reg[2][17]  ( .D(blocktag_next[17]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][17] ) );
  EDFFX1 \blocktag_reg[6][17]  ( .D(blocktag_next[17]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][17] ) );
  EDFFX1 \blocktag_reg[2][5]  ( .D(blocktag_next[5]), .E(n1192), .CK(clk), 
        .QN(n576) );
  EDFFX1 \blocktag_reg[2][14]  ( .D(blocktag_next[14]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][14] ) );
  EDFFX1 \blocktag_reg[6][5]  ( .D(blocktag_next[5]), .E(n1115), .CK(clk), 
        .QN(n580) );
  EDFFX1 \blocktag_reg[2][22]  ( .D(blocktag_next[22]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][22] ) );
  EDFFX1 \blocktag_reg[6][14]  ( .D(blocktag_next[14]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][14] ) );
  EDFFX1 \blocktag_reg[6][22]  ( .D(blocktag_next[22]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][22] ) );
  EDFFX1 \blocktag_reg[2][16]  ( .D(blocktag_next[16]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][16] ) );
  EDFFX1 \blocktag_reg[6][16]  ( .D(blocktag_next[16]), .E(n1116), .CK(clk), 
        .Q(n247) );
  EDFFX1 \blocktag_reg[2][10]  ( .D(blocktag_next[10]), .E(n1192), .CK(clk), 
        .Q(\blocktag[2][10] ) );
  EDFFX1 \blocktag_reg[6][10]  ( .D(blocktag_next[10]), .E(n1115), .CK(clk), 
        .Q(\blocktag[6][10] ) );
  EDFFX1 \blocktag_reg[2][7]  ( .D(n3), .E(n1192), .CK(clk), .Q(n243) );
  EDFFX1 \blocktag_reg[6][7]  ( .D(n3), .E(n1115), .CK(clk), .Q(n239) );
  EDFFX1 \blocktag_reg[2][15]  ( .D(blocktag_next[15]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][15] ) );
  EDFFX1 \blocktag_reg[2][8]  ( .D(blocktag_next[8]), .E(n1192), .CK(clk), .Q(
        n235) );
  EDFFX1 \blocktag_reg[6][15]  ( .D(blocktag_next[15]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][15] ) );
  EDFFX1 \blocktag_reg[6][8]  ( .D(blocktag_next[8]), .E(n1115), .CK(clk), .Q(
        n231) );
  EDFFX1 \blocktag_reg[2][13]  ( .D(blocktag_next[13]), .E(n1193), .CK(clk), 
        .Q(\blocktag[2][13] ) );
  EDFFX1 \blocktag_reg[6][13]  ( .D(blocktag_next[13]), .E(n1116), .CK(clk), 
        .Q(\blocktag[6][13] ) );
  EDFFX1 \blocktag_reg[6][9]  ( .D(blocktag_next[9]), .E(n1115), .CK(clk), .Q(
        \blocktag[6][9] ) );
  EDFFX1 \blocktag_reg[2][9]  ( .D(blocktag_next[9]), .E(n1192), .CK(clk), .Q(
        \blocktag[2][9] ) );
  EDFFX1 \blocktag_reg[5][9]  ( .D(blocktag_next[9]), .E(n1135), .CK(clk), .Q(
        \blocktag[5][9] ) );
  EDFFX1 \blocktag_reg[1][9]  ( .D(blocktag_next[9]), .E(n1211), .CK(clk), .Q(
        \blocktag[1][9] ) );
  EDFFX1 \blocktag_reg[7][9]  ( .D(blocktag_next[9]), .E(n1100), .CK(clk), .Q(
        \blocktag[7][9] ) );
  EDFFX1 \blocktag_reg[3][9]  ( .D(blocktag_next[9]), .E(n1173), .CK(clk), .Q(
        \blocktag[3][9] ) );
  EDFFX1 \blocktag_reg[5][4]  ( .D(blocktag_next[4]), .E(n1135), .CK(clk), .Q(
        \blocktag[5][4] ) );
  EDFFX1 \blocktag_reg[1][4]  ( .D(blocktag_next[4]), .E(n1211), .CK(clk), .Q(
        \blocktag[1][4] ) );
  EDFFX1 \blocktag_reg[4][4]  ( .D(blocktag_next[4]), .E(n1154), .CK(clk), .Q(
        \blocktag[4][4] ) );
  EDFFX1 \blocktag_reg[0][4]  ( .D(blocktag_next[4]), .E(n1230), .CK(clk), .Q(
        \blocktag[0][4] ) );
  EDFFX1 \blocktag_reg[4][9]  ( .D(blocktag_next[9]), .E(n1154), .CK(clk), .Q(
        \blocktag[4][9] ) );
  EDFFX1 \blocktag_reg[0][9]  ( .D(blocktag_next[9]), .E(n1230), .CK(clk), .Q(
        \blocktag[0][9] ) );
  EDFFX1 \blocktag_reg[6][4]  ( .D(blocktag_next[4]), .E(n1115), .CK(clk), .Q(
        \blocktag[6][4] ) );
  EDFFX1 \blocktag_reg[2][4]  ( .D(blocktag_next[4]), .E(n1192), .CK(clk), .Q(
        \blocktag[2][4] ) );
  EDFFX1 \blocktag_reg[7][4]  ( .D(blocktag_next[4]), .E(n1100), .CK(clk), .Q(
        \blocktag[7][4] ) );
  EDFFX1 \blocktag_reg[3][4]  ( .D(blocktag_next[4]), .E(n1173), .CK(clk), .Q(
        \blocktag[3][4] ) );
  EDFFX1 \blocktag_reg[3][21]  ( .D(blocktag_next[21]), .E(n1174), .CK(clk), 
        .Q(\blocktag[3][21] ) );
  EDFFX1 \blocktag_reg[5][6]  ( .D(blocktag_next[6]), .E(n1135), .CK(clk), 
        .QN(n262) );
  EDFFX1 \blocktag_reg[1][6]  ( .D(blocktag_next[6]), .E(n1211), .CK(clk), 
        .QN(n258) );
  EDFFX1 \blocktag_reg[4][6]  ( .D(blocktag_next[6]), .E(n1154), .CK(clk), 
        .QN(n261) );
  EDFFX1 \blocktag_reg[0][6]  ( .D(blocktag_next[6]), .E(n1230), .CK(clk), 
        .QN(n257) );
  EDFFX1 \blocktag_reg[6][6]  ( .D(blocktag_next[6]), .E(n1115), .CK(clk), 
        .QN(n263) );
  EDFFX1 \blocktag_reg[2][6]  ( .D(blocktag_next[6]), .E(n1192), .CK(clk), 
        .QN(n259) );
  EDFFX1 \blocktag_reg[7][6]  ( .D(blocktag_next[6]), .E(n1100), .CK(clk), 
        .QN(n264) );
  EDFFX1 \blocktag_reg[3][6]  ( .D(blocktag_next[6]), .E(n1173), .CK(clk), 
        .QN(n260) );
  EDFFXL \blocktag_reg[7][21]  ( .D(blocktag_next[21]), .E(n1101), .CK(clk), 
        .QN(n605) );
  EDFFXL \blocktag_reg[6][21]  ( .D(blocktag_next[21]), .E(n1116), .CK(clk), 
        .QN(n604) );
  EDFFXL \blocktag_reg[5][21]  ( .D(blocktag_next[21]), .E(n1136), .CK(clk), 
        .QN(n603) );
  EDFFXL \blocktag_reg[4][21]  ( .D(blocktag_next[21]), .E(n1155), .CK(clk), 
        .QN(n602) );
  DFFSRXL \blockvalid_reg[2]  ( .D(n1721), .CK(clk), .SN(1'b1), .RN(n1260), 
        .Q(blockvalid[2]), .QN(n1737) );
  DFFSRX4 \blockvalid_reg[3]  ( .D(n1720), .CK(clk), .SN(1'b1), .RN(n1260), 
        .Q(blockvalid[3]), .QN(n1736) );
  DFFSRX4 \blockvalid_reg[1]  ( .D(n1722), .CK(clk), .SN(1'b1), .RN(n1260), 
        .Q(blockvalid[1]), .QN(n1738) );
  DFFSRX4 \blockvalid_reg[4]  ( .D(n1719), .CK(clk), .SN(1'b1), .RN(n1260), 
        .QN(n1735) );
  DFFSRX4 \blockvalid_reg[5]  ( .D(n1718), .CK(clk), .SN(1'b1), .RN(n1260), 
        .QN(n1734) );
  DFFSRX4 \blockvalid_reg[7]  ( .D(n1716), .CK(clk), .SN(1'b1), .RN(n1260), 
        .QN(n1732) );
  XOR2X2 U3 ( .A(n1515), .B(proc_addr[15]), .Y(n1278) );
  NAND4X4 U4 ( .A(n1280), .B(n1279), .C(n1278), .D(n1277), .Y(n1284) );
  NAND2X6 U5 ( .A(tag[16]), .B(proc_addr[21]), .Y(n223) );
  BUFX20 U6 ( .A(n963), .Y(n978) );
  BUFX4 U7 ( .A(n1752), .Y(mem_read) );
  CLKINVX8 U8 ( .A(n1500), .Y(n214) );
  NAND4X4 U9 ( .A(n1272), .B(n1271), .C(n1270), .D(n1269), .Y(n1276) );
  INVX8 U10 ( .A(n1541), .Y(n1299) );
  BUFX6 U11 ( .A(n1), .Y(n1067) );
  MX4X2 U12 ( .A(\blocktag[0][24] ), .B(\blocktag[1][24] ), .C(
        \blocktag[2][24] ), .D(\blocktag[3][24] ), .S0(n1044), .S1(n1011), .Y(
        n610) );
  MX4X2 U13 ( .A(\blocktag[4][24] ), .B(\blocktag[5][24] ), .C(
        \blocktag[6][24] ), .D(\blocktag[7][24] ), .S0(n1044), .S1(n1011), .Y(
        n611) );
  INVX3 U14 ( .A(blockdata[3]), .Y(n1571) );
  AO22X1 U15 ( .A0(proc_addr[12]), .A1(mem_read), .B0(tag[7]), .B1(mem_write), 
        .Y(n1771) );
  AO22X1 U16 ( .A0(proc_addr[14]), .A1(mem_read), .B0(tag[9]), .B1(mem_write), 
        .Y(n1769) );
  AO22X1 U17 ( .A0(proc_addr[16]), .A1(mem_read), .B0(tag[11]), .B1(mem_write), 
        .Y(n1767) );
  AO22X1 U18 ( .A0(proc_addr[17]), .A1(mem_read), .B0(tag[12]), .B1(mem_write), 
        .Y(n1766) );
  MXI2X4 U19 ( .A(n1522), .B(n1521), .S0(n1068), .Y(n3) );
  INVX1 U20 ( .A(tag[7]), .Y(n1522) );
  NAND4X6 U21 ( .A(n1296), .B(n1295), .C(n1294), .D(n1293), .Y(n1541) );
  NOR2X6 U22 ( .A(n1284), .B(n1283), .Y(n1294) );
  NOR2X4 U23 ( .A(n1276), .B(n1275), .Y(n1295) );
  AND2X4 U24 ( .A(n1337), .B(n1336), .Y(n568) );
  INVX6 U25 ( .A(n1551), .Y(n1548) );
  INVX6 U26 ( .A(n2), .Y(n1485) );
  CLKAND2X3 U27 ( .A(n1255), .B(blockdata[8]), .Y(n1849) );
  CLKAND2X3 U28 ( .A(n1255), .B(blockdata[16]), .Y(n1842) );
  CLKAND2X3 U29 ( .A(n1255), .B(blockdata[17]), .Y(n1841) );
  CLKAND2X3 U30 ( .A(n1255), .B(blockdata[18]), .Y(n1840) );
  CLKAND2X3 U31 ( .A(n1255), .B(blockdata[19]), .Y(n1839) );
  CLKAND2X3 U32 ( .A(n1255), .B(blockdata[20]), .Y(n1838) );
  CLKAND2X3 U33 ( .A(n1255), .B(blockdata[21]), .Y(n1837) );
  CLKAND2X3 U34 ( .A(n1255), .B(blockdata[22]), .Y(n1836) );
  CLKAND2X3 U35 ( .A(n1255), .B(blockdata[23]), .Y(n1835) );
  CLKAND2X3 U36 ( .A(n1255), .B(blockdata[24]), .Y(n1834) );
  CLKAND2X3 U37 ( .A(n1255), .B(blockdata[25]), .Y(n1833) );
  CLKAND2X3 U38 ( .A(n1255), .B(blockdata[32]), .Y(n1828) );
  CLKAND2X3 U39 ( .A(n1254), .B(blockdata[48]), .Y(n1813) );
  CLKAND2X3 U40 ( .A(n1254), .B(blockdata[49]), .Y(n1812) );
  CLKAND2X3 U41 ( .A(n1254), .B(blockdata[50]), .Y(n1811) );
  CLKAND2X3 U42 ( .A(n1254), .B(blockdata[51]), .Y(n1810) );
  CLKAND2X3 U43 ( .A(n1254), .B(blockdata[52]), .Y(n1809) );
  CLKAND2X3 U44 ( .A(n1254), .B(blockdata[53]), .Y(n1808) );
  CLKAND2X3 U45 ( .A(n1254), .B(blockdata[54]), .Y(n1807) );
  CLKAND2X3 U46 ( .A(n1254), .B(blockdata[55]), .Y(n1806) );
  CLKAND2X3 U47 ( .A(n1254), .B(blockdata[56]), .Y(n1805) );
  CLKAND2X3 U48 ( .A(n1254), .B(blockdata[57]), .Y(n1804) );
  CLKAND2X3 U49 ( .A(n1254), .B(blockdata[64]), .Y(n1799) );
  CLKAND2X3 U50 ( .A(n1254), .B(blockdata[65]), .Y(n1798) );
  CLKAND2X3 U51 ( .A(n1254), .B(blockdata[66]), .Y(n1797) );
  CLKAND2X3 U52 ( .A(n1254), .B(blockdata[67]), .Y(n1796) );
  CLKAND2X3 U53 ( .A(n1254), .B(blockdata[68]), .Y(n1795) );
  CLKAND2X3 U54 ( .A(n1254), .B(blockdata[80]), .Y(n1783) );
  CLKAND2X3 U55 ( .A(n1254), .B(blockdata[81]), .Y(n1782) );
  CLKAND2X3 U56 ( .A(n1254), .B(blockdata[82]), .Y(n1781) );
  AO22X1 U57 ( .A0(proc_addr[5]), .A1(mem_read), .B0(tag[0]), .B1(mem_write), 
        .Y(n1778) );
  AO22X1 U58 ( .A0(proc_addr[7]), .A1(mem_read), .B0(tag[2]), .B1(mem_write), 
        .Y(n1776) );
  AO22X1 U59 ( .A0(proc_addr[8]), .A1(mem_read), .B0(tag[3]), .B1(mem_write), 
        .Y(n1775) );
  AO22X1 U60 ( .A0(proc_addr[9]), .A1(mem_read), .B0(tag[4]), .B1(mem_write), 
        .Y(n1774) );
  AO22X1 U61 ( .A0(proc_addr[11]), .A1(mem_read), .B0(tag[6]), .B1(mem_write), 
        .Y(n1772) );
  AO22X1 U62 ( .A0(proc_addr[13]), .A1(mem_read), .B0(tag[8]), .B1(mem_write), 
        .Y(n1770) );
  AO22X1 U63 ( .A0(proc_addr[15]), .A1(mem_read), .B0(tag[10]), .B1(mem_write), 
        .Y(n1768) );
  AO22X1 U64 ( .A0(proc_addr[18]), .A1(mem_read), .B0(tag[13]), .B1(mem_write), 
        .Y(n1765) );
  AO22X1 U65 ( .A0(proc_addr[20]), .A1(mem_read), .B0(tag[15]), .B1(mem_write), 
        .Y(n1763) );
  AO22X1 U66 ( .A0(proc_addr[22]), .A1(mem_read), .B0(tag[17]), .B1(mem_write), 
        .Y(n1761) );
  AO22X1 U67 ( .A0(proc_addr[23]), .A1(mem_read), .B0(tag[18]), .B1(mem_write), 
        .Y(n1760) );
  AO22X1 U68 ( .A0(proc_addr[24]), .A1(mem_read), .B0(tag[19]), .B1(mem_write), 
        .Y(n1759) );
  AO22X1 U69 ( .A0(proc_addr[25]), .A1(mem_read), .B0(tag[20]), .B1(mem_write), 
        .Y(n1758) );
  AO22X1 U70 ( .A0(proc_addr[27]), .A1(mem_read), .B0(tag[22]), .B1(mem_write), 
        .Y(n1756) );
  AO22X1 U71 ( .A0(proc_addr[28]), .A1(mem_read), .B0(tag[23]), .B1(mem_write), 
        .Y(n1755) );
  CLKINVX2 U72 ( .A(tag[22]), .Y(n1482) );
  CLKINVX3 U73 ( .A(tag[24]), .Y(n1476) );
  MXI2X4 U74 ( .A(n1536), .B(n1535), .S0(n1068), .Y(n4) );
  INVXL U75 ( .A(tag[0]), .Y(n1536) );
  CLKINVX3 U76 ( .A(tag[19]), .Y(n1491) );
  NAND2XL U77 ( .A(mem_rdata[91]), .B(n1074), .Y(n1343) );
  NAND2XL U78 ( .A(mem_rdata[90]), .B(n1074), .Y(n1344) );
  NAND2X2 U79 ( .A(mem_rdata[3]), .B(n1070), .Y(n1462) );
  BUFX2 U80 ( .A(n982), .Y(n990) );
  BUFX8 U81 ( .A(N32), .Y(n984) );
  BUFX2 U82 ( .A(n1019), .Y(n1023) );
  BUFX8 U83 ( .A(N31), .Y(n1048) );
  INVX2 U84 ( .A(N32), .Y(n1247) );
  BUFX2 U85 ( .A(n1048), .Y(n1016) );
  BUFX2 U86 ( .A(n1015), .Y(n1024) );
  AND2XL U87 ( .A(n739), .B(proc_stall), .Y(n1) );
  INVX16 U88 ( .A(N31), .Y(n1246) );
  CLKINVX3 U89 ( .A(n1062), .Y(n1061) );
  CLKINVX3 U90 ( .A(n1062), .Y(n1060) );
  BUFX2 U91 ( .A(n1014), .Y(n981) );
  BUFX8 U92 ( .A(n1067), .Y(n1079) );
  CLKINVX8 U93 ( .A(n210), .Y(tag[16]) );
  CLKBUFX8 U94 ( .A(n985), .Y(n982) );
  BUFX2 U95 ( .A(n984), .Y(n987) );
  CLKBUFX3 U96 ( .A(n560), .Y(n1131) );
  AND2X6 U97 ( .A(n212), .B(n213), .Y(n2) );
  BUFX2 U98 ( .A(n1017), .Y(n1020) );
  AND2X6 U99 ( .A(n558), .B(n1405), .Y(n553) );
  BUFX16 U100 ( .A(n553), .Y(n1064) );
  BUFX16 U101 ( .A(n553), .Y(n1063) );
  AND2X4 U102 ( .A(n558), .B(n1066), .Y(n559) );
  BUFX12 U103 ( .A(n559), .Y(n1059) );
  BUFX12 U104 ( .A(n559), .Y(n1058) );
  BUFX2 U105 ( .A(n1248), .Y(n966) );
  INVX3 U106 ( .A(proc_addr[21]), .Y(n221) );
  BUFX20 U107 ( .A(n1080), .Y(n1070) );
  BUFX20 U108 ( .A(n1067), .Y(n1080) );
  OAI221X4 U109 ( .A0(n1059), .A1(n1562), .B0(n1465), .B1(n1060), .C0(n1402), 
        .Y(block_next[34]) );
  NAND2X4 U110 ( .A(mem_rdata[48]), .B(n1072), .Y(n1388) );
  NAND2X4 U111 ( .A(mem_rdata[49]), .B(n1072), .Y(n1387) );
  NAND2X4 U112 ( .A(mem_rdata[50]), .B(n1072), .Y(n1386) );
  NAND2X4 U113 ( .A(mem_rdata[51]), .B(n1072), .Y(n1385) );
  NAND2X4 U114 ( .A(mem_rdata[52]), .B(n1072), .Y(n1384) );
  NAND2X4 U115 ( .A(mem_rdata[40]), .B(n1072), .Y(n1396) );
  NAND2X4 U116 ( .A(mem_rdata[46]), .B(n1072), .Y(n1390) );
  BUFX20 U117 ( .A(n1070), .Y(n1072) );
  NAND2X4 U118 ( .A(mem_rdata[66]), .B(n1073), .Y(n1368) );
  NAND2X4 U119 ( .A(mem_rdata[67]), .B(n1073), .Y(n1367) );
  NAND2X4 U120 ( .A(mem_rdata[68]), .B(n1073), .Y(n1366) );
  NAND2X4 U121 ( .A(mem_rdata[71]), .B(n1073), .Y(n1363) );
  NAND2X4 U122 ( .A(mem_rdata[69]), .B(n1073), .Y(n1365) );
  NAND2X4 U123 ( .A(mem_rdata[72]), .B(n1073), .Y(n1362) );
  NAND2X4 U124 ( .A(mem_rdata[73]), .B(n1073), .Y(n1361) );
  BUFX20 U125 ( .A(n1070), .Y(n1073) );
  BUFX20 U126 ( .A(n1079), .Y(n1075) );
  OAI221X4 U127 ( .A0(n1054), .A1(n1673), .B0(n1421), .B1(n1057), .C0(n1346), 
        .Y(block_next[88]) );
  OAI221X4 U128 ( .A0(n1054), .A1(n1668), .B0(n1423), .B1(n1057), .C0(n1347), 
        .Y(block_next[87]) );
  OAI221X4 U129 ( .A0(n1054), .A1(n1678), .B0(n1419), .B1(n1057), .C0(n1345), 
        .Y(block_next[89]) );
  OAI221X4 U130 ( .A0(n1055), .A1(n1628), .B0(n1439), .B1(n1372), .C0(n1355), 
        .Y(block_next[79]) );
  OAI221X4 U131 ( .A0(n1055), .A1(n1633), .B0(n1437), .B1(n1057), .C0(n1354), 
        .Y(block_next[80]) );
  OAI221X4 U132 ( .A0(n1054), .A1(n1683), .B0(n1417), .B1(n1057), .C0(n1344), 
        .Y(block_next[90]) );
  OAI221X4 U133 ( .A0(n1054), .A1(n1663), .B0(n1425), .B1(n1056), .C0(n1348), 
        .Y(block_next[86]) );
  OAI221X4 U134 ( .A0(n1054), .A1(n1658), .B0(n1427), .B1(n1057), .C0(n1349), 
        .Y(block_next[85]) );
  OAI221X4 U135 ( .A0(n1054), .A1(n1653), .B0(n1429), .B1(n1056), .C0(n1350), 
        .Y(block_next[84]) );
  OAI221X4 U136 ( .A0(n1055), .A1(n1648), .B0(n1431), .B1(n1056), .C0(n1351), 
        .Y(block_next[83]) );
  OAI221X4 U137 ( .A0(n1055), .A1(n1643), .B0(n1433), .B1(n1057), .C0(n1352), 
        .Y(block_next[82]) );
  OAI221X4 U138 ( .A0(n1055), .A1(n1638), .B0(n1435), .B1(n1056), .C0(n1353), 
        .Y(block_next[81]) );
  OAI221X4 U139 ( .A0(n1054), .A1(n1688), .B0(n1415), .B1(n1057), .C0(n1343), 
        .Y(block_next[91]) );
  BUFX20 U140 ( .A(n1371), .Y(n1054) );
  OAI221X4 U141 ( .A0(n1051), .A1(n1580), .B0(n1459), .B1(n1052), .C0(n1330), 
        .Y(block_next[101]) );
  OAI221X4 U142 ( .A0(n1051), .A1(n1590), .B0(n1455), .B1(n1053), .C0(n1328), 
        .Y(block_next[103]) );
  OAI221X4 U143 ( .A0(n1051), .A1(n1595), .B0(n1453), .B1(n1053), .C0(n1327), 
        .Y(block_next[104]) );
  BUFX20 U144 ( .A(n569), .Y(n1051) );
  OAI221X4 U145 ( .A0(n1066), .A1(n1435), .B0(n1064), .B1(n1641), .C0(n1434), 
        .Y(block_next[17]) );
  OAI221X4 U146 ( .A0(n1065), .A1(n1463), .B0(n1064), .B1(n1571), .C0(n1462), 
        .Y(block_next[3]) );
  OAI221X4 U147 ( .A0(n1066), .A1(n1429), .B0(n1063), .B1(n1656), .C0(n1428), 
        .Y(block_next[20]) );
  OAI221X4 U148 ( .A0(n1066), .A1(n1431), .B0(n1064), .B1(n1651), .C0(n1430), 
        .Y(block_next[19]) );
  OAI221X4 U149 ( .A0(n1066), .A1(n1443), .B0(n1063), .B1(n1621), .C0(n1442), 
        .Y(block_next[13]) );
  OAI221X4 U150 ( .A0(n1065), .A1(n1451), .B0(n1064), .B1(n1601), .C0(n1450), 
        .Y(block_next[9]) );
  OAI221X4 U151 ( .A0(n1066), .A1(n1419), .B0(n1063), .B1(n1681), .C0(n1418), 
        .Y(block_next[25]) );
  OAI221X4 U152 ( .A0(n1066), .A1(n1421), .B0(n1063), .B1(n1676), .C0(n1420), 
        .Y(block_next[24]) );
  OAI221X4 U153 ( .A0(n1066), .A1(n1423), .B0(n1063), .B1(n1671), .C0(n1422), 
        .Y(block_next[23]) );
  OAI221X4 U154 ( .A0(n1066), .A1(n1425), .B0(n1063), .B1(n1666), .C0(n1424), 
        .Y(block_next[22]) );
  OAI221X4 U155 ( .A0(n1065), .A1(n1449), .B0(n1063), .B1(n1606), .C0(n1448), 
        .Y(block_next[10]) );
  OAI221X4 U156 ( .A0(n1065), .A1(n1445), .B0(n1064), .B1(n1616), .C0(n1444), 
        .Y(block_next[12]) );
  OAI221X4 U157 ( .A0(n1065), .A1(n1459), .B0(n1064), .B1(n1581), .C0(n1458), 
        .Y(block_next[5]) );
  OAI221X4 U158 ( .A0(n1066), .A1(n1427), .B0(n1063), .B1(n1661), .C0(n1426), 
        .Y(block_next[21]) );
  OAI221X4 U159 ( .A0(n1066), .A1(n1439), .B0(n1064), .B1(n1631), .C0(n1438), 
        .Y(block_next[15]) );
  OAI221X4 U160 ( .A0(n1065), .A1(n1447), .B0(n553), .B1(n1611), .C0(n1446), 
        .Y(block_next[11]) );
  OAI221X4 U161 ( .A0(n1065), .A1(n1457), .B0(n1064), .B1(n1586), .C0(n1456), 
        .Y(block_next[6]) );
  OAI221X4 U162 ( .A0(n1065), .A1(n1455), .B0(n1064), .B1(n1591), .C0(n1454), 
        .Y(block_next[7]) );
  OAI221X4 U163 ( .A0(n1066), .A1(n1433), .B0(n1064), .B1(n1646), .C0(n1432), 
        .Y(block_next[18]) );
  OAI221X4 U164 ( .A0(n1066), .A1(n1437), .B0(n1064), .B1(n1636), .C0(n1436), 
        .Y(block_next[16]) );
  OAI221X4 U165 ( .A0(n1065), .A1(n1461), .B0(n1064), .B1(n1576), .C0(n1460), 
        .Y(block_next[4]) );
  OAI221X4 U166 ( .A0(n1065), .A1(n1465), .B0(n1064), .B1(n1566), .C0(n1464), 
        .Y(block_next[2]) );
  OAI221X4 U167 ( .A0(n1065), .A1(n1467), .B0(n1064), .B1(n1561), .C0(n1466), 
        .Y(block_next[1]) );
  OAI221X4 U168 ( .A0(n1066), .A1(n1441), .B0(n1064), .B1(n1626), .C0(n1440), 
        .Y(block_next[14]) );
  OAI221X4 U169 ( .A0(n1066), .A1(n1417), .B0(n1063), .B1(n1686), .C0(n1416), 
        .Y(block_next[26]) );
  OAI221X4 U170 ( .A0(n1065), .A1(n1453), .B0(n1064), .B1(n1596), .C0(n1452), 
        .Y(block_next[8]) );
  BUFX20 U171 ( .A(n1078), .Y(n1077) );
  CLKBUFX4 U172 ( .A(n1067), .Y(n1078) );
  NAND2X4 U173 ( .A(mem_rdata[122]), .B(n1077), .Y(n1309) );
  OAI221X4 U174 ( .A0(n1050), .A1(n1665), .B0(n1425), .B1(n1052), .C0(n1313), 
        .Y(block_next[118]) );
  OAI221X4 U175 ( .A0(n1050), .A1(n1680), .B0(n1419), .B1(n1052), .C0(n1310), 
        .Y(block_next[121]) );
  OAI221X4 U176 ( .A0(n1050), .A1(n1675), .B0(n1421), .B1(n1052), .C0(n1311), 
        .Y(block_next[120]) );
  OAI221X4 U177 ( .A0(n1050), .A1(n1670), .B0(n1423), .B1(n1052), .C0(n1312), 
        .Y(block_next[119]) );
  OAI221X4 U178 ( .A0(n1050), .A1(n1685), .B0(n1417), .B1(n1052), .C0(n1309), 
        .Y(block_next[122]) );
  OAI221X4 U179 ( .A0(n1050), .A1(n1712), .B0(n1407), .B1(n1052), .C0(n1304), 
        .Y(block_next[127]) );
  NAND2X4 U180 ( .A(mem_rdata[127]), .B(n1077), .Y(n1304) );
  OAI221X4 U181 ( .A0(n1050), .A1(n1695), .B0(n1413), .B1(n1052), .C0(n1307), 
        .Y(block_next[124]) );
  NAND2X4 U182 ( .A(mem_rdata[124]), .B(n1077), .Y(n1307) );
  OAI221X4 U183 ( .A0(n1050), .A1(n1690), .B0(n1415), .B1(n1052), .C0(n1308), 
        .Y(block_next[123]) );
  NAND2X4 U184 ( .A(mem_rdata[123]), .B(n1077), .Y(n1308) );
  OAI221X4 U185 ( .A0(n1050), .A1(n1705), .B0(n1409), .B1(n1052), .C0(n1305), 
        .Y(block_next[126]) );
  NAND2X4 U186 ( .A(mem_rdata[126]), .B(n1077), .Y(n1305) );
  OAI221X4 U187 ( .A0(n1050), .A1(n1700), .B0(n1411), .B1(n1052), .C0(n1306), 
        .Y(block_next[125]) );
  BUFX20 U188 ( .A(n569), .Y(n1050) );
  NAND2X4 U189 ( .A(mem_rdata[125]), .B(n1077), .Y(n1306) );
  OAI221X4 U190 ( .A0(n1059), .A1(n1602), .B0(n1449), .B1(n1060), .C0(n1394), 
        .Y(block_next[42]) );
  OAI221X4 U191 ( .A0(n1059), .A1(n1622), .B0(n1441), .B1(n1061), .C0(n1390), 
        .Y(block_next[46]) );
  OAI221X4 U192 ( .A0(n1059), .A1(n1632), .B0(n1437), .B1(n1061), .C0(n1388), 
        .Y(block_next[48]) );
  OAI221X4 U193 ( .A0(n1059), .A1(n1642), .B0(n1433), .B1(n1061), .C0(n1386), 
        .Y(block_next[50]) );
  OAI221X4 U194 ( .A0(n1059), .A1(n1637), .B0(n1435), .B1(n1061), .C0(n1387), 
        .Y(block_next[49]) );
  OAI221X4 U195 ( .A0(n1059), .A1(n1607), .B0(n1447), .B1(n1060), .C0(n1393), 
        .Y(block_next[43]) );
  OAI221X4 U196 ( .A0(n1059), .A1(n1617), .B0(n1443), .B1(n1061), .C0(n1391), 
        .Y(block_next[45]) );
  OAI221X4 U197 ( .A0(n1059), .A1(n1597), .B0(n1451), .B1(n1060), .C0(n1395), 
        .Y(block_next[41]) );
  OAI221X4 U198 ( .A0(n1059), .A1(n1592), .B0(n1453), .B1(n1060), .C0(n1396), 
        .Y(block_next[40]) );
  OAI221X4 U199 ( .A0(n1059), .A1(n1647), .B0(n1431), .B1(n1061), .C0(n1385), 
        .Y(block_next[51]) );
  OAI221X4 U200 ( .A0(n1058), .A1(n1652), .B0(n1429), .B1(n1061), .C0(n1384), 
        .Y(block_next[52]) );
  OAI221X4 U201 ( .A0(n1059), .A1(n1612), .B0(n1445), .B1(n1060), .C0(n1392), 
        .Y(block_next[44]) );
  OAI221X4 U202 ( .A0(n1058), .A1(n1687), .B0(n1415), .B1(n1405), .C0(n1377), 
        .Y(block_next[59]) );
  NAND2X4 U203 ( .A(mem_rdata[59]), .B(n1077), .Y(n1377) );
  OAI221X4 U204 ( .A0(n1055), .A1(n1558), .B0(n1467), .B1(n1056), .C0(n1369), 
        .Y(block_next[65]) );
  OAI221X4 U205 ( .A0(n1058), .A1(n1702), .B0(n1409), .B1(n1060), .C0(n1374), 
        .Y(block_next[62]) );
  NAND2X4 U206 ( .A(mem_rdata[62]), .B(n1077), .Y(n1374) );
  OAI221X4 U207 ( .A0(n1058), .A1(n1697), .B0(n1411), .B1(n1060), .C0(n1375), 
        .Y(block_next[61]) );
  NAND2X4 U208 ( .A(mem_rdata[61]), .B(n1077), .Y(n1375) );
  OAI221X4 U209 ( .A0(n1058), .A1(n1677), .B0(n1419), .B1(n1060), .C0(n1379), 
        .Y(block_next[57]) );
  OAI221X4 U210 ( .A0(n1058), .A1(n1682), .B0(n1417), .B1(n1061), .C0(n1378), 
        .Y(block_next[58]) );
  OAI221X4 U211 ( .A0(n1058), .A1(n1657), .B0(n1427), .B1(n1061), .C0(n1383), 
        .Y(block_next[53]) );
  OAI221X4 U212 ( .A0(n1058), .A1(n1667), .B0(n1423), .B1(n1061), .C0(n1381), 
        .Y(block_next[55]) );
  OAI221X4 U213 ( .A0(n1058), .A1(n1662), .B0(n1425), .B1(n1061), .C0(n1382), 
        .Y(block_next[54]) );
  OAI221X4 U214 ( .A0(n1055), .A1(n1603), .B0(n1449), .B1(n1056), .C0(n1360), 
        .Y(block_next[74]) );
  OAI221X4 U215 ( .A0(n1055), .A1(n1623), .B0(n1441), .B1(n1057), .C0(n1356), 
        .Y(block_next[78]) );
  OAI221X4 U216 ( .A0(n1055), .A1(n1608), .B0(n1447), .B1(n1056), .C0(n1359), 
        .Y(block_next[75]) );
  OAI221X4 U217 ( .A0(n1055), .A1(n1618), .B0(n1443), .B1(n1056), .C0(n1357), 
        .Y(block_next[77]) );
  OAI221X4 U218 ( .A0(n1055), .A1(n1593), .B0(n1453), .B1(n1056), .C0(n1362), 
        .Y(block_next[72]) );
  OAI221X4 U219 ( .A0(n1054), .A1(n1588), .B0(n1455), .B1(n1057), .C0(n1363), 
        .Y(block_next[71]) );
  OAI221X4 U220 ( .A0(n1055), .A1(n1573), .B0(n1461), .B1(n1056), .C0(n1366), 
        .Y(block_next[68]) );
  OAI221X4 U221 ( .A0(n1055), .A1(n1613), .B0(n1445), .B1(n1056), .C0(n1358), 
        .Y(block_next[76]) );
  OAI221X4 U222 ( .A0(n1055), .A1(n1568), .B0(n1463), .B1(n1056), .C0(n1367), 
        .Y(block_next[67]) );
  OAI221X4 U223 ( .A0(n1055), .A1(n1598), .B0(n1451), .B1(n1056), .C0(n1361), 
        .Y(block_next[73]) );
  OAI221X4 U224 ( .A0(n1054), .A1(n1578), .B0(n1459), .B1(n1056), .C0(n1365), 
        .Y(block_next[69]) );
  OAI221X4 U225 ( .A0(n1055), .A1(n1563), .B0(n1465), .B1(n1056), .C0(n1368), 
        .Y(block_next[66]) );
  OAI221X4 U226 ( .A0(n1055), .A1(n1583), .B0(n1457), .B1(n1056), .C0(n1364), 
        .Y(block_next[70]) );
  NAND2X4 U227 ( .A(mem_rdata[70]), .B(n1073), .Y(n1364) );
  OAI221X4 U228 ( .A0(n1058), .A1(n1672), .B0(n1421), .B1(n1061), .C0(n1380), 
        .Y(block_next[56]) );
  OAI221X4 U229 ( .A0(n1059), .A1(n1627), .B0(n1439), .B1(n1061), .C0(n1389), 
        .Y(block_next[47]) );
  NAND2X8 U230 ( .A(valid), .B(n1299), .Y(n1303) );
  BUFX20 U231 ( .A(n1081), .Y(n1069) );
  BUFX20 U232 ( .A(n1079), .Y(n1081) );
  BUFX20 U233 ( .A(n1081), .Y(n1068) );
  INVX4 U234 ( .A(n1528), .Y(blocktag_next[3]) );
  XOR2X4 U235 ( .A(n1479), .B(proc_addr[28]), .Y(n1287) );
  CLKINVX6 U236 ( .A(tag[23]), .Y(n1479) );
  AO22X1 U237 ( .A0(proc_addr[19]), .A1(mem_read), .B0(tag[14]), .B1(mem_write), .Y(n1764) );
  OAI221X2 U238 ( .A0(n1094), .A1(n1576), .B0(n1091), .B1(n1575), .C0(n1574), 
        .Y(proc_rdata[4]) );
  BUFX20 U239 ( .A(N32), .Y(n983) );
  BUFX20 U240 ( .A(n1260), .Y(n1259) );
  INVX4 U241 ( .A(proc_reset), .Y(n1260) );
  CLKINVX8 U242 ( .A(n1778), .Y(n5) );
  INVX20 U243 ( .A(n5), .Y(mem_addr[3]) );
  CLKINVX8 U244 ( .A(n1776), .Y(n7) );
  INVX20 U245 ( .A(n7), .Y(mem_addr[5]) );
  CLKINVX8 U246 ( .A(n1775), .Y(n9) );
  INVX20 U247 ( .A(n9), .Y(mem_addr[6]) );
  CLKINVX8 U248 ( .A(n1774), .Y(n11) );
  INVX20 U249 ( .A(n11), .Y(mem_addr[7]) );
  CLKINVX8 U250 ( .A(n1772), .Y(n13) );
  INVX20 U251 ( .A(n13), .Y(mem_addr[9]) );
  CLKINVX8 U252 ( .A(n1771), .Y(n15) );
  INVX20 U253 ( .A(n15), .Y(mem_addr[10]) );
  CLKINVX8 U254 ( .A(n1770), .Y(n17) );
  INVX20 U255 ( .A(n17), .Y(mem_addr[11]) );
  CLKINVX8 U256 ( .A(n1769), .Y(n19) );
  INVX20 U257 ( .A(n19), .Y(mem_addr[12]) );
  CLKINVX8 U258 ( .A(n1768), .Y(n21) );
  INVX20 U259 ( .A(n21), .Y(mem_addr[13]) );
  CLKINVX8 U260 ( .A(n1767), .Y(n23) );
  INVX20 U261 ( .A(n23), .Y(mem_addr[14]) );
  CLKINVX8 U262 ( .A(n1766), .Y(n25) );
  INVX20 U263 ( .A(n25), .Y(mem_addr[15]) );
  CLKINVX8 U264 ( .A(n1765), .Y(n27) );
  INVX20 U265 ( .A(n27), .Y(mem_addr[16]) );
  CLKINVX8 U266 ( .A(n1764), .Y(n29) );
  INVX20 U267 ( .A(n29), .Y(mem_addr[17]) );
  CLKINVX8 U268 ( .A(n1763), .Y(n31) );
  INVX20 U269 ( .A(n31), .Y(mem_addr[18]) );
  CLKINVX6 U270 ( .A(n1762), .Y(n33) );
  INVX20 U271 ( .A(n33), .Y(mem_addr[19]) );
  AO22X1 U272 ( .A0(proc_addr[21]), .A1(mem_read), .B0(tag[16]), .B1(mem_write), .Y(n1762) );
  CLKINVX8 U273 ( .A(n1761), .Y(n35) );
  INVX20 U274 ( .A(n35), .Y(mem_addr[20]) );
  CLKINVX8 U275 ( .A(n1760), .Y(n37) );
  INVX20 U276 ( .A(n37), .Y(mem_addr[21]) );
  CLKINVX8 U277 ( .A(n1759), .Y(n39) );
  INVX20 U278 ( .A(n39), .Y(mem_addr[22]) );
  CLKINVX8 U279 ( .A(n1758), .Y(n41) );
  INVX20 U280 ( .A(n41), .Y(mem_addr[23]) );
  CLKINVX6 U281 ( .A(n1757), .Y(n43) );
  INVX20 U282 ( .A(n43), .Y(mem_addr[24]) );
  AO22X1 U283 ( .A0(proc_addr[26]), .A1(mem_read), .B0(n2), .B1(mem_write), 
        .Y(n1757) );
  CLKINVX8 U284 ( .A(n1756), .Y(n45) );
  INVX20 U285 ( .A(n45), .Y(mem_addr[25]) );
  CLKINVX8 U286 ( .A(n1755), .Y(n47) );
  INVX20 U287 ( .A(n47), .Y(mem_addr[26]) );
  CLKINVX6 U288 ( .A(n1754), .Y(n49) );
  INVX20 U289 ( .A(n49), .Y(mem_addr[27]) );
  AO22X1 U290 ( .A0(proc_addr[29]), .A1(mem_read), .B0(tag[24]), .B1(mem_write), .Y(n1754) );
  CLKINVX8 U291 ( .A(n1851), .Y(n51) );
  CLKINVX20 U292 ( .A(n51), .Y(mem_wdata[5]) );
  CLKINVX8 U293 ( .A(n1850), .Y(n53) );
  CLKINVX20 U294 ( .A(n53), .Y(mem_wdata[7]) );
  CLKINVX8 U295 ( .A(n1849), .Y(n55) );
  CLKINVX20 U296 ( .A(n55), .Y(mem_wdata[8]) );
  CLKINVX8 U297 ( .A(n1848), .Y(n57) );
  CLKINVX20 U298 ( .A(n57), .Y(mem_wdata[9]) );
  CLKINVX8 U299 ( .A(n1847), .Y(n59) );
  CLKINVX20 U300 ( .A(n59), .Y(mem_wdata[10]) );
  CLKINVX8 U301 ( .A(n1846), .Y(n61) );
  CLKINVX20 U302 ( .A(n61), .Y(mem_wdata[11]) );
  CLKINVX8 U303 ( .A(n1845), .Y(n63) );
  CLKINVX20 U304 ( .A(n63), .Y(mem_wdata[12]) );
  CLKINVX8 U305 ( .A(n1844), .Y(n65) );
  CLKINVX20 U306 ( .A(n65), .Y(mem_wdata[13]) );
  CLKINVX8 U307 ( .A(n1843), .Y(n67) );
  CLKINVX20 U308 ( .A(n67), .Y(mem_wdata[15]) );
  CLKINVX8 U309 ( .A(n1842), .Y(n69) );
  CLKINVX20 U310 ( .A(n69), .Y(mem_wdata[16]) );
  CLKINVX8 U311 ( .A(n1841), .Y(n71) );
  CLKINVX20 U312 ( .A(n71), .Y(mem_wdata[17]) );
  CLKINVX8 U313 ( .A(n1840), .Y(n73) );
  CLKINVX20 U314 ( .A(n73), .Y(mem_wdata[18]) );
  CLKINVX8 U315 ( .A(n1839), .Y(n75) );
  CLKINVX20 U316 ( .A(n75), .Y(mem_wdata[19]) );
  CLKINVX8 U317 ( .A(n1838), .Y(n77) );
  CLKINVX20 U318 ( .A(n77), .Y(mem_wdata[20]) );
  CLKINVX8 U319 ( .A(n1837), .Y(n79) );
  CLKINVX20 U320 ( .A(n79), .Y(mem_wdata[21]) );
  CLKINVX8 U321 ( .A(n1836), .Y(n81) );
  CLKINVX20 U322 ( .A(n81), .Y(mem_wdata[22]) );
  CLKINVX8 U323 ( .A(n1835), .Y(n83) );
  CLKINVX20 U324 ( .A(n83), .Y(mem_wdata[23]) );
  CLKINVX8 U325 ( .A(n1834), .Y(n85) );
  CLKINVX20 U326 ( .A(n85), .Y(mem_wdata[24]) );
  CLKINVX8 U327 ( .A(n1833), .Y(n87) );
  CLKINVX20 U328 ( .A(n87), .Y(mem_wdata[25]) );
  CLKINVX8 U329 ( .A(n1832), .Y(n89) );
  CLKINVX20 U330 ( .A(n89), .Y(mem_wdata[26]) );
  CLKINVX8 U331 ( .A(n1831), .Y(n91) );
  CLKINVX20 U332 ( .A(n91), .Y(mem_wdata[27]) );
  CLKINVX8 U333 ( .A(n1830), .Y(n93) );
  CLKINVX20 U334 ( .A(n93), .Y(mem_wdata[29]) );
  CLKINVX8 U335 ( .A(n1829), .Y(n95) );
  CLKINVX20 U336 ( .A(n95), .Y(mem_wdata[30]) );
  CLKINVX8 U337 ( .A(n1828), .Y(n97) );
  CLKINVX20 U338 ( .A(n97), .Y(mem_wdata[32]) );
  CLKINVX8 U339 ( .A(n1827), .Y(n99) );
  CLKINVX20 U340 ( .A(n99), .Y(mem_wdata[33]) );
  CLKINVX8 U341 ( .A(n1826), .Y(n101) );
  CLKINVX20 U342 ( .A(n101), .Y(mem_wdata[34]) );
  CLKINVX8 U343 ( .A(n1825), .Y(n103) );
  CLKINVX20 U344 ( .A(n103), .Y(mem_wdata[35]) );
  CLKINVX8 U345 ( .A(n1824), .Y(n105) );
  CLKINVX20 U346 ( .A(n105), .Y(mem_wdata[36]) );
  CLKINVX8 U347 ( .A(n1823), .Y(n107) );
  CLKINVX20 U348 ( .A(n107), .Y(mem_wdata[37]) );
  CLKINVX8 U349 ( .A(n1822), .Y(n109) );
  CLKINVX20 U350 ( .A(n109), .Y(mem_wdata[38]) );
  CLKINVX8 U351 ( .A(n1821), .Y(n111) );
  CLKINVX20 U352 ( .A(n111), .Y(mem_wdata[39]) );
  CLKINVX8 U353 ( .A(n1820), .Y(n113) );
  CLKINVX20 U354 ( .A(n113), .Y(mem_wdata[40]) );
  CLKINVX8 U355 ( .A(n1819), .Y(n115) );
  CLKINVX20 U356 ( .A(n115), .Y(mem_wdata[41]) );
  CLKINVX8 U357 ( .A(n1818), .Y(n117) );
  CLKINVX20 U358 ( .A(n117), .Y(mem_wdata[42]) );
  CLKINVX8 U359 ( .A(n1817), .Y(n119) );
  CLKINVX20 U360 ( .A(n119), .Y(mem_wdata[43]) );
  CLKINVX8 U361 ( .A(n1816), .Y(n121) );
  CLKINVX20 U362 ( .A(n121), .Y(mem_wdata[44]) );
  CLKINVX8 U363 ( .A(n1815), .Y(n123) );
  CLKINVX20 U364 ( .A(n123), .Y(mem_wdata[45]) );
  CLKINVX8 U365 ( .A(n1814), .Y(n125) );
  CLKINVX20 U366 ( .A(n125), .Y(mem_wdata[47]) );
  CLKINVX8 U367 ( .A(n1813), .Y(n127) );
  CLKINVX20 U368 ( .A(n127), .Y(mem_wdata[48]) );
  CLKINVX8 U369 ( .A(n1812), .Y(n129) );
  CLKINVX20 U370 ( .A(n129), .Y(mem_wdata[49]) );
  CLKINVX8 U371 ( .A(n1811), .Y(n131) );
  CLKINVX20 U372 ( .A(n131), .Y(mem_wdata[50]) );
  CLKINVX8 U373 ( .A(n1810), .Y(n133) );
  CLKINVX20 U374 ( .A(n133), .Y(mem_wdata[51]) );
  CLKINVX8 U375 ( .A(n1809), .Y(n135) );
  CLKINVX20 U376 ( .A(n135), .Y(mem_wdata[52]) );
  CLKINVX8 U377 ( .A(n1808), .Y(n137) );
  CLKINVX20 U378 ( .A(n137), .Y(mem_wdata[53]) );
  CLKINVX8 U379 ( .A(n1807), .Y(n139) );
  CLKINVX20 U380 ( .A(n139), .Y(mem_wdata[54]) );
  CLKINVX8 U381 ( .A(n1806), .Y(n141) );
  CLKINVX20 U382 ( .A(n141), .Y(mem_wdata[55]) );
  CLKINVX8 U383 ( .A(n1805), .Y(n143) );
  CLKINVX20 U384 ( .A(n143), .Y(mem_wdata[56]) );
  CLKINVX8 U385 ( .A(n1804), .Y(n145) );
  CLKINVX20 U386 ( .A(n145), .Y(mem_wdata[57]) );
  CLKINVX8 U387 ( .A(n1803), .Y(n147) );
  CLKINVX20 U388 ( .A(n147), .Y(mem_wdata[58]) );
  CLKINVX8 U389 ( .A(n1802), .Y(n149) );
  CLKINVX20 U390 ( .A(n149), .Y(mem_wdata[59]) );
  CLKINVX8 U391 ( .A(n1801), .Y(n151) );
  CLKINVX20 U392 ( .A(n151), .Y(mem_wdata[61]) );
  CLKINVX8 U393 ( .A(n1800), .Y(n153) );
  CLKINVX20 U394 ( .A(n153), .Y(mem_wdata[62]) );
  CLKINVX8 U395 ( .A(n1799), .Y(n155) );
  CLKINVX20 U396 ( .A(n155), .Y(mem_wdata[64]) );
  CLKINVX8 U397 ( .A(n1798), .Y(n157) );
  CLKINVX20 U398 ( .A(n157), .Y(mem_wdata[65]) );
  CLKINVX8 U399 ( .A(n1797), .Y(n159) );
  CLKINVX20 U400 ( .A(n159), .Y(mem_wdata[66]) );
  CLKINVX8 U401 ( .A(n1796), .Y(n161) );
  CLKINVX20 U402 ( .A(n161), .Y(mem_wdata[67]) );
  CLKINVX8 U403 ( .A(n1795), .Y(n163) );
  CLKINVX20 U404 ( .A(n163), .Y(mem_wdata[68]) );
  CLKINVX8 U405 ( .A(n1794), .Y(n165) );
  CLKINVX20 U406 ( .A(n165), .Y(mem_wdata[69]) );
  CLKINVX8 U407 ( .A(n1793), .Y(n167) );
  CLKINVX20 U408 ( .A(n167), .Y(mem_wdata[70]) );
  CLKINVX8 U409 ( .A(n1792), .Y(n169) );
  CLKINVX20 U410 ( .A(n169), .Y(mem_wdata[71]) );
  CLKINVX8 U411 ( .A(n1791), .Y(n171) );
  CLKINVX20 U412 ( .A(n171), .Y(mem_wdata[72]) );
  CLKINVX8 U413 ( .A(n1790), .Y(n173) );
  CLKINVX20 U414 ( .A(n173), .Y(mem_wdata[73]) );
  CLKINVX8 U415 ( .A(n1789), .Y(n175) );
  CLKINVX20 U416 ( .A(n175), .Y(mem_wdata[74]) );
  CLKINVX8 U417 ( .A(n1788), .Y(n177) );
  CLKINVX20 U418 ( .A(n177), .Y(mem_wdata[75]) );
  CLKINVX8 U419 ( .A(n1787), .Y(n179) );
  CLKINVX20 U420 ( .A(n179), .Y(mem_wdata[76]) );
  CLKINVX8 U421 ( .A(n1786), .Y(n181) );
  CLKINVX20 U422 ( .A(n181), .Y(mem_wdata[77]) );
  CLKINVX8 U423 ( .A(n1785), .Y(n183) );
  CLKINVX20 U424 ( .A(n183), .Y(mem_wdata[78]) );
  CLKINVX8 U425 ( .A(n1784), .Y(n185) );
  CLKINVX20 U426 ( .A(n185), .Y(mem_wdata[79]) );
  CLKINVX8 U427 ( .A(n1783), .Y(n187) );
  CLKINVX20 U428 ( .A(n187), .Y(mem_wdata[80]) );
  CLKINVX8 U429 ( .A(n1782), .Y(n189) );
  CLKINVX20 U430 ( .A(n189), .Y(mem_wdata[81]) );
  CLKINVX8 U431 ( .A(n1781), .Y(n191) );
  CLKINVX20 U432 ( .A(n191), .Y(mem_wdata[82]) );
  INVX3 U433 ( .A(n1780), .Y(n193) );
  INVX20 U434 ( .A(n193), .Y(mem_addr[1]) );
  AND2XL U435 ( .A(n1544), .B(N32), .Y(n1780) );
  CLKINVX8 U436 ( .A(n1779), .Y(n195) );
  INVX20 U437 ( .A(n195), .Y(mem_addr[2]) );
  NAND4X2 U444 ( .A(n1547), .B(n1546), .C(n1550), .D(proc_addr[0]), .Y(n1708)
         );
  CLKINVX8 U445 ( .A(proc_addr[1]), .Y(n1550) );
  XNOR2X4 U446 ( .A(tag[19]), .B(proc_addr[24]), .Y(n1289) );
  OR2X4 U447 ( .A(proc_addr[26]), .B(n2), .Y(n219) );
  XNOR2X4 U448 ( .A(tag[22]), .B(proc_addr[27]), .Y(n1279) );
  XNOR2X4 U449 ( .A(tag[24]), .B(proc_addr[29]), .Y(n1286) );
  MXI4X1 U450 ( .A(n257), .B(n258), .C(n259), .D(n260), .S0(n1047), .S1(n1012), 
        .Y(n598) );
  NAND4X6 U451 ( .A(n1264), .B(n1263), .C(n1262), .D(n1261), .Y(n1268) );
  XNOR2X2 U452 ( .A(proc_addr[23]), .B(tag[18]), .Y(n1264) );
  MXI4X1 U453 ( .A(n229), .B(n230), .C(n231), .D(n232), .S0(n1016), .S1(n1012), 
        .Y(n951) );
  MXI4X1 U454 ( .A(\blocktag[4][4] ), .B(\blocktag[5][4] ), .C(
        \blocktag[6][4] ), .D(\blocktag[7][4] ), .S0(n1047), .S1(n1013), .Y(
        n266) );
  XOR2X4 U455 ( .A(tag[0]), .B(n1535), .Y(n1288) );
  CLKINVX2 U456 ( .A(proc_addr[5]), .Y(n1535) );
  MXI4X1 U457 ( .A(\blocktag[0][4] ), .B(\blocktag[1][4] ), .C(
        \blocktag[2][4] ), .D(\blocktag[3][4] ), .S0(n1047), .S1(n1013), .Y(
        n265) );
  MXI4X2 U458 ( .A(\blocktag[0][16] ), .B(\blocktag[1][16] ), .C(
        \blocktag[2][16] ), .D(\blocktag[3][16] ), .S0(n1045), .S1(n984), .Y(
        n936) );
  BUFX20 U459 ( .A(N32), .Y(n985) );
  XOR2X4 U460 ( .A(tag[9]), .B(proc_addr[14]), .Y(n1267) );
  MX2X6 U461 ( .A(n600), .B(n601), .S0(n979), .Y(tag[9]) );
  CLKMX2X4 U462 ( .A(n618), .B(n619), .S0(n978), .Y(tag[20]) );
  MX4X1 U463 ( .A(\blocktag[4][20] ), .B(\blocktag[5][20] ), .C(
        \blocktag[6][20] ), .D(\blocktag[7][20] ), .S0(n1044), .S1(n983), .Y(
        n619) );
  MXI4XL U464 ( .A(n203), .B(n204), .C(n205), .D(n206), .S0(n1246), .S1(n983), 
        .Y(n618) );
  NOR4X8 U465 ( .A(n1268), .B(n1267), .C(n1266), .D(n1265), .Y(n1296) );
  XOR2X4 U466 ( .A(tag[7]), .B(n1521), .Y(n1274) );
  CLKINVX2 U467 ( .A(proc_addr[12]), .Y(n1521) );
  MX2X6 U468 ( .A(n598), .B(n599), .S0(n979), .Y(tag[6]) );
  MX4X1 U469 ( .A(n606), .B(n607), .C(n608), .D(n609), .S0(n1047), .S1(n1013), 
        .Y(n961) );
  INVX12 U470 ( .A(n1249), .Y(n1248) );
  MXI4X4 U471 ( .A(\blocktag[0][15] ), .B(\blocktag[1][15] ), .C(
        \blocktag[2][15] ), .D(\blocktag[3][15] ), .S0(n1045), .S1(n1011), .Y(
        n938) );
  MXI4X4 U472 ( .A(\blocktag[4][15] ), .B(\blocktag[5][15] ), .C(
        \blocktag[6][15] ), .D(\blocktag[7][15] ), .S0(n1045), .S1(n1011), .Y(
        n939) );
  MXI4X4 U473 ( .A(n245), .B(n246), .C(n247), .D(n248), .S0(n1045), .S1(n985), 
        .Y(n937) );
  MXI4X1 U474 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n1046), .S1(n1012), 
        .Y(n952) );
  CLKINVX6 U475 ( .A(n1303), .Y(n1297) );
  BUFX8 U476 ( .A(n1248), .Y(n962) );
  BUFX12 U477 ( .A(n1708), .Y(n1082) );
  INVX6 U478 ( .A(tag[1]), .Y(n1533) );
  MXI4X1 U479 ( .A(\blocktag[0][1] ), .B(\blocktag[1][1] ), .C(
        \blocktag[2][1] ), .D(\blocktag[3][1] ), .S0(n1047), .S1(n1013), .Y(
        n960) );
  MXI4X1 U480 ( .A(blockvalid[0]), .B(blockvalid[1]), .C(blockvalid[2]), .D(
        blockvalid[3]), .S0(n1043), .S1(n1011), .Y(n924) );
  BUFX20 U481 ( .A(n1019), .Y(n1043) );
  INVX8 U482 ( .A(tag[15]), .Y(n1500) );
  MX4X1 U483 ( .A(n574), .B(n575), .C(n576), .D(n577), .S0(n1047), .S1(n1013), 
        .Y(n954) );
  MX4X1 U484 ( .A(n578), .B(n579), .C(n580), .D(n581), .S0(n1047), .S1(n1013), 
        .Y(n955) );
  OA22X4 U485 ( .A0(n1088), .A1(n1613), .B0(n1084), .B1(n1612), .Y(n1614) );
  BUFX12 U486 ( .A(n1089), .Y(n1088) );
  MX4X1 U487 ( .A(n582), .B(n583), .C(n584), .D(n585), .S0(n1047), .S1(n1013), 
        .Y(n956) );
  MX4X1 U488 ( .A(n586), .B(n587), .C(n588), .D(n589), .S0(n1047), .S1(n1013), 
        .Y(n957) );
  BUFX20 U489 ( .A(n1085), .Y(n1084) );
  OA22X4 U490 ( .A0(n1089), .A1(n1698), .B0(n1085), .B1(n1697), .Y(n1699) );
  XNOR2X4 U491 ( .A(proc_addr[7]), .B(tag[2]), .Y(n1261) );
  MXI4X1 U492 ( .A(\blocktag[4][2] ), .B(\blocktag[5][2] ), .C(
        \blocktag[6][2] ), .D(\blocktag[7][2] ), .S0(n1047), .S1(n1013), .Y(
        n959) );
  MX2X6 U493 ( .A(n616), .B(n617), .S0(n978), .Y(tag[19]) );
  NOR2X6 U494 ( .A(n1292), .B(n1291), .Y(n1293) );
  NAND2X8 U495 ( .A(n1547), .B(n1546), .Y(n1551) );
  CLKINVX8 U496 ( .A(n1298), .Y(n1547) );
  NAND2X4 U497 ( .A(proc_read), .B(n1297), .Y(n1298) );
  MXI4X4 U498 ( .A(\blocktag[0][21] ), .B(\blocktag[1][21] ), .C(
        \blocktag[2][21] ), .D(\blocktag[3][21] ), .S0(n1044), .S1(n986), .Y(
        n930) );
  CLKINVX6 U499 ( .A(tag[20]), .Y(n1488) );
  MXI4X1 U500 ( .A(\blocktag[0][2] ), .B(\blocktag[1][2] ), .C(
        \blocktag[2][2] ), .D(\blocktag[3][2] ), .S0(n1047), .S1(n1013), .Y(
        n958) );
  MXI4X1 U501 ( .A(\blocktag[4][22] ), .B(\blocktag[5][22] ), .C(
        \blocktag[6][22] ), .D(\blocktag[7][22] ), .S0(n1044), .S1(n986), .Y(
        n929) );
  MX2X6 U502 ( .A(n614), .B(n615), .S0(n979), .Y(tag[0]) );
  OA22X4 U503 ( .A0(n1089), .A1(n1688), .B0(n1085), .B1(n1687), .Y(n1689) );
  MX4X4 U504 ( .A(n590), .B(n591), .C(n592), .D(n593), .S0(n1045), .S1(n983), 
        .Y(n932) );
  MX2X6 U505 ( .A(n610), .B(n611), .S0(n977), .Y(tag[24]) );
  OR2X6 U506 ( .A(n1092), .B(n1700), .Y(n225) );
  AND2XL U507 ( .A(n1253), .B(blockdata[83]), .Y(mem_wdata[83]) );
  AND2XL U508 ( .A(n1253), .B(blockdata[84]), .Y(mem_wdata[84]) );
  AND2XL U509 ( .A(n1253), .B(blockdata[85]), .Y(mem_wdata[85]) );
  AND2XL U510 ( .A(n1253), .B(blockdata[86]), .Y(mem_wdata[86]) );
  AND2XL U511 ( .A(n1253), .B(blockdata[87]), .Y(mem_wdata[87]) );
  AND2XL U512 ( .A(n1253), .B(blockdata[88]), .Y(mem_wdata[88]) );
  AND2XL U513 ( .A(n1253), .B(blockdata[89]), .Y(mem_wdata[89]) );
  AND2XL U514 ( .A(n1253), .B(blockdata[94]), .Y(mem_wdata[94]) );
  AND2XL U515 ( .A(n1253), .B(blockdata[96]), .Y(mem_wdata[96]) );
  AND2XL U516 ( .A(n1253), .B(blockdata[97]), .Y(mem_wdata[97]) );
  AND2XL U517 ( .A(n1253), .B(blockdata[98]), .Y(mem_wdata[98]) );
  AND2XL U518 ( .A(n1253), .B(blockdata[99]), .Y(mem_wdata[99]) );
  AND2XL U519 ( .A(n1253), .B(blockdata[100]), .Y(mem_wdata[100]) );
  AND2XL U520 ( .A(n1253), .B(blockdata[101]), .Y(mem_wdata[101]) );
  AND2XL U521 ( .A(n1253), .B(blockdata[102]), .Y(mem_wdata[102]) );
  AND2XL U522 ( .A(n1253), .B(blockdata[103]), .Y(mem_wdata[103]) );
  AND2XL U523 ( .A(n1253), .B(blockdata[104]), .Y(mem_wdata[104]) );
  AND2XL U524 ( .A(n1253), .B(blockdata[105]), .Y(mem_wdata[105]) );
  AND2XL U525 ( .A(N31), .B(n1544), .Y(mem_addr[0]) );
  AND2XL U526 ( .A(n1253), .B(blockdata[106]), .Y(mem_wdata[106]) );
  AND2XL U527 ( .A(n1253), .B(blockdata[107]), .Y(mem_wdata[107]) );
  AND2XL U528 ( .A(n1253), .B(blockdata[108]), .Y(mem_wdata[108]) );
  AND2XL U529 ( .A(n1253), .B(blockdata[109]), .Y(mem_wdata[109]) );
  AND2XL U530 ( .A(n1253), .B(blockdata[110]), .Y(mem_wdata[110]) );
  AND2XL U531 ( .A(n1253), .B(blockdata[112]), .Y(mem_wdata[112]) );
  AND2XL U532 ( .A(n1253), .B(blockdata[113]), .Y(mem_wdata[113]) );
  AND2XL U533 ( .A(n1253), .B(blockdata[114]), .Y(mem_wdata[114]) );
  AND2XL U534 ( .A(n1253), .B(blockdata[115]), .Y(mem_wdata[115]) );
  AND2XL U535 ( .A(n1253), .B(blockdata[116]), .Y(mem_wdata[116]) );
  AND2XL U536 ( .A(n1253), .B(blockdata[117]), .Y(mem_wdata[117]) );
  AND2XL U537 ( .A(n1253), .B(blockdata[118]), .Y(mem_wdata[118]) );
  AND2XL U538 ( .A(n1253), .B(blockdata[119]), .Y(mem_wdata[119]) );
  AND2XL U539 ( .A(n1253), .B(blockdata[120]), .Y(mem_wdata[120]) );
  AND2XL U540 ( .A(mem_write), .B(blockdata[0]), .Y(mem_wdata[0]) );
  AND2XL U541 ( .A(mem_write), .B(blockdata[121]), .Y(mem_wdata[121]) );
  MXI4X1 U542 ( .A(\blocktag[0][22] ), .B(\blocktag[1][22] ), .C(
        \blocktag[2][22] ), .D(\blocktag[3][22] ), .S0(n1044), .S1(n983), .Y(
        n928) );
  AND2XL U543 ( .A(mem_write), .B(blockdata[125]), .Y(mem_wdata[125]) );
  AND2XL U544 ( .A(mem_write), .B(blockdata[126]), .Y(mem_wdata[126]) );
  CLKINVX6 U545 ( .A(proc_addr[0]), .Y(n1549) );
  OA22X4 U546 ( .A0(n1089), .A1(n1683), .B0(n1085), .B1(n1682), .Y(n1684) );
  OAI221X2 U547 ( .A0(n1096), .A1(n1686), .B0(n1092), .B1(n1685), .C0(n1684), 
        .Y(proc_rdata[26]) );
  BUFX20 U548 ( .A(n963), .Y(n977) );
  BUFX12 U549 ( .A(N33), .Y(n963) );
  BUFX6 U550 ( .A(n1710), .Y(n1086) );
  NAND3BX4 U551 ( .AN(n1551), .B(proc_addr[1]), .C(n1549), .Y(n1710) );
  MXI4X1 U552 ( .A(n233), .B(n234), .C(n235), .D(n236), .S0(n1046), .S1(n1012), 
        .Y(n950) );
  BUFX20 U553 ( .A(n1018), .Y(n1046) );
  NAND4X4 U554 ( .A(n1288), .B(n1287), .C(n1286), .D(n1285), .Y(n1292) );
  NAND2X6 U555 ( .A(n219), .B(n220), .Y(n1285) );
  OA22X4 U556 ( .A0(n1089), .A1(n1703), .B0(n1085), .B1(n1702), .Y(n1704) );
  MX4X2 U557 ( .A(n602), .B(n604), .C(n603), .D(n605), .S0(n983), .S1(n1044), 
        .Y(n931) );
  BUFX20 U558 ( .A(n1018), .Y(n1044) );
  OAI221X2 U559 ( .A0(n1096), .A1(n1706), .B0(n1092), .B1(n1705), .C0(n1704), 
        .Y(proc_rdata[30]) );
  BUFX20 U560 ( .A(n985), .Y(n1013) );
  BUFX20 U561 ( .A(n1018), .Y(n1047) );
  OR2X4 U562 ( .A(n1096), .B(n1701), .Y(n224) );
  MX4X2 U563 ( .A(n594), .B(n595), .C(n596), .D(n597), .S0(n1045), .S1(n983), 
        .Y(n933) );
  BUFX20 U564 ( .A(n1018), .Y(n1045) );
  BUFX8 U565 ( .A(N31), .Y(n1018) );
  NAND2X4 U566 ( .A(n936), .B(n207), .Y(n208) );
  NAND2X2 U567 ( .A(n937), .B(n978), .Y(n209) );
  NAND2X6 U568 ( .A(n208), .B(n209), .Y(n210) );
  INVX1 U569 ( .A(n978), .Y(n207) );
  NAND2X2 U570 ( .A(n930), .B(n211), .Y(n212) );
  NAND2X2 U571 ( .A(n931), .B(n978), .Y(n213) );
  CLKINVX1 U572 ( .A(n978), .Y(n211) );
  NAND2X4 U573 ( .A(n1500), .B(n215), .Y(n216) );
  NAND2X8 U574 ( .A(n214), .B(proc_addr[20]), .Y(n217) );
  NAND2X8 U575 ( .A(n216), .B(n217), .Y(n1282) );
  INVX4 U576 ( .A(proc_addr[20]), .Y(n215) );
  NAND2X8 U577 ( .A(n1282), .B(n1281), .Y(n1283) );
  NAND2X6 U578 ( .A(n218), .B(proc_addr[26]), .Y(n220) );
  INVX4 U579 ( .A(n1485), .Y(n218) );
  NAND2X4 U580 ( .A(n210), .B(n221), .Y(n222) );
  NAND2X8 U581 ( .A(n222), .B(n223), .Y(n1270) );
  NAND3X4 U582 ( .A(n224), .B(n225), .C(n1699), .Y(proc_rdata[29]) );
  INVX3 U583 ( .A(blockdata[29]), .Y(n1701) );
  INVX3 U584 ( .A(blockdata[125]), .Y(n1700) );
  BUFX20 U585 ( .A(n985), .Y(n1012) );
  CLKBUFX2 U586 ( .A(N32), .Y(n986) );
  CLKBUFX2 U587 ( .A(N32), .Y(n1014) );
  BUFX8 U588 ( .A(n984), .Y(n980) );
  AND2X4 U589 ( .A(proc_addr[0]), .B(proc_addr[1]), .Y(n692) );
  BUFX20 U590 ( .A(n1250), .Y(n1254) );
  INVX4 U591 ( .A(blockdata[6]), .Y(n1586) );
  MXI2X1 U592 ( .A(n912), .B(n913), .S0(n977), .Y(blockdata[6]) );
  BUFX20 U593 ( .A(n1250), .Y(n1255) );
  BUFX3 U594 ( .A(n1753), .Y(n1250) );
  INVX4 U595 ( .A(blockdata[4]), .Y(n1576) );
  MXI2X1 U596 ( .A(n914), .B(n915), .S0(n977), .Y(blockdata[4]) );
  INVX4 U597 ( .A(blockdata[1]), .Y(n1561) );
  MXI2X2 U598 ( .A(n920), .B(n921), .S0(n977), .Y(blockdata[1]) );
  CLKAND2X12 U599 ( .A(n1256), .B(blockdata[6]), .Y(mem_wdata[6]) );
  MXI2X1 U600 ( .A(n916), .B(n917), .S0(n977), .Y(blockdata[3]) );
  CLKAND2X12 U601 ( .A(n1256), .B(blockdata[4]), .Y(mem_wdata[4]) );
  INVX4 U602 ( .A(blockdata[2]), .Y(n1566) );
  MXI2X2 U603 ( .A(n918), .B(n919), .S0(n977), .Y(blockdata[2]) );
  CLKAND2X12 U604 ( .A(n1256), .B(blockdata[3]), .Y(mem_wdata[3]) );
  NAND3BX4 U605 ( .AN(proc_addr[0]), .B(n1548), .C(n1550), .Y(n1715) );
  CLKINVX6 U606 ( .A(n1773), .Y(n226) );
  INVX20 U607 ( .A(n226), .Y(mem_addr[8]) );
  AO22X1 U608 ( .A0(proc_addr[10]), .A1(mem_read), .B0(tag[5]), .B1(mem_write), 
        .Y(n1773) );
  BUFX20 U609 ( .A(n1777), .Y(mem_addr[4]) );
  AO22XL U610 ( .A0(proc_addr[6]), .A1(mem_read), .B0(tag[1]), .B1(mem_write), 
        .Y(n1777) );
  CLKAND2X12 U611 ( .A(n1256), .B(blockdata[2]), .Y(mem_wdata[2]) );
  CLKAND2X12 U612 ( .A(n1256), .B(blockdata[1]), .Y(mem_wdata[1]) );
  BUFX3 U613 ( .A(n1251), .Y(n1256) );
  CLKAND2X12 U614 ( .A(mem_write), .B(blockdata[127]), .Y(mem_wdata[127]) );
  CLKAND2X12 U615 ( .A(mem_write), .B(blockdata[124]), .Y(mem_wdata[124]) );
  CLKAND2X12 U616 ( .A(mem_write), .B(blockdata[123]), .Y(mem_wdata[123]) );
  CLKAND2X12 U617 ( .A(mem_write), .B(blockdata[122]), .Y(mem_wdata[122]) );
  CLKAND2X12 U618 ( .A(n1254), .B(blockdata[63]), .Y(mem_wdata[63]) );
  CLKAND2X12 U619 ( .A(n1254), .B(blockdata[60]), .Y(mem_wdata[60]) );
  CLKAND2X12 U620 ( .A(n1254), .B(blockdata[46]), .Y(mem_wdata[46]) );
  CLKAND2X12 U621 ( .A(n1255), .B(blockdata[31]), .Y(mem_wdata[31]) );
  CLKAND2X12 U622 ( .A(n1255), .B(blockdata[28]), .Y(mem_wdata[28]) );
  CLKAND2X12 U623 ( .A(n1255), .B(blockdata[14]), .Y(mem_wdata[14]) );
  CLKAND2X12 U624 ( .A(n1253), .B(blockdata[111]), .Y(mem_wdata[111]) );
  CLKAND2X12 U625 ( .A(n1253), .B(blockdata[95]), .Y(mem_wdata[95]) );
  CLKAND2X12 U626 ( .A(n1253), .B(blockdata[93]), .Y(mem_wdata[93]) );
  CLKAND2X12 U627 ( .A(n1253), .B(blockdata[92]), .Y(mem_wdata[92]) );
  CLKAND2X12 U628 ( .A(n1253), .B(blockdata[91]), .Y(mem_wdata[91]) );
  CLKAND2X12 U629 ( .A(n1253), .B(blockdata[90]), .Y(mem_wdata[90]) );
  BUFX12 U630 ( .A(n988), .Y(n1007) );
  BUFX12 U631 ( .A(n990), .Y(n1002) );
  BUFX8 U632 ( .A(n989), .Y(n1005) );
  BUFX12 U633 ( .A(n1005), .Y(n1001) );
  CLKBUFX2 U634 ( .A(n989), .Y(n1006) );
  CLKBUFX2 U635 ( .A(n988), .Y(n1008) );
  CLKBUFX2 U636 ( .A(n987), .Y(n1000) );
  BUFX12 U637 ( .A(n991), .Y(n993) );
  CLKBUFX8 U638 ( .A(n1753), .Y(n1253) );
  BUFX12 U639 ( .A(n1078), .Y(n1076) );
  BUFX12 U640 ( .A(n966), .Y(n967) );
  CLKBUFX2 U641 ( .A(n991), .Y(n992) );
  BUFX12 U642 ( .A(n1092), .Y(n1091) );
  BUFX12 U643 ( .A(n1096), .Y(n1094) );
  BUFX12 U644 ( .A(n1085), .Y(n1083) );
  BUFX12 U645 ( .A(n1089), .Y(n1087) );
  OAI221X4 U646 ( .A0(n1094), .A1(n1571), .B0(n1091), .B1(n1570), .C0(n1569), 
        .Y(proc_rdata[3]) );
  OAI221X4 U647 ( .A0(n1094), .A1(n1561), .B0(n1091), .B1(n1560), .C0(n1559), 
        .Y(proc_rdata[1]) );
  CLKBUFX2 U648 ( .A(n1096), .Y(n1095) );
  AND4X6 U649 ( .A(n1337), .B(n1057), .C(n1061), .D(n1065), .Y(n569) );
  INVX2 U650 ( .A(blockdata[116]), .Y(n1655) );
  MXI4X1 U651 ( .A(n253), .B(n254), .C(n255), .D(n256), .S0(n1046), .S1(n982), 
        .Y(n944) );
  MXI4X1 U652 ( .A(n249), .B(n250), .C(n251), .D(n252), .S0(n1046), .S1(n982), 
        .Y(n945) );
  MXI4XL U653 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(n1039), .S1(n1008), 
        .Y(n676) );
  MXI4XL U654 ( .A(n295), .B(n296), .C(n297), .D(n298), .S0(n1039), .S1(n1008), 
        .Y(n677) );
  MXI4XL U655 ( .A(n369), .B(n370), .C(n371), .D(n372), .S0(n1036), .S1(n1005), 
        .Y(n759) );
  OAI221X2 U656 ( .A0(n1094), .A1(n1581), .B0(n1091), .B1(n1580), .C0(n1579), 
        .Y(proc_rdata[5]) );
  OA22X2 U657 ( .A0(n1087), .A1(n1578), .B0(n1083), .B1(n1577), .Y(n1579) );
  MXI4X2 U658 ( .A(n267), .B(n268), .C(n269), .D(n270), .S0(n1024), .S1(n1002), 
        .Y(n678) );
  MX4X1 U659 ( .A(\block[4][94] ), .B(\block[5][94] ), .C(\block[6][94] ), .D(
        \block[7][94] ), .S0(n1031), .S1(n997), .Y(n687) );
  BUFX8 U660 ( .A(n1715), .Y(n1093) );
  INVX3 U661 ( .A(blockdata[94]), .Y(n1703) );
  INVX2 U662 ( .A(blockdata[8]), .Y(n1596) );
  INVX3 U663 ( .A(blockdata[10]), .Y(n1606) );
  INVX3 U664 ( .A(blockdata[106]), .Y(n1605) );
  INVX3 U665 ( .A(blockdata[74]), .Y(n1603) );
  INVX3 U666 ( .A(blockdata[42]), .Y(n1602) );
  MXI4X1 U667 ( .A(\block[0][15] ), .B(\block[1][15] ), .C(\block[2][15] ), 
        .D(\block[3][15] ), .S0(n1041), .S1(n1009), .Y(n908) );
  MX4X1 U668 ( .A(\block[4][40] ), .B(\block[5][40] ), .C(\block[6][40] ), .D(
        \block[7][40] ), .S0(n1037), .S1(n1005), .Y(n714) );
  CLKMX2X4 U669 ( .A(n713), .B(n714), .S0(n974), .Y(blockdata[40]) );
  MX4X1 U670 ( .A(\block[4][46] ), .B(\block[5][46] ), .C(\block[6][46] ), .D(
        \block[7][46] ), .S0(n1036), .S1(n1004), .Y(n722) );
  CLKMX2X4 U671 ( .A(n721), .B(n722), .S0(n973), .Y(blockdata[46]) );
  MXI4XL U672 ( .A(n421), .B(n422), .C(n423), .D(n424), .S0(n1033), .S1(n1000), 
        .Y(n772) );
  MXI4XL U673 ( .A(n537), .B(n538), .C(n539), .D(n540), .S0(n1041), .S1(n1004), 
        .Y(n729) );
  AND2X4 U674 ( .A(n564), .B(n1259), .Y(n557) );
  AND2X6 U675 ( .A(n567), .B(n1259), .Y(n556) );
  AND2X4 U676 ( .A(n566), .B(n1259), .Y(n555) );
  AND2X4 U677 ( .A(n565), .B(n1259), .Y(n554) );
  OAI221X1 U678 ( .A0(n1094), .A1(n1596), .B0(n1091), .B1(n1595), .C0(n1594), 
        .Y(proc_rdata[8]) );
  OA22XL U679 ( .A0(n1087), .A1(n1593), .B0(n1083), .B1(n1592), .Y(n1594) );
  AND2X8 U680 ( .A(n570), .B(n1259), .Y(n563) );
  INVX4 U681 ( .A(blockdata[59]), .Y(n1687) );
  MXI2X4 U682 ( .A(n265), .B(n266), .S0(n979), .Y(tag[4]) );
  MXI4XL U683 ( .A(n237), .B(n238), .C(n239), .D(n240), .S0(n1046), .S1(n1012), 
        .Y(n953) );
  MX2X2 U684 ( .A(n682), .B(n683), .S0(n969), .Y(blockdata[93]) );
  MX2X2 U685 ( .A(n697), .B(n698), .S0(n972), .Y(blockdata[61]) );
  MXI4X2 U686 ( .A(n279), .B(n280), .C(n281), .D(n282), .S0(n1031), .S1(n997), 
        .Y(n686) );
  MX4XL U687 ( .A(\block[4][125] ), .B(\block[5][125] ), .C(\block[6][125] ), 
        .D(\block[7][125] ), .S0(n1026), .S1(n992), .Y(n689) );
  CLKMX2X4 U688 ( .A(n744), .B(n745), .S0(n971), .Y(blockdata[69]) );
  MXI4XL U689 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(n1034), .S1(n1001), 
        .Y(n760) );
  MX2X1 U690 ( .A(n699), .B(n700), .S0(n974), .Y(blockdata[34]) );
  MXI4X1 U691 ( .A(n313), .B(n314), .C(n315), .D(n316), .S0(n1042), .S1(n1010), 
        .Y(n751) );
  MX2X2 U692 ( .A(n719), .B(n720), .S0(n971), .Y(blockdata[72]) );
  MX4XL U693 ( .A(\block[4][72] ), .B(\block[5][72] ), .C(\block[6][72] ), .D(
        \block[7][72] ), .S0(n1034), .S1(n1001), .Y(n720) );
  MXI4XL U694 ( .A(n337), .B(n338), .C(n339), .D(n340), .S0(n1034), .S1(n1000), 
        .Y(n779) );
  MXI4XL U695 ( .A(n333), .B(n334), .C(n335), .D(n336), .S0(n1034), .S1(n1000), 
        .Y(n778) );
  MXI4X1 U696 ( .A(n465), .B(n466), .C(n502), .D(n504), .S0(n1028), .S1(n995), 
        .Y(n736) );
  MXI4XL U697 ( .A(n549), .B(n550), .C(n551), .D(n552), .S0(n1036), .S1(n1004), 
        .Y(n775) );
  MXI4XL U698 ( .A(n545), .B(n546), .C(n547), .D(n548), .S0(n1036), .S1(n1004), 
        .Y(n774) );
  BUFX16 U699 ( .A(n984), .Y(n1011) );
  BUFX12 U700 ( .A(n987), .Y(n997) );
  BUFX12 U701 ( .A(n981), .Y(n998) );
  CLKBUFX2 U702 ( .A(n1014), .Y(n996) );
  CLKBUFX2 U703 ( .A(n1014), .Y(n1010) );
  BUFX8 U704 ( .A(n1005), .Y(n1004) );
  CLKBUFX2 U705 ( .A(n987), .Y(n994) );
  CLKBUFX2 U706 ( .A(n987), .Y(n1009) );
  CLKBUFX2 U707 ( .A(n981), .Y(n999) );
  CLKBUFX2 U708 ( .A(n987), .Y(n1003) );
  CLKBUFX4 U709 ( .A(n1170), .Y(n1183) );
  CLKBUFX4 U710 ( .A(n1132), .Y(n1145) );
  CLKBUFX4 U711 ( .A(n1208), .Y(n1221) );
  CLKBUFX4 U712 ( .A(n1189), .Y(n1202) );
  CLKBUFX4 U713 ( .A(n1151), .Y(n1164) );
  CLKBUFX4 U714 ( .A(n1227), .Y(n1240) );
  BUFX4 U715 ( .A(n1172), .Y(n1188) );
  BUFX4 U716 ( .A(n1134), .Y(n1150) );
  CLKBUFX2 U717 ( .A(n1172), .Y(n1187) );
  CLKBUFX2 U718 ( .A(n1134), .Y(n1149) );
  BUFX4 U719 ( .A(n1210), .Y(n1226) );
  CLKBUFX2 U720 ( .A(n1210), .Y(n1225) );
  BUFX4 U721 ( .A(n1099), .Y(n1112) );
  BUFX20 U722 ( .A(n962), .Y(n979) );
  BUFX8 U723 ( .A(n1017), .Y(n1019) );
  BUFX8 U724 ( .A(n1016), .Y(n1021) );
  BUFX8 U725 ( .A(n1015), .Y(n1025) );
  BUFX8 U726 ( .A(n1248), .Y(n964) );
  BUFX8 U727 ( .A(n1045), .Y(n1022) );
  CLKBUFX2 U728 ( .A(n1248), .Y(n965) );
  BUFX4 U729 ( .A(n1191), .Y(n1207) );
  BUFX4 U730 ( .A(n1153), .Y(n1169) );
  CLKBUFX2 U731 ( .A(n1191), .Y(n1206) );
  CLKBUFX2 U732 ( .A(n1153), .Y(n1168) );
  BUFX4 U733 ( .A(n1229), .Y(n1245) );
  CLKBUFX2 U734 ( .A(n1229), .Y(n1244) );
  INVX3 U735 ( .A(n1472), .Y(proc_stall) );
  BUFX8 U736 ( .A(n1713), .Y(n1090) );
  OAI221X4 U737 ( .A0(n1096), .A1(n1691), .B0(n1092), .B1(n1690), .C0(n1689), 
        .Y(proc_rdata[27]) );
  OA22XL U738 ( .A0(n1087), .A1(n1573), .B0(n1083), .B1(n1572), .Y(n1574) );
  OA22XL U739 ( .A0(n1087), .A1(n1558), .B0(n1083), .B1(n1557), .Y(n1559) );
  OA22XL U740 ( .A0(n1087), .A1(n1568), .B0(n1083), .B1(n1567), .Y(n1569) );
  OA22XL U741 ( .A0(n1087), .A1(n1563), .B0(n1083), .B1(n1562), .Y(n1564) );
  OA22XL U742 ( .A0(n1087), .A1(n1588), .B0(n1083), .B1(n1587), .Y(n1589) );
  OA22XL U743 ( .A0(n1088), .A1(n1643), .B0(n1084), .B1(n1642), .Y(n1644) );
  OA22XL U744 ( .A0(n1088), .A1(n1653), .B0(n1084), .B1(n1652), .Y(n1654) );
  OA22XL U745 ( .A0(n1088), .A1(n1663), .B0(n1084), .B1(n1662), .Y(n1664) );
  OA22XL U746 ( .A0(n1088), .A1(n1638), .B0(n1084), .B1(n1637), .Y(n1639) );
  OA22XL U747 ( .A0(n1088), .A1(n1648), .B0(n1084), .B1(n1647), .Y(n1649) );
  OA22XL U748 ( .A0(n1088), .A1(n1658), .B0(n1084), .B1(n1657), .Y(n1659) );
  OA22XL U749 ( .A0(n1088), .A1(n1668), .B0(n1084), .B1(n1667), .Y(n1669) );
  OA22XL U750 ( .A0(n1088), .A1(n1633), .B0(n1084), .B1(n1632), .Y(n1634) );
  INVX3 U751 ( .A(n1543), .Y(n1753) );
  NOR2XL U752 ( .A(n1248), .B(N32), .Y(n1748) );
  AND2XL U753 ( .A(n1749), .B(N31), .Y(n566) );
  AND2XL U754 ( .A(n1750), .B(N31), .Y(n567) );
  AND2XL U755 ( .A(n1748), .B(N31), .Y(n564) );
  AND2XL U756 ( .A(n1751), .B(N31), .Y(n565) );
  AND2X8 U757 ( .A(n572), .B(n1259), .Y(n561) );
  AND2X8 U758 ( .A(n573), .B(n1259), .Y(n562) );
  AND2X4 U759 ( .A(n571), .B(n1259), .Y(n560) );
  INVX6 U760 ( .A(blockdata[27]), .Y(n1691) );
  INVX3 U761 ( .A(blockdata[30]), .Y(n1706) );
  INVX4 U762 ( .A(blockdata[26]), .Y(n1686) );
  INVX3 U763 ( .A(blockdata[126]), .Y(n1705) );
  INVX4 U764 ( .A(blockdata[122]), .Y(n1685) );
  INVX4 U765 ( .A(blockdata[91]), .Y(n1688) );
  INVX4 U766 ( .A(blockdata[90]), .Y(n1683) );
  INVX3 U767 ( .A(blockdata[62]), .Y(n1702) );
  INVX4 U768 ( .A(blockdata[58]), .Y(n1682) );
  NAND2X1 U769 ( .A(n1543), .B(n1545), .Y(n1544) );
  INVX2 U770 ( .A(blockdata[104]), .Y(n1595) );
  INVX2 U771 ( .A(blockdata[32]), .Y(n1552) );
  INVX2 U772 ( .A(blockdata[98]), .Y(n1565) );
  INVX2 U773 ( .A(blockdata[0]), .Y(n1556) );
  INVX2 U774 ( .A(blockdata[97]), .Y(n1560) );
  INVX2 U775 ( .A(blockdata[96]), .Y(n1555) );
  INVX2 U776 ( .A(blockdata[102]), .Y(n1585) );
  INVX2 U777 ( .A(blockdata[66]), .Y(n1563) );
  INVX2 U778 ( .A(blockdata[67]), .Y(n1568) );
  INVX2 U779 ( .A(blockdata[65]), .Y(n1558) );
  INVX2 U780 ( .A(blockdata[68]), .Y(n1573) );
  INVX2 U781 ( .A(blockdata[64]), .Y(n1553) );
  INVX3 U782 ( .A(blockdata[103]), .Y(n1590) );
  INVX3 U783 ( .A(blockdata[7]), .Y(n1591) );
  INVX3 U784 ( .A(blockdata[5]), .Y(n1581) );
  INVX3 U785 ( .A(blockdata[99]), .Y(n1570) );
  INVX3 U786 ( .A(blockdata[100]), .Y(n1575) );
  INVX3 U787 ( .A(blockdata[101]), .Y(n1580) );
  INVX3 U788 ( .A(blockdata[9]), .Y(n1601) );
  INVX3 U789 ( .A(blockdata[11]), .Y(n1611) );
  INVX3 U790 ( .A(blockdata[12]), .Y(n1616) );
  INVX3 U791 ( .A(blockdata[13]), .Y(n1621) );
  INVX3 U792 ( .A(blockdata[107]), .Y(n1610) );
  INVX3 U793 ( .A(blockdata[105]), .Y(n1600) );
  INVX3 U794 ( .A(blockdata[110]), .Y(n1625) );
  INVX3 U795 ( .A(blockdata[108]), .Y(n1615) );
  INVX3 U796 ( .A(blockdata[109]), .Y(n1620) );
  INVX3 U797 ( .A(blockdata[73]), .Y(n1598) );
  INVX3 U798 ( .A(blockdata[75]), .Y(n1608) );
  INVX3 U799 ( .A(blockdata[78]), .Y(n1623) );
  INVX3 U800 ( .A(blockdata[76]), .Y(n1613) );
  INVX3 U801 ( .A(blockdata[77]), .Y(n1618) );
  INVX3 U802 ( .A(blockdata[79]), .Y(n1628) );
  INVX3 U803 ( .A(blockdata[41]), .Y(n1597) );
  INVX3 U804 ( .A(blockdata[43]), .Y(n1607) );
  INVX3 U805 ( .A(blockdata[44]), .Y(n1612) );
  INVX3 U806 ( .A(blockdata[47]), .Y(n1627) );
  INVX3 U807 ( .A(blockdata[45]), .Y(n1617) );
  INVX4 U808 ( .A(blockdata[36]), .Y(n1572) );
  INVX2 U809 ( .A(blockdata[25]), .Y(n1681) );
  INVX2 U810 ( .A(blockdata[22]), .Y(n1666) );
  INVX2 U811 ( .A(blockdata[21]), .Y(n1661) );
  INVX2 U812 ( .A(blockdata[23]), .Y(n1671) );
  INVX2 U813 ( .A(blockdata[24]), .Y(n1676) );
  INVX2 U814 ( .A(blockdata[117]), .Y(n1660) );
  INVX2 U815 ( .A(blockdata[121]), .Y(n1680) );
  INVX2 U816 ( .A(blockdata[119]), .Y(n1670) );
  INVX2 U817 ( .A(blockdata[120]), .Y(n1675) );
  INVX2 U818 ( .A(blockdata[118]), .Y(n1665) );
  INVX2 U819 ( .A(blockdata[57]), .Y(n1677) );
  INVX2 U820 ( .A(blockdata[87]), .Y(n1668) );
  INVX2 U821 ( .A(blockdata[89]), .Y(n1678) );
  INVX2 U822 ( .A(blockdata[88]), .Y(n1673) );
  INVX2 U823 ( .A(blockdata[82]), .Y(n1643) );
  INVX2 U824 ( .A(blockdata[81]), .Y(n1638) );
  INVX2 U825 ( .A(blockdata[83]), .Y(n1648) );
  INVX2 U826 ( .A(blockdata[84]), .Y(n1653) );
  INVX2 U827 ( .A(blockdata[86]), .Y(n1663) );
  INVX2 U828 ( .A(blockdata[85]), .Y(n1658) );
  NAND3BXL U829 ( .AN(n1550), .B(n1302), .C(n1549), .Y(n1372) );
  NAND2XL U830 ( .A(n1302), .B(n692), .Y(n1336) );
  MXI2X4 U831 ( .A(n958), .B(n959), .S0(n979), .Y(tag[2]) );
  MX4XL U832 ( .A(n1735), .B(n1734), .C(n1733), .D(n1732), .S0(n1043), .S1(
        n1011), .Y(n925) );
  MXI4XL U833 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n1046), .S1(n1012), 
        .Y(n599) );
  MX4XL U834 ( .A(\blocktag[0][9] ), .B(\blocktag[1][9] ), .C(\blocktag[2][9] ), .D(\blocktag[3][9] ), .S0(n1046), .S1(n1012), .Y(n600) );
  MX4XL U835 ( .A(\blocktag[4][9] ), .B(\blocktag[5][9] ), .C(\blocktag[6][9] ), .D(\blocktag[7][9] ), .S0(n1046), .S1(n1012), .Y(n601) );
  MX4XL U836 ( .A(\blocktag[0][0] ), .B(\blocktag[1][0] ), .C(\blocktag[2][0] ), .D(\blocktag[3][0] ), .S0(n1047), .S1(n1013), .Y(n614) );
  MX4XL U837 ( .A(\blocktag[4][0] ), .B(\blocktag[5][0] ), .C(\blocktag[6][0] ), .D(\blocktag[7][0] ), .S0(n1047), .S1(n1013), .Y(n615) );
  CLKINVX8 U838 ( .A(N33), .Y(n1249) );
  XOR2X4 U839 ( .A(tag[6]), .B(proc_addr[11]), .Y(n1265) );
  XOR2X4 U840 ( .A(tag[4]), .B(proc_addr[9]), .Y(n1266) );
  CLKMX2X4 U841 ( .A(n680), .B(n681), .S0(n975), .Y(blockdata[29]) );
  CLKMX2X4 U842 ( .A(n688), .B(n689), .S0(n967), .Y(blockdata[125]) );
  MXI4X1 U843 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(n1026), .S1(n992), 
        .Y(n690) );
  MXI4X1 U844 ( .A(n275), .B(n276), .C(n277), .D(n278), .S0(n1026), .S1(n992), 
        .Y(n691) );
  MX4XL U845 ( .A(\block[0][59] ), .B(\block[1][59] ), .C(\block[2][59] ), .D(
        \block[3][59] ), .S0(n1022), .S1(n1002), .Y(n695) );
  MX4XL U846 ( .A(\block[4][59] ), .B(\block[5][59] ), .C(\block[6][59] ), .D(
        \block[7][59] ), .S0(n1022), .S1(n1002), .Y(n696) );
  MX4XL U847 ( .A(\block[0][27] ), .B(\block[1][27] ), .C(\block[2][27] ), .D(
        \block[3][27] ), .S0(n1039), .S1(n1007), .Y(n670) );
  MX4XL U848 ( .A(\block[4][27] ), .B(\block[5][27] ), .C(\block[6][27] ), .D(
        \block[7][27] ), .S0(n1039), .S1(n1007), .Y(n671) );
  MXI4XL U849 ( .A(n283), .B(n284), .C(n285), .D(n286), .S0(n1022), .S1(n1002), 
        .Y(n672) );
  MXI4XL U850 ( .A(n287), .B(n288), .C(n289), .D(n290), .S0(n1022), .S1(n1002), 
        .Y(n673) );
  MXI2X2 U851 ( .A(n299), .B(n300), .S0(n967), .Y(blockdata[123]) );
  MXI4XL U852 ( .A(\block[0][123] ), .B(\block[1][123] ), .C(\block[2][123] ), 
        .D(\block[3][123] ), .S0(n1026), .S1(n992), .Y(n299) );
  MXI4XL U853 ( .A(\block[4][123] ), .B(\block[5][123] ), .C(\block[6][123] ), 
        .D(\block[7][123] ), .S0(n1026), .S1(n992), .Y(n300) );
  MX4XL U854 ( .A(\block[0][122] ), .B(\block[1][122] ), .C(\block[2][122] ), 
        .D(\block[3][122] ), .S0(n1027), .S1(n993), .Y(n693) );
  MX4XL U855 ( .A(\block[0][91] ), .B(\block[1][91] ), .C(\block[2][91] ), .D(
        \block[3][91] ), .S0(n1031), .S1(n998), .Y(n668) );
  MX4XL U856 ( .A(\block[4][91] ), .B(\block[5][91] ), .C(\block[6][91] ), .D(
        \block[7][91] ), .S0(n1031), .S1(n998), .Y(n669) );
  MXI4XL U857 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(n1031), .S1(n998), 
        .Y(n674) );
  MXI4XL U858 ( .A(n305), .B(n306), .C(n307), .D(n308), .S0(n1031), .S1(n998), 
        .Y(n675) );
  MXI2XL U859 ( .A(tag[3]), .B(proc_addr[8]), .S0(n1068), .Y(n1528) );
  MXI2XL U860 ( .A(tag[4]), .B(proc_addr[9]), .S0(n1068), .Y(n1527) );
  MXI2XL U861 ( .A(tag[6]), .B(proc_addr[11]), .S0(n1068), .Y(n1523) );
  MXI2XL U862 ( .A(tag[9]), .B(proc_addr[14]), .S0(n1068), .Y(n1517) );
  MX4XL U863 ( .A(n620), .B(n621), .C(n622), .D(n623), .S0(n1022), .S1(n1014), 
        .Y(n859) );
  MXI4XL U864 ( .A(\block[0][63] ), .B(\block[1][63] ), .C(\block[2][63] ), 
        .D(\block[3][63] ), .S0(n1022), .S1(n990), .Y(n858) );
  MX4XL U865 ( .A(n632), .B(n633), .C(n634), .D(n635), .S0(n1039), .S1(n1007), 
        .Y(n884) );
  MXI4XL U866 ( .A(\block[4][31] ), .B(\block[5][31] ), .C(\block[6][31] ), 
        .D(\block[7][31] ), .S0(n1038), .S1(n1007), .Y(n885) );
  MX4XL U867 ( .A(n640), .B(n641), .C(n642), .D(n643), .S0(n1022), .S1(n1002), 
        .Y(n861) );
  MX4XL U868 ( .A(n636), .B(n637), .C(n638), .D(n639), .S0(n1022), .S1(n1002), 
        .Y(n860) );
  MX4XL U869 ( .A(n664), .B(n665), .C(n666), .D(n667), .S0(n1039), .S1(n1007), 
        .Y(n887) );
  MX4XL U870 ( .A(n660), .B(n661), .C(n662), .D(n663), .S0(n1039), .S1(n1007), 
        .Y(n886) );
  MX4XL U871 ( .A(n628), .B(n629), .C(n630), .D(n631), .S0(n1026), .S1(n992), 
        .Y(n791) );
  MXI4XL U872 ( .A(\block[0][127] ), .B(\block[1][127] ), .C(\block[2][127] ), 
        .D(\block[3][127] ), .S0(n1026), .S1(n992), .Y(n790) );
  MX4XL U873 ( .A(n656), .B(n657), .C(n658), .D(n659), .S0(n1026), .S1(n992), 
        .Y(n793) );
  MX4XL U874 ( .A(n652), .B(n653), .C(n654), .D(n655), .S0(n1026), .S1(n992), 
        .Y(n792) );
  MX4XL U875 ( .A(n648), .B(n649), .C(n650), .D(n651), .S0(n1031), .S1(n998), 
        .Y(n827) );
  MX4XL U876 ( .A(n644), .B(n645), .C(n646), .D(n647), .S0(n1031), .S1(n998), 
        .Y(n826) );
  MX4XL U877 ( .A(n624), .B(n625), .C(n626), .D(n627), .S0(n1031), .S1(n997), 
        .Y(n825) );
  MXI4XL U878 ( .A(\block[0][95] ), .B(\block[1][95] ), .C(\block[2][95] ), 
        .D(\block[3][95] ), .S0(n1031), .S1(n997), .Y(n824) );
  NAND2XL U879 ( .A(mem_rdata[8]), .B(n1070), .Y(n1452) );
  NAND2XL U880 ( .A(mem_rdata[14]), .B(n1071), .Y(n1440) );
  NAND2XL U881 ( .A(mem_rdata[27]), .B(n1070), .Y(n1414) );
  NAND2XL U882 ( .A(mem_rdata[0]), .B(n1069), .Y(n1468) );
  MXI2X2 U883 ( .A(n908), .B(n909), .S0(n976), .Y(blockdata[15]) );
  MXI4XL U884 ( .A(n309), .B(n310), .C(n311), .D(n312), .S0(n1043), .S1(n1010), 
        .Y(n750) );
  MX2XL U885 ( .A(n701), .B(n702), .S0(n974), .Y(blockdata[35]) );
  MXI4XL U886 ( .A(n317), .B(n318), .C(n319), .D(n320), .S0(n1038), .S1(n1006), 
        .Y(n705) );
  MXI4XL U887 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n1038), .S1(n1006), 
        .Y(n706) );
  CLKMX2X2 U888 ( .A(n707), .B(n708), .S0(n974), .Y(blockdata[37]) );
  NAND2XL U889 ( .A(mem_rdata[105]), .B(n1076), .Y(n1326) );
  NAND2XL U890 ( .A(mem_rdata[79]), .B(n1074), .Y(n1355) );
  NAND2XL U891 ( .A(mem_rdata[92]), .B(n1075), .Y(n1342) );
  NAND2XL U892 ( .A(mem_rdata[53]), .B(n1077), .Y(n1383) );
  NAND2XL U893 ( .A(mem_rdata[118]), .B(n1077), .Y(n1313) );
  MX4XL U894 ( .A(\block[0][69] ), .B(\block[1][69] ), .C(\block[2][69] ), .D(
        \block[3][69] ), .S0(n1040), .S1(n1001), .Y(n744) );
  MX4XL U895 ( .A(\block[4][69] ), .B(\block[5][69] ), .C(\block[6][69] ), .D(
        \block[7][69] ), .S0(n1028), .S1(n1001), .Y(n745) );
  MXI4XL U896 ( .A(n325), .B(n326), .C(n327), .D(n328), .S0(n1034), .S1(n1001), 
        .Y(n723) );
  MXI4XL U897 ( .A(n329), .B(n330), .C(n331), .D(n332), .S0(n1034), .S1(n1001), 
        .Y(n724) );
  MXI4XL U898 ( .A(n345), .B(n346), .C(n347), .D(n348), .S0(n1034), .S1(n1001), 
        .Y(n761) );
  MXI4XL U899 ( .A(n349), .B(n350), .C(n351), .D(n352), .S0(n1037), .S1(n1005), 
        .Y(n766) );
  MXI4XL U900 ( .A(n353), .B(n354), .C(n355), .D(n356), .S0(n1037), .S1(n1005), 
        .Y(n767) );
  MXI4XL U901 ( .A(n357), .B(n358), .C(n359), .D(n360), .S0(n1037), .S1(n1005), 
        .Y(n715) );
  MXI4XL U902 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(n1037), .S1(n1005), 
        .Y(n716) );
  MXI4XL U903 ( .A(n365), .B(n366), .C(n367), .D(n368), .S0(n1037), .S1(n1005), 
        .Y(n758) );
  MXI4XL U904 ( .A(n373), .B(n374), .C(n375), .D(n376), .S0(n1029), .S1(n995), 
        .Y(n776) );
  MXI4XL U905 ( .A(n377), .B(n378), .C(n379), .D(n380), .S0(n1029), .S1(n995), 
        .Y(n777) );
  MXI4XL U906 ( .A(n381), .B(n382), .C(n383), .D(n384), .S0(n1029), .S1(n995), 
        .Y(n786) );
  MXI4XL U907 ( .A(n385), .B(n386), .C(n387), .D(n388), .S0(n1029), .S1(n995), 
        .Y(n787) );
  MXI4XL U908 ( .A(n389), .B(n390), .C(n391), .D(n392), .S0(n1029), .S1(n995), 
        .Y(n725) );
  MXI4XL U909 ( .A(n393), .B(n394), .C(n395), .D(n396), .S0(n1029), .S1(n995), 
        .Y(n726) );
  MXI4XL U910 ( .A(n397), .B(n398), .C(n399), .D(n400), .S0(n1029), .S1(n995), 
        .Y(n733) );
  MXI4XL U911 ( .A(n401), .B(n402), .C(n403), .D(n404), .S0(n1029), .S1(n995), 
        .Y(n734) );
  MXI4X1 U912 ( .A(n405), .B(n406), .C(n407), .D(n408), .S0(n1036), .S1(n1004), 
        .Y(n762) );
  MXI4X1 U913 ( .A(n409), .B(n410), .C(n411), .D(n412), .S0(n1036), .S1(n1004), 
        .Y(n763) );
  MXI4XL U914 ( .A(n413), .B(n414), .C(n415), .D(n416), .S0(n1033), .S1(n1000), 
        .Y(n731) );
  MXI4XL U915 ( .A(n417), .B(n418), .C(n419), .D(n420), .S0(n1033), .S1(n1000), 
        .Y(n732) );
  MXI4XL U916 ( .A(n425), .B(n426), .C(n427), .D(n428), .S0(n1033), .S1(n1000), 
        .Y(n773) );
  CLKMX2X4 U917 ( .A(n780), .B(n781), .S0(n976), .Y(blockdata[14]) );
  MX4XL U918 ( .A(\block[0][14] ), .B(\block[1][14] ), .C(\block[2][14] ), .D(
        \block[3][14] ), .S0(n1041), .S1(n1004), .Y(n780) );
  MX4XL U919 ( .A(\block[4][14] ), .B(\block[5][14] ), .C(\block[6][14] ), .D(
        \block[7][14] ), .S0(n1041), .S1(n1004), .Y(n781) );
  MXI4XL U920 ( .A(n429), .B(n430), .C(n431), .D(n432), .S0(n1028), .S1(n995), 
        .Y(n784) );
  MXI4XL U921 ( .A(n433), .B(n434), .C(n435), .D(n436), .S0(n1028), .S1(n995), 
        .Y(n785) );
  MX2XL U922 ( .A(n711), .B(n712), .S0(n971), .Y(blockdata[70]) );
  MX4XL U923 ( .A(\block[0][70] ), .B(\block[1][70] ), .C(\block[2][70] ), .D(
        \block[3][70] ), .S0(n1022), .S1(n1001), .Y(n711) );
  MX4XL U924 ( .A(\block[4][70] ), .B(\block[5][70] ), .C(\block[6][70] ), .D(
        \block[7][70] ), .S0(n1034), .S1(n1001), .Y(n712) );
  MX4XL U925 ( .A(\block[0][99] ), .B(\block[1][99] ), .C(\block[2][99] ), .D(
        \block[3][99] ), .S0(n1030), .S1(n996), .Y(n703) );
  MX4XL U926 ( .A(\block[4][99] ), .B(\block[5][99] ), .C(\block[6][99] ), .D(
        \block[7][99] ), .S0(n1030), .S1(n996), .Y(n704) );
  MX4XL U927 ( .A(\block[0][100] ), .B(\block[1][100] ), .C(\block[2][100] ), 
        .D(\block[3][100] ), .S0(n1030), .S1(n996), .Y(n742) );
  MX4XL U928 ( .A(\block[4][100] ), .B(\block[5][100] ), .C(\block[6][100] ), 
        .D(\block[7][100] ), .S0(n1030), .S1(n996), .Y(n743) );
  MX2XL U929 ( .A(n709), .B(n710), .S0(n974), .Y(blockdata[38]) );
  MX4XL U930 ( .A(\block[0][38] ), .B(\block[1][38] ), .C(\block[2][38] ), .D(
        \block[3][38] ), .S0(n1037), .S1(n1006), .Y(n709) );
  MX4XL U931 ( .A(\block[4][38] ), .B(\block[5][38] ), .C(\block[6][38] ), .D(
        \block[7][38] ), .S0(n1037), .S1(n1006), .Y(n710) );
  MXI4XL U932 ( .A(n437), .B(n438), .C(n439), .D(n440), .S0(n1037), .S1(n1005), 
        .Y(n717) );
  MXI4XL U933 ( .A(n441), .B(n442), .C(n443), .D(n444), .S0(n1037), .S1(n1005), 
        .Y(n718) );
  MXI4XL U934 ( .A(n445), .B(n446), .C(n447), .D(n448), .S0(n1034), .S1(n1000), 
        .Y(n768) );
  MXI4XL U935 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n1034), .S1(n1000), 
        .Y(n769) );
  MXI4XL U936 ( .A(n453), .B(n454), .C(n455), .D(n456), .S0(n1033), .S1(n1000), 
        .Y(n782) );
  MXI4XL U937 ( .A(n457), .B(n458), .C(n459), .D(n460), .S0(n1033), .S1(n1000), 
        .Y(n783) );
  MXI4XL U938 ( .A(n461), .B(n462), .C(n463), .D(n464), .S0(n1029), .S1(n995), 
        .Y(n735) );
  CLKMX2X4 U939 ( .A(n788), .B(n789), .S0(n968), .Y(blockdata[111]) );
  MXI4XL U940 ( .A(n505), .B(n506), .C(n507), .D(n508), .S0(n1042), .S1(n1004), 
        .Y(n770) );
  MXI4XL U941 ( .A(n509), .B(n510), .C(n511), .D(n512), .S0(n1042), .S1(n1004), 
        .Y(n771) );
  MXI4XL U942 ( .A(n513), .B(n514), .C(n515), .D(n516), .S0(n1042), .S1(n1004), 
        .Y(n737) );
  MXI4XL U943 ( .A(n517), .B(n518), .C(n519), .D(n520), .S0(n1042), .S1(n1004), 
        .Y(n738) );
  MXI4XL U944 ( .A(n521), .B(n522), .C(n523), .D(n524), .S0(n1042), .S1(n1004), 
        .Y(n764) );
  MXI4XL U945 ( .A(n525), .B(n526), .C(n527), .D(n528), .S0(n1042), .S1(n1004), 
        .Y(n765) );
  MXI4XL U946 ( .A(n529), .B(n530), .C(n531), .D(n532), .S0(n1041), .S1(n1004), 
        .Y(n727) );
  MXI4XL U947 ( .A(n533), .B(n534), .C(n535), .D(n536), .S0(n1041), .S1(n1004), 
        .Y(n728) );
  MXI4XL U948 ( .A(n541), .B(n542), .C(n543), .D(n544), .S0(n1041), .S1(n1004), 
        .Y(n730) );
  MX2X1 U949 ( .A(n740), .B(n741), .S0(n974), .Y(blockdata[33]) );
  MX2XL U950 ( .A(n748), .B(n749), .S0(n974), .Y(blockdata[39]) );
  MX4XL U951 ( .A(\block[0][39] ), .B(\block[1][39] ), .C(\block[2][39] ), .D(
        \block[3][39] ), .S0(n1037), .S1(n1005), .Y(n748) );
  MX4XL U952 ( .A(\block[4][39] ), .B(\block[5][39] ), .C(\block[6][39] ), .D(
        \block[7][39] ), .S0(n1037), .S1(n1005), .Y(n749) );
  MX2XL U953 ( .A(n752), .B(n753), .S0(n971), .Y(blockdata[71]) );
  MX4XL U954 ( .A(\block[0][71] ), .B(\block[1][71] ), .C(\block[2][71] ), .D(
        \block[3][71] ), .S0(n1034), .S1(n1001), .Y(n752) );
  MX4XL U955 ( .A(\block[4][71] ), .B(\block[5][71] ), .C(\block[6][71] ), .D(
        \block[7][71] ), .S0(n1034), .S1(n1001), .Y(n753) );
  MXI2XL U956 ( .A(n846), .B(n847), .S0(n971), .Y(blockdata[80]) );
  MXI4XL U957 ( .A(\block[4][80] ), .B(\block[5][80] ), .C(\block[6][80] ), 
        .D(\block[7][80] ), .S0(n1033), .S1(n1000), .Y(n847) );
  MXI4XL U958 ( .A(\block[0][80] ), .B(\block[1][80] ), .C(\block[2][80] ), 
        .D(\block[3][80] ), .S0(n1033), .S1(n1000), .Y(n846) );
  MXI2XL U959 ( .A(n808), .B(n809), .S0(n968), .Y(blockdata[114]) );
  MXI4XL U960 ( .A(\block[4][114] ), .B(\block[5][114] ), .C(\block[6][114] ), 
        .D(\block[7][114] ), .S0(n1028), .S1(n994), .Y(n809) );
  MXI4XL U961 ( .A(\block[0][114] ), .B(\block[1][114] ), .C(\block[2][114] ), 
        .D(\block[3][114] ), .S0(n1028), .S1(n994), .Y(n808) );
  MXI2XL U962 ( .A(n810), .B(n811), .S0(n968), .Y(blockdata[113]) );
  MXI4XL U963 ( .A(\block[4][113] ), .B(\block[5][113] ), .C(\block[6][113] ), 
        .D(\block[7][113] ), .S0(n1028), .S1(n994), .Y(n811) );
  MXI4XL U964 ( .A(\block[0][113] ), .B(\block[1][113] ), .C(\block[2][113] ), 
        .D(\block[3][113] ), .S0(n1028), .S1(n994), .Y(n810) );
  MXI2XL U965 ( .A(n806), .B(n807), .S0(n968), .Y(blockdata[115]) );
  MXI4XL U966 ( .A(\block[4][115] ), .B(\block[5][115] ), .C(\block[6][115] ), 
        .D(\block[7][115] ), .S0(n1028), .S1(n994), .Y(n807) );
  MXI4XL U967 ( .A(\block[0][115] ), .B(\block[1][115] ), .C(\block[2][115] ), 
        .D(\block[3][115] ), .S0(n1028), .S1(n994), .Y(n806) );
  MXI2XL U968 ( .A(n812), .B(n813), .S0(n968), .Y(blockdata[112]) );
  MXI4XL U969 ( .A(\block[4][112] ), .B(\block[5][112] ), .C(\block[6][112] ), 
        .D(\block[7][112] ), .S0(n1028), .S1(n994), .Y(n813) );
  MXI4XL U970 ( .A(\block[0][112] ), .B(\block[1][112] ), .C(\block[2][112] ), 
        .D(\block[3][112] ), .S0(n1028), .S1(n994), .Y(n812) );
  MXI2XL U971 ( .A(n904), .B(n905), .S0(n976), .Y(blockdata[17]) );
  MXI4XL U972 ( .A(\block[4][17] ), .B(\block[5][17] ), .C(\block[6][17] ), 
        .D(\block[7][17] ), .S0(n1041), .S1(n1009), .Y(n905) );
  MXI4XL U973 ( .A(\block[0][17] ), .B(\block[1][17] ), .C(\block[2][17] ), 
        .D(\block[3][17] ), .S0(n1041), .S1(n1009), .Y(n904) );
  MXI2XL U974 ( .A(n902), .B(n903), .S0(n976), .Y(blockdata[18]) );
  MXI4XL U975 ( .A(\block[4][18] ), .B(\block[5][18] ), .C(\block[6][18] ), 
        .D(\block[7][18] ), .S0(n1040), .S1(n1009), .Y(n903) );
  MXI4XL U976 ( .A(\block[0][18] ), .B(\block[1][18] ), .C(\block[2][18] ), 
        .D(\block[3][18] ), .S0(n1041), .S1(n1009), .Y(n902) );
  MXI2XL U977 ( .A(n898), .B(n899), .S0(n976), .Y(blockdata[20]) );
  MXI4XL U978 ( .A(\block[4][20] ), .B(\block[5][20] ), .C(\block[6][20] ), 
        .D(\block[7][20] ), .S0(n1040), .S1(n1009), .Y(n899) );
  MXI4XL U979 ( .A(\block[0][20] ), .B(\block[1][20] ), .C(\block[2][20] ), 
        .D(\block[3][20] ), .S0(n1040), .S1(n1009), .Y(n898) );
  MXI2XL U980 ( .A(n900), .B(n901), .S0(n976), .Y(blockdata[19]) );
  MXI4XL U981 ( .A(\block[4][19] ), .B(\block[5][19] ), .C(\block[6][19] ), 
        .D(\block[7][19] ), .S0(n1040), .S1(n1009), .Y(n901) );
  MXI4XL U982 ( .A(\block[0][19] ), .B(\block[1][19] ), .C(\block[2][19] ), 
        .D(\block[3][19] ), .S0(n1040), .S1(n1009), .Y(n900) );
  MXI2XL U983 ( .A(n876), .B(n877), .S0(n973), .Y(blockdata[50]) );
  MXI4XL U984 ( .A(\block[4][50] ), .B(\block[5][50] ), .C(\block[6][50] ), 
        .D(\block[7][50] ), .S0(n1036), .S1(n1004), .Y(n877) );
  MXI4XL U985 ( .A(\block[0][50] ), .B(\block[1][50] ), .C(\block[2][50] ), 
        .D(\block[3][50] ), .S0(n1036), .S1(n1004), .Y(n876) );
  MXI2XL U986 ( .A(n878), .B(n879), .S0(n973), .Y(blockdata[49]) );
  MXI4XL U987 ( .A(\block[4][49] ), .B(\block[5][49] ), .C(\block[6][49] ), 
        .D(\block[7][49] ), .S0(n1036), .S1(n1004), .Y(n879) );
  MXI4XL U988 ( .A(\block[0][49] ), .B(\block[1][49] ), .C(\block[2][49] ), 
        .D(\block[3][49] ), .S0(n1036), .S1(n1004), .Y(n878) );
  MXI2XL U989 ( .A(n872), .B(n873), .S0(n973), .Y(blockdata[52]) );
  MXI4XL U990 ( .A(\block[4][52] ), .B(\block[5][52] ), .C(\block[6][52] ), 
        .D(\block[7][52] ), .S0(n1035), .S1(n1003), .Y(n873) );
  MXI4XL U991 ( .A(\block[0][52] ), .B(\block[1][52] ), .C(\block[2][52] ), 
        .D(\block[3][52] ), .S0(n1035), .S1(n1003), .Y(n872) );
  MXI2XL U992 ( .A(n868), .B(n869), .S0(n973), .Y(blockdata[54]) );
  MXI4XL U993 ( .A(\block[4][54] ), .B(\block[5][54] ), .C(\block[6][54] ), 
        .D(\block[7][54] ), .S0(n1035), .S1(n1003), .Y(n869) );
  MXI4XL U994 ( .A(\block[0][54] ), .B(\block[1][54] ), .C(\block[2][54] ), 
        .D(\block[3][54] ), .S0(n1035), .S1(n1003), .Y(n868) );
  MXI2XL U995 ( .A(n874), .B(n875), .S0(n973), .Y(blockdata[51]) );
  MXI4XL U996 ( .A(\block[4][51] ), .B(\block[5][51] ), .C(\block[6][51] ), 
        .D(\block[7][51] ), .S0(n1035), .S1(n1003), .Y(n875) );
  MXI4XL U997 ( .A(\block[0][51] ), .B(\block[1][51] ), .C(\block[2][51] ), 
        .D(\block[3][51] ), .S0(n1035), .S1(n1003), .Y(n874) );
  MXI2XL U998 ( .A(n866), .B(n867), .S0(n973), .Y(blockdata[55]) );
  MXI4XL U999 ( .A(\block[4][55] ), .B(\block[5][55] ), .C(\block[6][55] ), 
        .D(\block[7][55] ), .S0(n1035), .S1(n1003), .Y(n867) );
  MXI4XL U1000 ( .A(\block[0][55] ), .B(\block[1][55] ), .C(\block[2][55] ), 
        .D(\block[3][55] ), .S0(n1035), .S1(n1003), .Y(n866) );
  MXI2XL U1001 ( .A(n864), .B(n865), .S0(n973), .Y(blockdata[56]) );
  MXI4XL U1002 ( .A(\block[4][56] ), .B(\block[5][56] ), .C(\block[6][56] ), 
        .D(\block[7][56] ), .S0(n1035), .S1(n1003), .Y(n865) );
  MXI4XL U1003 ( .A(\block[0][56] ), .B(\block[1][56] ), .C(\block[2][56] ), 
        .D(\block[3][56] ), .S0(n1035), .S1(n1003), .Y(n864) );
  MXI2XL U1004 ( .A(n870), .B(n871), .S0(n973), .Y(blockdata[53]) );
  MXI4XL U1005 ( .A(\block[4][53] ), .B(\block[5][53] ), .C(\block[6][53] ), 
        .D(\block[7][53] ), .S0(n1035), .S1(n1003), .Y(n871) );
  MXI4XL U1006 ( .A(\block[0][53] ), .B(\block[1][53] ), .C(\block[2][53] ), 
        .D(\block[3][53] ), .S0(n1035), .S1(n1003), .Y(n870) );
  MXI2XL U1007 ( .A(n880), .B(n881), .S0(n973), .Y(blockdata[48]) );
  MXI4XL U1008 ( .A(\block[4][48] ), .B(\block[5][48] ), .C(\block[6][48] ), 
        .D(\block[7][48] ), .S0(n1036), .S1(n1004), .Y(n881) );
  MXI4XL U1009 ( .A(\block[0][48] ), .B(\block[1][48] ), .C(\block[2][48] ), 
        .D(\block[3][48] ), .S0(n1036), .S1(n1004), .Y(n880) );
  MXI2XL U1010 ( .A(n906), .B(n907), .S0(n976), .Y(blockdata[16]) );
  MXI4XL U1011 ( .A(\block[4][16] ), .B(\block[5][16] ), .C(\block[6][16] ), 
        .D(\block[7][16] ), .S0(n1041), .S1(n1009), .Y(n907) );
  MXI4XL U1012 ( .A(\block[0][16] ), .B(\block[1][16] ), .C(\block[2][16] ), 
        .D(\block[3][16] ), .S0(n1041), .S1(n1009), .Y(n906) );
  MXI2XL U1013 ( .A(n1735), .B(n1537), .S0(n573), .Y(n1719) );
  MXI2XL U1014 ( .A(n1734), .B(n1537), .S0(n567), .Y(n1718) );
  MXI2XL U1015 ( .A(n1733), .B(n1537), .S0(n571), .Y(n1717) );
  MXI2XL U1016 ( .A(n1732), .B(n1537), .S0(n565), .Y(n1716) );
  NAND3BXL U1017 ( .AN(proc_addr[0]), .B(n1302), .C(n1550), .Y(n1470) );
  CLKBUFX3 U1018 ( .A(n1005), .Y(n995) );
  CLKBUFX3 U1019 ( .A(n1098), .Y(n1102) );
  CLKBUFX3 U1020 ( .A(n1097), .Y(n1103) );
  CLKBUFX3 U1021 ( .A(n1098), .Y(n1104) );
  CLKBUFX3 U1022 ( .A(n1098), .Y(n1105) );
  CLKBUFX3 U1023 ( .A(n1098), .Y(n1106) );
  CLKBUFX3 U1024 ( .A(n1098), .Y(n1107) );
  CLKBUFX3 U1025 ( .A(n1097), .Y(n1108) );
  CLKBUFX3 U1026 ( .A(n1097), .Y(n1109) );
  CLKBUFX3 U1027 ( .A(n1097), .Y(n1110) );
  CLKBUFX3 U1028 ( .A(n1112), .Y(n1100) );
  CLKBUFX3 U1029 ( .A(n1112), .Y(n1101) );
  CLKBUFX3 U1030 ( .A(n1187), .Y(n1175) );
  CLKBUFX3 U1031 ( .A(n1187), .Y(n1176) );
  CLKBUFX3 U1032 ( .A(n1186), .Y(n1177) );
  CLKBUFX3 U1033 ( .A(n1186), .Y(n1178) );
  CLKBUFX3 U1034 ( .A(n1185), .Y(n1179) );
  CLKBUFX3 U1035 ( .A(n1185), .Y(n1180) );
  CLKBUFX3 U1036 ( .A(n1170), .Y(n1181) );
  CLKBUFX3 U1037 ( .A(n1170), .Y(n1182) );
  CLKBUFX3 U1038 ( .A(n1188), .Y(n1173) );
  CLKBUFX3 U1039 ( .A(n1188), .Y(n1174) );
  CLKBUFX3 U1040 ( .A(n1149), .Y(n1137) );
  CLKBUFX3 U1041 ( .A(n1149), .Y(n1138) );
  CLKBUFX3 U1042 ( .A(n1148), .Y(n1139) );
  CLKBUFX3 U1043 ( .A(n1148), .Y(n1140) );
  CLKBUFX3 U1044 ( .A(n1147), .Y(n1141) );
  CLKBUFX3 U1045 ( .A(n1147), .Y(n1142) );
  CLKBUFX3 U1046 ( .A(n1132), .Y(n1143) );
  CLKBUFX3 U1047 ( .A(n1132), .Y(n1144) );
  CLKBUFX3 U1048 ( .A(n1150), .Y(n1135) );
  CLKBUFX3 U1049 ( .A(n1150), .Y(n1136) );
  CLKBUFX3 U1050 ( .A(n1225), .Y(n1213) );
  CLKBUFX3 U1051 ( .A(n1225), .Y(n1214) );
  CLKBUFX3 U1052 ( .A(n1224), .Y(n1215) );
  CLKBUFX3 U1053 ( .A(n1224), .Y(n1216) );
  CLKBUFX3 U1054 ( .A(n1223), .Y(n1217) );
  CLKBUFX3 U1055 ( .A(n1223), .Y(n1218) );
  CLKBUFX3 U1056 ( .A(n1208), .Y(n1219) );
  CLKBUFX3 U1057 ( .A(n1208), .Y(n1220) );
  CLKBUFX3 U1058 ( .A(n1226), .Y(n1211) );
  CLKBUFX3 U1059 ( .A(n1226), .Y(n1212) );
  CLKBUFX3 U1060 ( .A(n1097), .Y(n1111) );
  CLKBUFX3 U1061 ( .A(n1170), .Y(n1184) );
  CLKBUFX3 U1062 ( .A(n1132), .Y(n1146) );
  CLKBUFX3 U1063 ( .A(n1208), .Y(n1222) );
  CLKBUFX3 U1064 ( .A(n1248), .Y(n972) );
  CLKBUFX3 U1065 ( .A(n964), .Y(n975) );
  CLKBUFX3 U1066 ( .A(n1248), .Y(n969) );
  CLKBUFX3 U1067 ( .A(n964), .Y(n970) );
  CLKBUFX3 U1068 ( .A(n1017), .Y(n1031) );
  CLKBUFX3 U1069 ( .A(n1021), .Y(n1039) );
  CLKBUFX3 U1070 ( .A(n1021), .Y(n1038) );
  CLKBUFX3 U1071 ( .A(n1025), .Y(n1027) );
  CLKBUFX3 U1072 ( .A(n1025), .Y(n1026) );
  CLKBUFX3 U1073 ( .A(n983), .Y(n988) );
  CLKBUFX3 U1074 ( .A(n965), .Y(n974) );
  CLKBUFX3 U1075 ( .A(n966), .Y(n971) );
  CLKBUFX3 U1076 ( .A(n964), .Y(n976) );
  CLKBUFX3 U1077 ( .A(n965), .Y(n973) );
  CLKBUFX3 U1078 ( .A(n1020), .Y(n1030) );
  CLKBUFX3 U1079 ( .A(n1019), .Y(n1042) );
  CLKBUFX3 U1080 ( .A(n1023), .Y(n1034) );
  CLKBUFX3 U1081 ( .A(n1020), .Y(n1037) );
  CLKBUFX3 U1082 ( .A(n1024), .Y(n1029) );
  CLKBUFX3 U1083 ( .A(n1020), .Y(n1041) );
  CLKBUFX3 U1084 ( .A(n1024), .Y(n1036) );
  CLKBUFX3 U1085 ( .A(n1020), .Y(n1033) );
  CLKBUFX3 U1086 ( .A(n1024), .Y(n1028) );
  CLKBUFX3 U1087 ( .A(n1022), .Y(n1035) );
  CLKBUFX3 U1088 ( .A(n1020), .Y(n1040) );
  CLKBUFX3 U1089 ( .A(n1020), .Y(n1032) );
  CLKBUFX3 U1090 ( .A(n983), .Y(n989) );
  CLKBUFX3 U1091 ( .A(n1131), .Y(n1117) );
  CLKBUFX3 U1092 ( .A(n1131), .Y(n1118) );
  CLKBUFX3 U1093 ( .A(n1130), .Y(n1119) );
  CLKBUFX3 U1094 ( .A(n1130), .Y(n1120) );
  CLKBUFX3 U1095 ( .A(n1129), .Y(n1121) );
  CLKBUFX3 U1096 ( .A(n1129), .Y(n1122) );
  CLKBUFX3 U1097 ( .A(n1128), .Y(n1123) );
  CLKBUFX3 U1098 ( .A(n1128), .Y(n1124) );
  CLKBUFX3 U1099 ( .A(n1127), .Y(n1125) );
  CLKBUFX3 U1100 ( .A(n1131), .Y(n1115) );
  CLKBUFX3 U1101 ( .A(n1131), .Y(n1116) );
  CLKBUFX3 U1102 ( .A(n1206), .Y(n1194) );
  CLKBUFX3 U1103 ( .A(n1206), .Y(n1195) );
  CLKBUFX3 U1104 ( .A(n1205), .Y(n1196) );
  CLKBUFX3 U1105 ( .A(n1205), .Y(n1197) );
  CLKBUFX3 U1106 ( .A(n1204), .Y(n1198) );
  CLKBUFX3 U1107 ( .A(n1204), .Y(n1199) );
  CLKBUFX3 U1108 ( .A(n1189), .Y(n1200) );
  CLKBUFX3 U1109 ( .A(n1189), .Y(n1201) );
  CLKBUFX3 U1110 ( .A(n1207), .Y(n1192) );
  CLKBUFX3 U1111 ( .A(n1207), .Y(n1193) );
  CLKBUFX3 U1112 ( .A(n1168), .Y(n1156) );
  CLKBUFX3 U1113 ( .A(n1168), .Y(n1157) );
  CLKBUFX3 U1114 ( .A(n1167), .Y(n1158) );
  CLKBUFX3 U1115 ( .A(n1167), .Y(n1159) );
  CLKBUFX3 U1116 ( .A(n1166), .Y(n1160) );
  CLKBUFX3 U1117 ( .A(n1166), .Y(n1161) );
  CLKBUFX3 U1118 ( .A(n1151), .Y(n1162) );
  CLKBUFX3 U1119 ( .A(n1151), .Y(n1163) );
  CLKBUFX3 U1120 ( .A(n1169), .Y(n1154) );
  CLKBUFX3 U1121 ( .A(n1169), .Y(n1155) );
  CLKBUFX3 U1122 ( .A(n1244), .Y(n1232) );
  CLKBUFX3 U1123 ( .A(n1244), .Y(n1233) );
  CLKBUFX3 U1124 ( .A(n1243), .Y(n1234) );
  CLKBUFX3 U1125 ( .A(n1243), .Y(n1235) );
  CLKBUFX3 U1126 ( .A(n1242), .Y(n1236) );
  CLKBUFX3 U1127 ( .A(n1242), .Y(n1237) );
  CLKBUFX3 U1128 ( .A(n1227), .Y(n1238) );
  CLKBUFX3 U1129 ( .A(n1227), .Y(n1239) );
  CLKBUFX3 U1130 ( .A(n1245), .Y(n1230) );
  CLKBUFX3 U1131 ( .A(n1245), .Y(n1231) );
  CLKBUFX3 U1132 ( .A(n1127), .Y(n1126) );
  CLKBUFX3 U1133 ( .A(n1189), .Y(n1203) );
  CLKBUFX3 U1134 ( .A(n1151), .Y(n1165) );
  CLKBUFX3 U1135 ( .A(n1227), .Y(n1241) );
  CLKBUFX3 U1136 ( .A(n1171), .Y(n1186) );
  CLKBUFX3 U1137 ( .A(n1171), .Y(n1185) );
  CLKBUFX3 U1138 ( .A(n1133), .Y(n1148) );
  CLKBUFX3 U1139 ( .A(n1133), .Y(n1147) );
  CLKBUFX3 U1140 ( .A(n1209), .Y(n1224) );
  CLKBUFX3 U1141 ( .A(n1209), .Y(n1223) );
  CLKBUFX6 U1142 ( .A(n1753), .Y(mem_write) );
  CLKBUFX3 U1143 ( .A(n966), .Y(n968) );
  CLKBUFX3 U1144 ( .A(n1080), .Y(n1071) );
  CLKBUFX3 U1145 ( .A(n1079), .Y(n1074) );
  CLKBUFX3 U1146 ( .A(n554), .Y(n1098) );
  CLKBUFX3 U1147 ( .A(n554), .Y(n1099) );
  CLKBUFX3 U1148 ( .A(n554), .Y(n1097) );
  CLKBUFX3 U1149 ( .A(n555), .Y(n1171) );
  CLKBUFX3 U1150 ( .A(n555), .Y(n1172) );
  CLKBUFX3 U1151 ( .A(n556), .Y(n1133) );
  CLKBUFX3 U1152 ( .A(n556), .Y(n1134) );
  CLKBUFX3 U1153 ( .A(n555), .Y(n1170) );
  CLKBUFX3 U1154 ( .A(n556), .Y(n1132) );
  CLKBUFX3 U1155 ( .A(n557), .Y(n1209) );
  CLKBUFX3 U1156 ( .A(n557), .Y(n1210) );
  CLKBUFX3 U1157 ( .A(n557), .Y(n1208) );
  CLKBUFX3 U1158 ( .A(n1114), .Y(n1130) );
  CLKBUFX3 U1159 ( .A(n1114), .Y(n1129) );
  CLKBUFX3 U1160 ( .A(n1113), .Y(n1128) );
  CLKBUFX3 U1161 ( .A(n1113), .Y(n1127) );
  CLKBUFX3 U1162 ( .A(n1190), .Y(n1205) );
  CLKBUFX3 U1163 ( .A(n1190), .Y(n1204) );
  CLKBUFX3 U1164 ( .A(n1152), .Y(n1167) );
  CLKBUFX3 U1165 ( .A(n1152), .Y(n1166) );
  CLKBUFX3 U1166 ( .A(n1228), .Y(n1243) );
  CLKBUFX3 U1167 ( .A(n1228), .Y(n1242) );
  CLKBUFX3 U1168 ( .A(n1048), .Y(n1017) );
  BUFX12 U1169 ( .A(n1371), .Y(n1055) );
  CLKBUFX3 U1170 ( .A(n1048), .Y(n1015) );
  CLKBUFX3 U1171 ( .A(n980), .Y(n991) );
  CLKBUFX3 U1172 ( .A(n1753), .Y(n1251) );
  CLKINVX1 U1173 ( .A(proc_read), .Y(n1049) );
  CLKBUFX3 U1174 ( .A(n560), .Y(n1114) );
  CLKBUFX3 U1175 ( .A(n560), .Y(n1113) );
  CLKBUFX3 U1176 ( .A(n561), .Y(n1190) );
  CLKBUFX3 U1177 ( .A(n561), .Y(n1191) );
  CLKBUFX3 U1178 ( .A(n562), .Y(n1152) );
  CLKBUFX3 U1179 ( .A(n562), .Y(n1153) );
  CLKBUFX3 U1180 ( .A(n561), .Y(n1189) );
  CLKBUFX3 U1181 ( .A(n562), .Y(n1151) );
  CLKBUFX3 U1182 ( .A(n563), .Y(n1228) );
  CLKBUFX3 U1183 ( .A(n563), .Y(n1229) );
  CLKBUFX3 U1184 ( .A(n563), .Y(n1227) );
  CLKBUFX3 U1185 ( .A(n1260), .Y(n1258) );
  CLKBUFX3 U1186 ( .A(n1336), .Y(n1053) );
  CLKBUFX3 U1187 ( .A(n1336), .Y(n1052) );
  CLKBUFX3 U1188 ( .A(n1372), .Y(n1056) );
  BUFX20 U1189 ( .A(n1090), .Y(n1092) );
  OAI221X1 U1190 ( .A0(n1094), .A1(n1556), .B0(n1091), .B1(n1555), .C0(n1554), 
        .Y(proc_rdata[0]) );
  OA22X1 U1191 ( .A0(n1087), .A1(n1553), .B0(n1083), .B1(n1552), .Y(n1554) );
  OAI221X1 U1192 ( .A0(n1094), .A1(n1601), .B0(n1091), .B1(n1600), .C0(n1599), 
        .Y(proc_rdata[9]) );
  OA22X1 U1193 ( .A0(n1087), .A1(n1598), .B0(n1083), .B1(n1597), .Y(n1599) );
  OAI221X1 U1194 ( .A0(n1095), .A1(n1616), .B0(n1091), .B1(n1615), .C0(n1614), 
        .Y(proc_rdata[12]) );
  OAI221X1 U1195 ( .A0(n1095), .A1(n1621), .B0(n1091), .B1(n1620), .C0(n1619), 
        .Y(proc_rdata[13]) );
  OA22X1 U1196 ( .A0(n1088), .A1(n1618), .B0(n1084), .B1(n1617), .Y(n1619) );
  OAI221X1 U1197 ( .A0(n1094), .A1(n1606), .B0(n1091), .B1(n1605), .C0(n1604), 
        .Y(proc_rdata[10]) );
  OA22X1 U1198 ( .A0(n1087), .A1(n1603), .B0(n1083), .B1(n1602), .Y(n1604) );
  OAI221XL U1199 ( .A0(n1095), .A1(n1646), .B0(n1091), .B1(n1645), .C0(n1644), 
        .Y(proc_rdata[18]) );
  OAI221XL U1200 ( .A0(n1095), .A1(n1656), .B0(n1091), .B1(n1655), .C0(n1654), 
        .Y(proc_rdata[20]) );
  OAI221XL U1201 ( .A0(n1095), .A1(n1666), .B0(n1091), .B1(n1665), .C0(n1664), 
        .Y(proc_rdata[22]) );
  OAI221XL U1202 ( .A0(n1095), .A1(n1641), .B0(n1091), .B1(n1640), .C0(n1639), 
        .Y(proc_rdata[17]) );
  OAI221XL U1203 ( .A0(n1095), .A1(n1651), .B0(n1091), .B1(n1650), .C0(n1649), 
        .Y(proc_rdata[19]) );
  OAI221XL U1204 ( .A0(n1095), .A1(n1661), .B0(n1091), .B1(n1660), .C0(n1659), 
        .Y(proc_rdata[21]) );
  OAI221XL U1205 ( .A0(n1095), .A1(n1671), .B0(n1091), .B1(n1670), .C0(n1669), 
        .Y(proc_rdata[23]) );
  OAI221XL U1206 ( .A0(n1096), .A1(n1681), .B0(n1092), .B1(n1680), .C0(n1679), 
        .Y(proc_rdata[25]) );
  OA22X1 U1207 ( .A0(n1089), .A1(n1678), .B0(n1085), .B1(n1677), .Y(n1679) );
  OAI221XL U1208 ( .A0(n1096), .A1(n1676), .B0(n1092), .B1(n1675), .C0(n1674), 
        .Y(proc_rdata[24]) );
  OA22X1 U1209 ( .A0(n1089), .A1(n1673), .B0(n1085), .B1(n1672), .Y(n1674) );
  OAI221XL U1210 ( .A0(n1095), .A1(n1636), .B0(n1091), .B1(n1635), .C0(n1634), 
        .Y(proc_rdata[16]) );
  NAND3BX1 U1211 ( .AN(n1062), .B(n568), .C(n1470), .Y(n1338) );
  NAND2XL U1212 ( .A(n1540), .B(n1303), .Y(n1472) );
  AND2X2 U1213 ( .A(n568), .B(n1057), .Y(n558) );
  OAI221X1 U1214 ( .A0(n1094), .A1(n1586), .B0(n1091), .B1(n1585), .C0(n1584), 
        .Y(proc_rdata[6]) );
  OA22X1 U1215 ( .A0(n1087), .A1(n1583), .B0(n1083), .B1(n1582), .Y(n1584) );
  OAI221X1 U1216 ( .A0(n1095), .A1(n1626), .B0(n1091), .B1(n1625), .C0(n1624), 
        .Y(proc_rdata[14]) );
  OA22X1 U1217 ( .A0(n1088), .A1(n1623), .B0(n1084), .B1(n1622), .Y(n1624) );
  OAI221X1 U1218 ( .A0(n1094), .A1(n1611), .B0(n1091), .B1(n1610), .C0(n1609), 
        .Y(proc_rdata[11]) );
  OA22X1 U1219 ( .A0(n1087), .A1(n1608), .B0(n1083), .B1(n1607), .Y(n1609) );
  OAI221X1 U1220 ( .A0(n1095), .A1(n1631), .B0(n1091), .B1(n1630), .C0(n1629), 
        .Y(proc_rdata[15]) );
  OA22X1 U1221 ( .A0(n1088), .A1(n1628), .B0(n1084), .B1(n1627), .Y(n1629) );
  CLKBUFX3 U1222 ( .A(n1470), .Y(n1065) );
  CLKBUFX3 U1223 ( .A(n1470), .Y(n1066) );
  CLKBUFX3 U1224 ( .A(n1372), .Y(n1057) );
  BUFX20 U1225 ( .A(n1093), .Y(n1096) );
  BUFX20 U1226 ( .A(n1086), .Y(n1089) );
  BUFX20 U1227 ( .A(n1082), .Y(n1085) );
  NAND2XL U1228 ( .A(dirty), .B(valid), .Y(n1542) );
  NAND4BXL U1229 ( .AN(n1542), .B(n1541), .C(n1540), .D(n1539), .Y(n1543) );
  CLKINVX1 U1230 ( .A(n1545), .Y(n1752) );
  CLKINVX1 U1231 ( .A(blockdata[123]), .Y(n1690) );
  CLKINVX1 U1232 ( .A(blockdata[61]), .Y(n1697) );
  CLKINVX1 U1233 ( .A(blockdata[93]), .Y(n1698) );
  CLKINVX1 U1234 ( .A(blockdata[14]), .Y(n1626) );
  CLKINVX1 U1235 ( .A(blockdata[15]), .Y(n1631) );
  CLKINVX1 U1236 ( .A(blockdata[111]), .Y(n1630) );
  CLKINVX1 U1237 ( .A(blockdata[34]), .Y(n1562) );
  CLKINVX1 U1238 ( .A(blockdata[35]), .Y(n1567) );
  CLKINVX1 U1239 ( .A(blockdata[33]), .Y(n1557) );
  CLKINVX1 U1240 ( .A(blockdata[37]), .Y(n1577) );
  CLKINVX1 U1241 ( .A(blockdata[39]), .Y(n1587) );
  CLKINVX1 U1242 ( .A(blockdata[38]), .Y(n1582) );
  CLKINVX1 U1243 ( .A(blockdata[40]), .Y(n1592) );
  CLKINVX1 U1244 ( .A(blockdata[46]), .Y(n1622) );
  CLKINVX1 U1245 ( .A(blockdata[69]), .Y(n1578) );
  CLKINVX1 U1246 ( .A(blockdata[71]), .Y(n1588) );
  CLKINVX1 U1247 ( .A(blockdata[70]), .Y(n1583) );
  CLKINVX1 U1248 ( .A(blockdata[72]), .Y(n1593) );
  AND2X2 U1249 ( .A(n1474), .B(n1473), .Y(n1538) );
  OAI21XL U1250 ( .A0(n1539), .A1(n1472), .B0(dirty), .Y(n1474) );
  AND2X2 U1251 ( .A(n1748), .B(n1246), .Y(n570) );
  CLKINVX1 U1252 ( .A(blockdata[18]), .Y(n1646) );
  CLKINVX1 U1253 ( .A(blockdata[20]), .Y(n1656) );
  CLKINVX1 U1254 ( .A(blockdata[17]), .Y(n1641) );
  CLKINVX1 U1255 ( .A(blockdata[19]), .Y(n1651) );
  CLKINVX1 U1256 ( .A(blockdata[114]), .Y(n1645) );
  CLKINVX1 U1257 ( .A(blockdata[113]), .Y(n1640) );
  CLKINVX1 U1258 ( .A(blockdata[115]), .Y(n1650) );
  CLKINVX1 U1259 ( .A(blockdata[112]), .Y(n1635) );
  CLKINVX1 U1260 ( .A(blockdata[16]), .Y(n1636) );
  CLKINVX1 U1261 ( .A(blockdata[50]), .Y(n1642) );
  CLKINVX1 U1262 ( .A(blockdata[52]), .Y(n1652) );
  CLKINVX1 U1263 ( .A(blockdata[54]), .Y(n1662) );
  CLKINVX1 U1264 ( .A(blockdata[49]), .Y(n1637) );
  CLKINVX1 U1265 ( .A(blockdata[51]), .Y(n1647) );
  CLKINVX1 U1266 ( .A(blockdata[53]), .Y(n1657) );
  CLKINVX1 U1267 ( .A(blockdata[55]), .Y(n1667) );
  CLKINVX1 U1268 ( .A(blockdata[56]), .Y(n1672) );
  CLKINVX1 U1269 ( .A(blockdata[48]), .Y(n1632) );
  CLKINVX1 U1270 ( .A(blockdata[80]), .Y(n1633) );
  NOR2X1 U1271 ( .A(n1249), .B(n1247), .Y(n1751) );
  NOR2XL U1272 ( .A(n1247), .B(n1248), .Y(n1749) );
  NOR2XL U1273 ( .A(n1249), .B(N32), .Y(n1750) );
  AND2X2 U1274 ( .A(n1751), .B(n1246), .Y(n571) );
  AND2X2 U1275 ( .A(n1749), .B(n1246), .Y(n572) );
  AND2X2 U1276 ( .A(n1750), .B(n1246), .Y(n573) );
  CLKINVX1 U1277 ( .A(n1473), .Y(n1302) );
  CLKINVX1 U1278 ( .A(n1405), .Y(n1062) );
  NAND3BXL U1279 ( .AN(n1549), .B(n1302), .C(n1550), .Y(n1405) );
  CLKMX2X4 U1280 ( .A(n612), .B(n613), .S0(n978), .Y(tag[23]) );
  MX4X1 U1281 ( .A(\blocktag[0][23] ), .B(\blocktag[1][23] ), .C(
        \blocktag[2][23] ), .D(\blocktag[3][23] ), .S0(n1044), .S1(n983), .Y(
        n612) );
  MX4X1 U1282 ( .A(\blocktag[4][23] ), .B(\blocktag[5][23] ), .C(
        \blocktag[6][23] ), .D(\blocktag[7][23] ), .S0(n1044), .S1(n983), .Y(
        n613) );
  MX4X1 U1283 ( .A(\blocktag[0][19] ), .B(\blocktag[1][19] ), .C(
        \blocktag[2][19] ), .D(\blocktag[3][19] ), .S0(n1045), .S1(n983), .Y(
        n616) );
  MX4X1 U1284 ( .A(\blocktag[4][19] ), .B(\blocktag[5][19] ), .C(
        \blocktag[6][19] ), .D(\blocktag[7][19] ), .S0(n1044), .S1(n983), .Y(
        n617) );
  NAND2XL U1285 ( .A(mem_rdata[9]), .B(n1070), .Y(n1450) );
  NAND2XL U1286 ( .A(mem_rdata[10]), .B(n1070), .Y(n1448) );
  NAND2XL U1287 ( .A(mem_rdata[11]), .B(n1070), .Y(n1446) );
  NAND2XL U1288 ( .A(mem_rdata[12]), .B(n1070), .Y(n1444) );
  NAND2XL U1289 ( .A(mem_rdata[13]), .B(n1070), .Y(n1442) );
  NAND2XL U1290 ( .A(mem_rdata[15]), .B(n1071), .Y(n1438) );
  NAND2XL U1291 ( .A(mem_rdata[16]), .B(n1071), .Y(n1436) );
  NAND2XL U1292 ( .A(mem_rdata[17]), .B(n1071), .Y(n1434) );
  NAND2XL U1293 ( .A(mem_rdata[18]), .B(n1071), .Y(n1432) );
  NAND2XL U1294 ( .A(mem_rdata[19]), .B(n1071), .Y(n1430) );
  NAND2XL U1295 ( .A(mem_rdata[20]), .B(n1071), .Y(n1428) );
  NAND2XL U1296 ( .A(mem_rdata[21]), .B(n1071), .Y(n1426) );
  NAND2XL U1297 ( .A(mem_rdata[22]), .B(n1071), .Y(n1424) );
  NAND2XL U1298 ( .A(mem_rdata[23]), .B(n1071), .Y(n1422) );
  NAND2XL U1299 ( .A(mem_rdata[24]), .B(n1071), .Y(n1420) );
  NAND2XL U1300 ( .A(mem_rdata[25]), .B(n1071), .Y(n1418) );
  NAND2XL U1301 ( .A(mem_rdata[26]), .B(n1071), .Y(n1416) );
  NAND2XL U1302 ( .A(mem_rdata[28]), .B(n1070), .Y(n1412) );
  NAND2XL U1303 ( .A(mem_rdata[29]), .B(n1070), .Y(n1410) );
  NAND2XL U1304 ( .A(mem_rdata[30]), .B(n1070), .Y(n1408) );
  NAND2XL U1305 ( .A(mem_rdata[31]), .B(n1070), .Y(n1406) );
  NAND2XL U1306 ( .A(mem_rdata[1]), .B(n1070), .Y(n1466) );
  NAND2XL U1307 ( .A(mem_rdata[2]), .B(n1070), .Y(n1464) );
  NAND2XL U1308 ( .A(mem_rdata[4]), .B(n1070), .Y(n1460) );
  NAND2XL U1309 ( .A(mem_rdata[5]), .B(n1070), .Y(n1458) );
  NAND2XL U1310 ( .A(mem_rdata[6]), .B(n1070), .Y(n1456) );
  NAND2XL U1311 ( .A(mem_rdata[7]), .B(n1070), .Y(n1454) );
  NAND2XL U1312 ( .A(mem_rdata[41]), .B(n1072), .Y(n1395) );
  NAND2XL U1313 ( .A(mem_rdata[42]), .B(n1072), .Y(n1394) );
  NAND2XL U1314 ( .A(mem_rdata[43]), .B(n1072), .Y(n1393) );
  NAND2XL U1315 ( .A(mem_rdata[44]), .B(n1072), .Y(n1392) );
  NAND2XL U1316 ( .A(mem_rdata[45]), .B(n1072), .Y(n1391) );
  NAND2XL U1317 ( .A(mem_rdata[47]), .B(n1072), .Y(n1389) );
  NAND2XL U1318 ( .A(mem_rdata[54]), .B(n1077), .Y(n1382) );
  NAND2XL U1319 ( .A(mem_rdata[55]), .B(n1077), .Y(n1381) );
  NAND2XL U1320 ( .A(mem_rdata[56]), .B(n1077), .Y(n1380) );
  NAND2XL U1321 ( .A(mem_rdata[57]), .B(n1077), .Y(n1379) );
  NAND2XL U1322 ( .A(mem_rdata[58]), .B(n1077), .Y(n1378) );
  NAND2XL U1323 ( .A(mem_rdata[60]), .B(n1075), .Y(n1376) );
  NAND2XL U1324 ( .A(mem_rdata[63]), .B(n1075), .Y(n1373) );
  NAND2XL U1325 ( .A(mem_rdata[32]), .B(n1070), .Y(n1404) );
  NAND2XL U1326 ( .A(mem_rdata[33]), .B(n1070), .Y(n1403) );
  NAND2XL U1327 ( .A(mem_rdata[34]), .B(n1077), .Y(n1402) );
  NAND2XL U1328 ( .A(mem_rdata[35]), .B(n1070), .Y(n1401) );
  NAND2XL U1329 ( .A(mem_rdata[36]), .B(n1070), .Y(n1400) );
  NAND2XL U1330 ( .A(mem_rdata[37]), .B(n1070), .Y(n1399) );
  NAND2XL U1331 ( .A(mem_rdata[38]), .B(n1070), .Y(n1398) );
  NAND2XL U1332 ( .A(mem_rdata[39]), .B(n1070), .Y(n1397) );
  NAND2XL U1333 ( .A(mem_rdata[74]), .B(n1073), .Y(n1360) );
  NAND2XL U1334 ( .A(mem_rdata[75]), .B(n1073), .Y(n1359) );
  NAND2XL U1335 ( .A(mem_rdata[76]), .B(n1073), .Y(n1358) );
  NAND2XL U1336 ( .A(mem_rdata[77]), .B(n1073), .Y(n1357) );
  NAND2XL U1337 ( .A(mem_rdata[78]), .B(n1073), .Y(n1356) );
  NAND2XL U1338 ( .A(mem_rdata[80]), .B(n1074), .Y(n1354) );
  NAND2XL U1339 ( .A(mem_rdata[81]), .B(n1074), .Y(n1353) );
  NAND2XL U1340 ( .A(mem_rdata[82]), .B(n1074), .Y(n1352) );
  NAND2XL U1341 ( .A(mem_rdata[83]), .B(n1074), .Y(n1351) );
  NAND2XL U1342 ( .A(mem_rdata[84]), .B(n1074), .Y(n1350) );
  NAND2XL U1343 ( .A(mem_rdata[85]), .B(n1074), .Y(n1349) );
  NAND2XL U1344 ( .A(mem_rdata[86]), .B(n1074), .Y(n1348) );
  NAND2XL U1345 ( .A(mem_rdata[87]), .B(n1074), .Y(n1347) );
  NAND2XL U1346 ( .A(mem_rdata[88]), .B(n1074), .Y(n1346) );
  NAND2XL U1347 ( .A(mem_rdata[89]), .B(n1074), .Y(n1345) );
  NAND2XL U1348 ( .A(mem_rdata[93]), .B(n1075), .Y(n1341) );
  NAND2XL U1349 ( .A(mem_rdata[94]), .B(n1075), .Y(n1340) );
  NAND2XL U1350 ( .A(mem_rdata[95]), .B(n1075), .Y(n1339) );
  NAND2XL U1351 ( .A(mem_rdata[64]), .B(n1075), .Y(n1370) );
  NAND2XL U1352 ( .A(mem_rdata[65]), .B(n1077), .Y(n1369) );
  OAI211XL U1353 ( .A0(mem_ready), .A1(valid), .B0(n1300), .C0(n1540), .Y(
        n1301) );
  AOI2BB1XL U1354 ( .A0N(n1299), .A1N(n739), .B0(n1547), .Y(n1300) );
  NAND3BXL U1355 ( .AN(mem_ready), .B(proc_stall), .C(n1542), .Y(n1545) );
  CLKMX2X4 U1356 ( .A(n668), .B(n669), .S0(n970), .Y(blockdata[91]) );
  CLKMX2X4 U1357 ( .A(n670), .B(n671), .S0(n975), .Y(blockdata[27]) );
  CLKMX2X4 U1358 ( .A(n672), .B(n673), .S0(n972), .Y(blockdata[58]) );
  CLKMX2X4 U1359 ( .A(n674), .B(n675), .S0(n970), .Y(blockdata[90]) );
  CLKMX2X4 U1360 ( .A(n676), .B(n677), .S0(n975), .Y(blockdata[26]) );
  CLKMX2X2 U1361 ( .A(n678), .B(n679), .S0(n972), .Y(blockdata[62]) );
  MX4X1 U1362 ( .A(\block[4][62] ), .B(\block[5][62] ), .C(\block[6][62] ), 
        .D(\block[7][62] ), .S0(n1022), .S1(n1002), .Y(n679) );
  MX4X1 U1363 ( .A(\block[0][29] ), .B(\block[1][29] ), .C(\block[2][29] ), 
        .D(\block[3][29] ), .S0(n1039), .S1(n1007), .Y(n680) );
  MX4X1 U1364 ( .A(\block[4][29] ), .B(\block[5][29] ), .C(\block[6][29] ), 
        .D(\block[7][29] ), .S0(n1039), .S1(n1007), .Y(n681) );
  MX4X1 U1365 ( .A(\block[0][93] ), .B(\block[1][93] ), .C(\block[2][93] ), 
        .D(\block[3][93] ), .S0(n1031), .S1(n997), .Y(n682) );
  MX4X1 U1366 ( .A(\block[4][93] ), .B(\block[5][93] ), .C(\block[6][93] ), 
        .D(\block[7][93] ), .S0(n1031), .S1(n997), .Y(n683) );
  CLKMX2X2 U1367 ( .A(n684), .B(n685), .S0(n975), .Y(blockdata[30]) );
  MX4X1 U1368 ( .A(\block[0][30] ), .B(\block[1][30] ), .C(\block[2][30] ), 
        .D(\block[3][30] ), .S0(n1039), .S1(n1007), .Y(n684) );
  MX4X1 U1369 ( .A(\block[4][30] ), .B(\block[5][30] ), .C(\block[6][30] ), 
        .D(\block[7][30] ), .S0(n1039), .S1(n1007), .Y(n685) );
  CLKMX2X2 U1370 ( .A(n686), .B(n687), .S0(n969), .Y(blockdata[94]) );
  MX4X1 U1371 ( .A(\block[0][125] ), .B(\block[1][125] ), .C(\block[2][125] ), 
        .D(\block[3][125] ), .S0(n1026), .S1(n992), .Y(n688) );
  CLKMX2X2 U1372 ( .A(n690), .B(n691), .S0(n967), .Y(blockdata[126]) );
  CLKMX2X4 U1373 ( .A(n693), .B(n694), .S0(n967), .Y(blockdata[122]) );
  MX4XL U1374 ( .A(\block[4][122] ), .B(\block[5][122] ), .C(\block[6][122] ), 
        .D(\block[7][122] ), .S0(n1026), .S1(n993), .Y(n694) );
  CLKMX2X4 U1375 ( .A(n695), .B(n696), .S0(n972), .Y(blockdata[59]) );
  MX4X1 U1376 ( .A(\block[0][61] ), .B(\block[1][61] ), .C(\block[2][61] ), 
        .D(\block[3][61] ), .S0(n1022), .S1(n1002), .Y(n697) );
  MX4X1 U1377 ( .A(\block[4][61] ), .B(\block[5][61] ), .C(\block[6][61] ), 
        .D(\block[7][61] ), .S0(n1022), .S1(n1002), .Y(n698) );
  NAND2XL U1378 ( .A(mem_rdata[104]), .B(n1075), .Y(n1327) );
  NAND2XL U1379 ( .A(mem_rdata[106]), .B(n1076), .Y(n1325) );
  NAND2XL U1380 ( .A(mem_rdata[107]), .B(n1076), .Y(n1324) );
  NAND2XL U1381 ( .A(mem_rdata[108]), .B(n1076), .Y(n1323) );
  NAND2XL U1382 ( .A(mem_rdata[109]), .B(n1076), .Y(n1322) );
  NAND2XL U1383 ( .A(mem_rdata[110]), .B(n1076), .Y(n1321) );
  NAND2XL U1384 ( .A(mem_rdata[111]), .B(n1076), .Y(n1320) );
  NAND2XL U1385 ( .A(mem_rdata[112]), .B(n1076), .Y(n1319) );
  NAND2XL U1386 ( .A(mem_rdata[113]), .B(n1076), .Y(n1318) );
  NAND2XL U1387 ( .A(mem_rdata[114]), .B(n1076), .Y(n1317) );
  NAND2XL U1388 ( .A(mem_rdata[115]), .B(n1076), .Y(n1316) );
  NAND2XL U1389 ( .A(mem_rdata[116]), .B(n1076), .Y(n1315) );
  NAND2XL U1390 ( .A(mem_rdata[117]), .B(n1076), .Y(n1314) );
  NAND2XL U1391 ( .A(mem_rdata[119]), .B(n1077), .Y(n1312) );
  NAND2XL U1392 ( .A(mem_rdata[120]), .B(n1077), .Y(n1311) );
  NAND2XL U1393 ( .A(mem_rdata[121]), .B(n1077), .Y(n1310) );
  NAND2XL U1394 ( .A(mem_rdata[96]), .B(n1075), .Y(n1335) );
  NAND2XL U1395 ( .A(mem_rdata[97]), .B(n1075), .Y(n1334) );
  NAND2XL U1396 ( .A(mem_rdata[98]), .B(n1075), .Y(n1333) );
  NAND2XL U1397 ( .A(mem_rdata[99]), .B(n1075), .Y(n1332) );
  NAND2XL U1398 ( .A(mem_rdata[100]), .B(n1075), .Y(n1331) );
  NAND2XL U1399 ( .A(mem_rdata[101]), .B(n1075), .Y(n1330) );
  NAND2XL U1400 ( .A(mem_rdata[102]), .B(n1075), .Y(n1329) );
  NAND2XL U1401 ( .A(mem_rdata[103]), .B(n1075), .Y(n1328) );
  MXI2X1 U1402 ( .A(n926), .B(n927), .S0(n977), .Y(dirty) );
  MXI4XL U1403 ( .A(blockdirty[4]), .B(blockdirty[5]), .C(blockdirty[6]), .D(
        blockdirty[7]), .S0(n1044), .S1(n1011), .Y(n927) );
  MXI4XL U1404 ( .A(blockdirty[0]), .B(blockdirty[1]), .C(blockdirty[2]), .D(
        blockdirty[3]), .S0(n1044), .S1(n1011), .Y(n926) );
  MX4XL U1405 ( .A(\block[0][34] ), .B(\block[1][34] ), .C(\block[2][34] ), 
        .D(\block[3][34] ), .S0(n1038), .S1(n1006), .Y(n699) );
  MX4XL U1406 ( .A(\block[4][34] ), .B(\block[5][34] ), .C(\block[6][34] ), 
        .D(\block[7][34] ), .S0(n1038), .S1(n1006), .Y(n700) );
  MX4XL U1407 ( .A(\block[0][35] ), .B(\block[1][35] ), .C(\block[2][35] ), 
        .D(\block[3][35] ), .S0(n1038), .S1(n1006), .Y(n701) );
  MX4XL U1408 ( .A(\block[4][35] ), .B(\block[5][35] ), .C(\block[6][35] ), 
        .D(\block[7][35] ), .S0(n1038), .S1(n1006), .Y(n702) );
  MXI2XL U1409 ( .A(n850), .B(n851), .S0(n972), .Y(blockdata[67]) );
  MXI4XL U1410 ( .A(\block[0][67] ), .B(\block[1][67] ), .C(\block[2][67] ), 
        .D(\block[3][67] ), .S0(n1022), .S1(N32), .Y(n850) );
  MXI4XL U1411 ( .A(\block[4][67] ), .B(\block[5][67] ), .C(\block[6][67] ), 
        .D(\block[7][67] ), .S0(n1022), .S1(n1004), .Y(n851) );
  MX2XL U1412 ( .A(n703), .B(n704), .S0(n969), .Y(blockdata[99]) );
  MXI2XL U1413 ( .A(n854), .B(n855), .S0(n972), .Y(blockdata[65]) );
  MXI4XL U1414 ( .A(\block[0][65] ), .B(\block[1][65] ), .C(\block[2][65] ), 
        .D(\block[3][65] ), .S0(n1022), .S1(n993), .Y(n854) );
  MXI4XL U1415 ( .A(\block[4][65] ), .B(\block[5][65] ), .C(\block[6][65] ), 
        .D(\block[7][65] ), .S0(n1022), .S1(n1005), .Y(n855) );
  MXI2XL U1416 ( .A(n820), .B(n821), .S0(n969), .Y(blockdata[97]) );
  MXI4XL U1417 ( .A(\block[0][97] ), .B(\block[1][97] ), .C(\block[2][97] ), 
        .D(\block[3][97] ), .S0(n1030), .S1(n997), .Y(n820) );
  MXI4XL U1418 ( .A(\block[4][97] ), .B(\block[5][97] ), .C(\block[6][97] ), 
        .D(\block[7][97] ), .S0(n1030), .S1(n997), .Y(n821) );
  MXI4XL U1419 ( .A(\block[0][1] ), .B(\block[1][1] ), .C(\block[2][1] ), .D(
        \block[3][1] ), .S0(n1043), .S1(n1011), .Y(n920) );
  MXI4XL U1420 ( .A(\block[4][1] ), .B(\block[5][1] ), .C(\block[6][1] ), .D(
        \block[7][1] ), .S0(n1043), .S1(n1011), .Y(n921) );
  CLKMX2X4 U1421 ( .A(n705), .B(n706), .S0(n974), .Y(blockdata[36]) );
  MX4XL U1422 ( .A(\block[0][37] ), .B(\block[1][37] ), .C(\block[2][37] ), 
        .D(\block[3][37] ), .S0(n1038), .S1(n1006), .Y(n707) );
  MX4XL U1423 ( .A(\block[4][37] ), .B(\block[5][37] ), .C(\block[6][37] ), 
        .D(\block[7][37] ), .S0(n1038), .S1(n1006), .Y(n708) );
  MXI2XL U1424 ( .A(n856), .B(n857), .S0(n972), .Y(blockdata[64]) );
  MXI4XL U1425 ( .A(\block[0][64] ), .B(\block[1][64] ), .C(\block[2][64] ), 
        .D(\block[3][64] ), .S0(n1022), .S1(n993), .Y(n856) );
  MXI4XL U1426 ( .A(\block[4][64] ), .B(\block[5][64] ), .C(\block[6][64] ), 
        .D(\block[7][64] ), .S0(n1022), .S1(n993), .Y(n857) );
  MXI2XL U1427 ( .A(n822), .B(n823), .S0(n969), .Y(blockdata[96]) );
  MXI4XL U1428 ( .A(\block[0][96] ), .B(\block[1][96] ), .C(\block[2][96] ), 
        .D(\block[3][96] ), .S0(n1031), .S1(n997), .Y(n822) );
  MXI4XL U1429 ( .A(\block[4][96] ), .B(\block[5][96] ), .C(\block[6][96] ), 
        .D(\block[7][96] ), .S0(n1030), .S1(n997), .Y(n823) );
  MXI2XL U1430 ( .A(n922), .B(n923), .S0(n977), .Y(blockdata[0]) );
  MXI4XL U1431 ( .A(\block[0][0] ), .B(\block[1][0] ), .C(\block[2][0] ), .D(
        \block[3][0] ), .S0(n1043), .S1(n1011), .Y(n922) );
  MXI4XL U1432 ( .A(\block[4][0] ), .B(\block[5][0] ), .C(\block[6][0] ), .D(
        \block[7][0] ), .S0(n1043), .S1(n1011), .Y(n923) );
  MX4X1 U1433 ( .A(\block[0][40] ), .B(\block[1][40] ), .C(\block[2][40] ), 
        .D(\block[3][40] ), .S0(n1037), .S1(n1005), .Y(n713) );
  CLKMX2X2 U1434 ( .A(n715), .B(n716), .S0(n974), .Y(blockdata[41]) );
  CLKMX2X2 U1435 ( .A(n717), .B(n718), .S0(n974), .Y(blockdata[42]) );
  MX4X1 U1436 ( .A(\block[0][72] ), .B(\block[1][72] ), .C(\block[2][72] ), 
        .D(\block[3][72] ), .S0(n1034), .S1(n1001), .Y(n719) );
  MXI2XL U1437 ( .A(n910), .B(n911), .S0(n977), .Y(blockdata[8]) );
  MXI4X1 U1438 ( .A(\block[0][8] ), .B(\block[1][8] ), .C(\block[2][8] ), .D(
        \block[3][8] ), .S0(n1042), .S1(n1010), .Y(n910) );
  MXI4X1 U1439 ( .A(\block[4][8] ), .B(\block[5][8] ), .C(\block[6][8] ), .D(
        \block[7][8] ), .S0(n1042), .S1(n1010), .Y(n911) );
  MX4X1 U1440 ( .A(\block[0][46] ), .B(\block[1][46] ), .C(\block[2][46] ), 
        .D(\block[3][46] ), .S0(n1036), .S1(n1004), .Y(n721) );
  MXI2XL U1441 ( .A(n814), .B(n815), .S0(n969), .Y(blockdata[104]) );
  MXI4X1 U1442 ( .A(\block[0][104] ), .B(\block[1][104] ), .C(\block[2][104] ), 
        .D(\block[3][104] ), .S0(n1029), .S1(n996), .Y(n814) );
  MXI4X1 U1443 ( .A(\block[4][104] ), .B(\block[5][104] ), .C(\block[6][104] ), 
        .D(\block[7][104] ), .S0(n1029), .S1(n996), .Y(n815) );
  CLKMX2X2 U1444 ( .A(n723), .B(n724), .S0(n971), .Y(blockdata[74]) );
  CLKMX2X2 U1445 ( .A(n725), .B(n726), .S0(n968), .Y(blockdata[105]) );
  CLKMX2X2 U1446 ( .A(n727), .B(n728), .S0(n976), .Y(blockdata[12]) );
  CLKMX2X2 U1447 ( .A(n729), .B(n730), .S0(n976), .Y(blockdata[13]) );
  CLKMX2X2 U1448 ( .A(n731), .B(n732), .S0(n971), .Y(blockdata[78]) );
  CLKMX2X2 U1449 ( .A(n733), .B(n734), .S0(n968), .Y(blockdata[108]) );
  CLKMX2X2 U1450 ( .A(n735), .B(n736), .S0(n968), .Y(blockdata[109]) );
  CLKMX2X2 U1451 ( .A(n737), .B(n738), .S0(n976), .Y(blockdata[11]) );
  MXI4X1 U1452 ( .A(\block[4][15] ), .B(\block[5][15] ), .C(\block[6][15] ), 
        .D(\block[7][15] ), .S0(n1041), .S1(n1009), .Y(n909) );
  MXI2XL U1453 ( .A(n862), .B(n863), .S0(n972), .Y(blockdata[57]) );
  MXI4XL U1454 ( .A(\block[4][57] ), .B(\block[5][57] ), .C(\block[6][57] ), 
        .D(\block[7][57] ), .S0(n1032), .S1(n1002), .Y(n863) );
  MXI4XL U1455 ( .A(\block[0][57] ), .B(\block[1][57] ), .C(\block[2][57] ), 
        .D(\block[3][57] ), .S0(n1035), .S1(n1002), .Y(n862) );
  MXI2XL U1456 ( .A(n842), .B(n843), .S0(n970), .Y(blockdata[82]) );
  MXI4X1 U1457 ( .A(\block[4][82] ), .B(\block[5][82] ), .C(\block[6][82] ), 
        .D(\block[7][82] ), .S0(n1033), .S1(n999), .Y(n843) );
  MXI4X1 U1458 ( .A(\block[0][82] ), .B(\block[1][82] ), .C(\block[2][82] ), 
        .D(\block[3][82] ), .S0(n1033), .S1(n999), .Y(n842) );
  MXI2XL U1459 ( .A(n838), .B(n839), .S0(n970), .Y(blockdata[84]) );
  MXI4X1 U1460 ( .A(\block[4][84] ), .B(\block[5][84] ), .C(\block[6][84] ), 
        .D(\block[7][84] ), .S0(n1032), .S1(n999), .Y(n839) );
  MXI4X1 U1461 ( .A(\block[0][84] ), .B(\block[1][84] ), .C(\block[2][84] ), 
        .D(\block[3][84] ), .S0(n1032), .S1(n999), .Y(n838) );
  MXI2XL U1462 ( .A(n834), .B(n835), .S0(n970), .Y(blockdata[86]) );
  MXI4X1 U1463 ( .A(\block[4][86] ), .B(\block[5][86] ), .C(\block[6][86] ), 
        .D(\block[7][86] ), .S0(n1032), .S1(n999), .Y(n835) );
  MXI4X1 U1464 ( .A(\block[0][86] ), .B(\block[1][86] ), .C(\block[2][86] ), 
        .D(\block[3][86] ), .S0(n1032), .S1(n999), .Y(n834) );
  MXI2XL U1465 ( .A(n844), .B(n845), .S0(n970), .Y(blockdata[81]) );
  MXI4X1 U1466 ( .A(\block[4][81] ), .B(\block[5][81] ), .C(\block[6][81] ), 
        .D(\block[7][81] ), .S0(n1033), .S1(n999), .Y(n845) );
  MXI4X1 U1467 ( .A(\block[0][81] ), .B(\block[1][81] ), .C(\block[2][81] ), 
        .D(\block[3][81] ), .S0(n1033), .S1(n999), .Y(n844) );
  MXI2XL U1468 ( .A(n840), .B(n841), .S0(n970), .Y(blockdata[83]) );
  MXI4X1 U1469 ( .A(\block[4][83] ), .B(\block[5][83] ), .C(\block[6][83] ), 
        .D(\block[7][83] ), .S0(n1032), .S1(n999), .Y(n841) );
  MXI4X1 U1470 ( .A(\block[0][83] ), .B(\block[1][83] ), .C(\block[2][83] ), 
        .D(\block[3][83] ), .S0(n1033), .S1(n999), .Y(n840) );
  MXI2XL U1471 ( .A(n836), .B(n837), .S0(n970), .Y(blockdata[85]) );
  MXI4X1 U1472 ( .A(\block[4][85] ), .B(\block[5][85] ), .C(\block[6][85] ), 
        .D(\block[7][85] ), .S0(n1032), .S1(n999), .Y(n837) );
  MXI4X1 U1473 ( .A(\block[0][85] ), .B(\block[1][85] ), .C(\block[2][85] ), 
        .D(\block[3][85] ), .S0(n1032), .S1(n999), .Y(n836) );
  MXI2XL U1474 ( .A(n832), .B(n833), .S0(n970), .Y(blockdata[87]) );
  MXI4XL U1475 ( .A(\block[4][87] ), .B(\block[5][87] ), .C(\block[6][87] ), 
        .D(\block[7][87] ), .S0(n1032), .S1(n998), .Y(n833) );
  MXI4XL U1476 ( .A(\block[0][87] ), .B(\block[1][87] ), .C(\block[2][87] ), 
        .D(\block[3][87] ), .S0(n1032), .S1(n998), .Y(n832) );
  MXI2XL U1477 ( .A(n828), .B(n829), .S0(n970), .Y(blockdata[89]) );
  MXI4XL U1478 ( .A(\block[4][89] ), .B(\block[5][89] ), .C(\block[6][89] ), 
        .D(\block[7][89] ), .S0(n1032), .S1(n998), .Y(n829) );
  MXI4XL U1479 ( .A(\block[0][89] ), .B(\block[1][89] ), .C(\block[2][89] ), 
        .D(\block[3][89] ), .S0(n1032), .S1(n998), .Y(n828) );
  MXI2XL U1480 ( .A(n830), .B(n831), .S0(n970), .Y(blockdata[88]) );
  MXI4XL U1481 ( .A(\block[4][88] ), .B(\block[5][88] ), .C(\block[6][88] ), 
        .D(\block[7][88] ), .S0(n1032), .S1(n998), .Y(n831) );
  MXI4XL U1482 ( .A(\block[0][88] ), .B(\block[1][88] ), .C(\block[2][88] ), 
        .D(\block[3][88] ), .S0(n1032), .S1(n998), .Y(n830) );
  MXI2XL U1483 ( .A(n894), .B(n895), .S0(n975), .Y(blockdata[22]) );
  MXI4XL U1484 ( .A(\block[4][22] ), .B(\block[5][22] ), .C(\block[6][22] ), 
        .D(\block[7][22] ), .S0(n1040), .S1(n1008), .Y(n895) );
  MXI4XL U1485 ( .A(\block[0][22] ), .B(\block[1][22] ), .C(\block[2][22] ), 
        .D(\block[3][22] ), .S0(n1040), .S1(n1008), .Y(n894) );
  MXI2XL U1486 ( .A(n896), .B(n897), .S0(n975), .Y(blockdata[21]) );
  MXI4XL U1487 ( .A(\block[4][21] ), .B(\block[5][21] ), .C(\block[6][21] ), 
        .D(\block[7][21] ), .S0(n1040), .S1(n1008), .Y(n897) );
  MXI4XL U1488 ( .A(\block[0][21] ), .B(\block[1][21] ), .C(\block[2][21] ), 
        .D(\block[3][21] ), .S0(n1040), .S1(n1008), .Y(n896) );
  MXI2XL U1489 ( .A(n892), .B(n893), .S0(n975), .Y(blockdata[23]) );
  MXI4XL U1490 ( .A(\block[4][23] ), .B(\block[5][23] ), .C(\block[6][23] ), 
        .D(\block[7][23] ), .S0(n1040), .S1(n1008), .Y(n893) );
  MXI4XL U1491 ( .A(\block[0][23] ), .B(\block[1][23] ), .C(\block[2][23] ), 
        .D(\block[3][23] ), .S0(n1040), .S1(n1008), .Y(n892) );
  MXI2XL U1492 ( .A(n888), .B(n889), .S0(n975), .Y(blockdata[25]) );
  MXI4XL U1493 ( .A(\block[4][25] ), .B(\block[5][25] ), .C(\block[6][25] ), 
        .D(\block[7][25] ), .S0(n1039), .S1(n1008), .Y(n889) );
  MXI4XL U1494 ( .A(\block[0][25] ), .B(\block[1][25] ), .C(\block[2][25] ), 
        .D(\block[3][25] ), .S0(n1039), .S1(n1008), .Y(n888) );
  MXI2XL U1495 ( .A(n890), .B(n891), .S0(n975), .Y(blockdata[24]) );
  MXI4XL U1496 ( .A(\block[4][24] ), .B(\block[5][24] ), .C(\block[6][24] ), 
        .D(\block[7][24] ), .S0(n1040), .S1(n1008), .Y(n891) );
  MXI4XL U1497 ( .A(\block[0][24] ), .B(\block[1][24] ), .C(\block[2][24] ), 
        .D(\block[3][24] ), .S0(n1040), .S1(n1008), .Y(n890) );
  MXI2X1 U1498 ( .A(n804), .B(n805), .S0(n968), .Y(blockdata[116]) );
  MXI4XL U1499 ( .A(\block[4][116] ), .B(\block[5][116] ), .C(\block[6][116] ), 
        .D(\block[7][116] ), .S0(n1027), .S1(n994), .Y(n805) );
  MXI4XL U1500 ( .A(\block[0][116] ), .B(\block[1][116] ), .C(\block[2][116] ), 
        .D(\block[3][116] ), .S0(n1027), .S1(n994), .Y(n804) );
  AND2XL U1501 ( .A(mem_ready), .B(n1542), .Y(n739) );
  MX2XL U1502 ( .A(n1482), .B(n1481), .S0(n1069), .Y(n1483) );
  INVXL U1503 ( .A(proc_addr[27]), .Y(n1481) );
  MX2XL U1504 ( .A(n1479), .B(n1478), .S0(n1069), .Y(n1480) );
  INVXL U1505 ( .A(proc_addr[28]), .Y(n1478) );
  MX2XL U1506 ( .A(n1519), .B(n1518), .S0(n1068), .Y(n1520) );
  INVXL U1507 ( .A(proc_addr[13]), .Y(n1518) );
  MX2XL U1508 ( .A(n1515), .B(n1514), .S0(n1068), .Y(n1516) );
  INVXL U1509 ( .A(proc_addr[15]), .Y(n1514) );
  MX2XL U1510 ( .A(n1512), .B(n1511), .S0(n1068), .Y(n1513) );
  INVXL U1511 ( .A(proc_addr[16]), .Y(n1511) );
  MX2XL U1512 ( .A(n1509), .B(n1508), .S0(n1068), .Y(n1510) );
  INVXL U1513 ( .A(proc_addr[17]), .Y(n1508) );
  MX2XL U1514 ( .A(n1506), .B(n1505), .S0(n1069), .Y(n1507) );
  INVXL U1515 ( .A(proc_addr[18]), .Y(n1505) );
  MX2XL U1516 ( .A(n1503), .B(n1502), .S0(n1069), .Y(n1504) );
  INVXL U1517 ( .A(proc_addr[19]), .Y(n1502) );
  MX2XL U1518 ( .A(n1500), .B(n215), .S0(n1069), .Y(n1501) );
  MX2XL U1519 ( .A(n210), .B(n221), .S0(n1069), .Y(n1499) );
  MX2XL U1520 ( .A(n1497), .B(n1496), .S0(n1069), .Y(n1498) );
  INVXL U1521 ( .A(proc_addr[22]), .Y(n1496) );
  MX2XL U1522 ( .A(n1491), .B(n1490), .S0(n1069), .Y(n1492) );
  INVXL U1523 ( .A(proc_addr[24]), .Y(n1490) );
  MX2XL U1524 ( .A(n1488), .B(n1487), .S0(n1069), .Y(n1489) );
  INVXL U1525 ( .A(proc_addr[25]), .Y(n1487) );
  MX2XL U1526 ( .A(n1530), .B(n1529), .S0(n1068), .Y(n1531) );
  INVXL U1527 ( .A(proc_addr[7]), .Y(n1529) );
  INVXL U1528 ( .A(tag[2]), .Y(n1530) );
  MX2XL U1529 ( .A(n1525), .B(n1524), .S0(n1068), .Y(n1526) );
  INVXL U1530 ( .A(proc_addr[10]), .Y(n1524) );
  INVXL U1531 ( .A(tag[5]), .Y(n1525) );
  MX2XL U1532 ( .A(n1494), .B(n1493), .S0(n1069), .Y(n1495) );
  INVXL U1533 ( .A(proc_addr[23]), .Y(n1493) );
  INVXL U1534 ( .A(tag[18]), .Y(n1494) );
  MX2XL U1535 ( .A(n1485), .B(n1484), .S0(n1069), .Y(n1486) );
  INVXL U1536 ( .A(proc_addr[26]), .Y(n1484) );
  MX2XL U1537 ( .A(n1533), .B(n1532), .S0(n1068), .Y(n1534) );
  INVXL U1538 ( .A(proc_addr[6]), .Y(n1532) );
  MX2XL U1539 ( .A(n1476), .B(n1475), .S0(n1069), .Y(n1477) );
  INVXL U1540 ( .A(proc_addr[29]), .Y(n1475) );
  MXI2XL U1541 ( .A(n800), .B(n801), .S0(n967), .Y(blockdata[118]) );
  MXI4XL U1542 ( .A(\block[4][118] ), .B(\block[5][118] ), .C(\block[6][118] ), 
        .D(\block[7][118] ), .S0(n1027), .S1(n993), .Y(n801) );
  MXI4XL U1543 ( .A(\block[0][118] ), .B(\block[1][118] ), .C(\block[2][118] ), 
        .D(\block[3][118] ), .S0(n1027), .S1(n993), .Y(n800) );
  MXI2XL U1544 ( .A(n798), .B(n799), .S0(n967), .Y(blockdata[119]) );
  MXI4XL U1545 ( .A(\block[4][119] ), .B(\block[5][119] ), .C(\block[6][119] ), 
        .D(\block[7][119] ), .S0(n1027), .S1(n993), .Y(n799) );
  MXI4XL U1546 ( .A(\block[0][119] ), .B(\block[1][119] ), .C(\block[2][119] ), 
        .D(\block[3][119] ), .S0(n1027), .S1(n993), .Y(n798) );
  MXI2XL U1547 ( .A(n794), .B(n795), .S0(n967), .Y(blockdata[121]) );
  MXI4XL U1548 ( .A(\block[4][121] ), .B(\block[5][121] ), .C(\block[6][121] ), 
        .D(\block[7][121] ), .S0(n1027), .S1(n993), .Y(n795) );
  MXI4XL U1549 ( .A(\block[0][121] ), .B(\block[1][121] ), .C(\block[2][121] ), 
        .D(\block[3][121] ), .S0(n1027), .S1(n993), .Y(n794) );
  MXI2XL U1550 ( .A(n796), .B(n797), .S0(n967), .Y(blockdata[120]) );
  MXI4XL U1551 ( .A(\block[4][120] ), .B(\block[5][120] ), .C(\block[6][120] ), 
        .D(\block[7][120] ), .S0(n1027), .S1(n993), .Y(n797) );
  MXI4XL U1552 ( .A(\block[0][120] ), .B(\block[1][120] ), .C(\block[2][120] ), 
        .D(\block[3][120] ), .S0(n1027), .S1(n993), .Y(n796) );
  MXI2XL U1553 ( .A(n802), .B(n803), .S0(n967), .Y(blockdata[117]) );
  MXI4XL U1554 ( .A(\block[4][117] ), .B(\block[5][117] ), .C(\block[6][117] ), 
        .D(\block[7][117] ), .S0(n1027), .S1(n993), .Y(n803) );
  MXI4XL U1555 ( .A(\block[0][117] ), .B(\block[1][117] ), .C(\block[2][117] ), 
        .D(\block[3][117] ), .S0(n1027), .S1(n993), .Y(n802) );
  MXI2XL U1556 ( .A(n852), .B(n853), .S0(n972), .Y(blockdata[66]) );
  MXI4XL U1557 ( .A(\block[0][66] ), .B(\block[1][66] ), .C(\block[2][66] ), 
        .D(\block[3][66] ), .S0(n1022), .S1(n993), .Y(n852) );
  MXI4XL U1558 ( .A(\block[4][66] ), .B(\block[5][66] ), .C(\block[6][66] ), 
        .D(\block[7][66] ), .S0(n1022), .S1(n993), .Y(n853) );
  MXI2XL U1559 ( .A(n818), .B(n819), .S0(n969), .Y(blockdata[98]) );
  MXI4XL U1560 ( .A(\block[0][98] ), .B(\block[1][98] ), .C(\block[2][98] ), 
        .D(\block[3][98] ), .S0(n1030), .S1(n997), .Y(n818) );
  MXI4XL U1561 ( .A(\block[4][98] ), .B(\block[5][98] ), .C(\block[6][98] ), 
        .D(\block[7][98] ), .S0(n1030), .S1(n997), .Y(n819) );
  MXI4XL U1562 ( .A(\block[0][2] ), .B(\block[1][2] ), .C(\block[2][2] ), .D(
        \block[3][2] ), .S0(n1043), .S1(n1011), .Y(n918) );
  MXI4XL U1563 ( .A(\block[4][2] ), .B(\block[5][2] ), .C(\block[6][2] ), .D(
        \block[7][2] ), .S0(n1043), .S1(n1011), .Y(n919) );
  MXI4XL U1564 ( .A(\block[0][3] ), .B(\block[1][3] ), .C(\block[2][3] ), .D(
        \block[3][3] ), .S0(n1043), .S1(n1010), .Y(n916) );
  MXI4XL U1565 ( .A(\block[4][3] ), .B(\block[5][3] ), .C(\block[6][3] ), .D(
        \block[7][3] ), .S0(n1043), .S1(n1010), .Y(n917) );
  MX4XL U1566 ( .A(\block[0][33] ), .B(\block[1][33] ), .C(\block[2][33] ), 
        .D(\block[3][33] ), .S0(n1038), .S1(n1006), .Y(n740) );
  MX4XL U1567 ( .A(\block[4][33] ), .B(\block[5][33] ), .C(\block[6][33] ), 
        .D(\block[7][33] ), .S0(n1038), .S1(n1006), .Y(n741) );
  MXI2XL U1568 ( .A(n848), .B(n849), .S0(n972), .Y(blockdata[68]) );
  MXI4XL U1569 ( .A(\block[0][68] ), .B(\block[1][68] ), .C(\block[2][68] ), 
        .D(\block[3][68] ), .S0(n1022), .S1(n1001), .Y(n848) );
  MXI4XL U1570 ( .A(\block[4][68] ), .B(\block[5][68] ), .C(\block[6][68] ), 
        .D(\block[7][68] ), .S0(n1022), .S1(n1007), .Y(n849) );
  MX2XL U1571 ( .A(n742), .B(n743), .S0(n969), .Y(blockdata[100]) );
  MXI4XL U1572 ( .A(\block[0][4] ), .B(\block[1][4] ), .C(\block[2][4] ), .D(
        \block[3][4] ), .S0(n1043), .S1(n1010), .Y(n914) );
  MXI4XL U1573 ( .A(\block[4][4] ), .B(\block[5][4] ), .C(\block[6][4] ), .D(
        \block[7][4] ), .S0(n1043), .S1(n1010), .Y(n915) );
  MX2XL U1574 ( .A(n746), .B(n747), .S0(n969), .Y(blockdata[101]) );
  MX4X1 U1575 ( .A(\block[0][101] ), .B(\block[1][101] ), .C(\block[2][101] ), 
        .D(\block[3][101] ), .S0(n1030), .S1(n996), .Y(n746) );
  MX4X1 U1576 ( .A(\block[4][101] ), .B(\block[5][101] ), .C(\block[6][101] ), 
        .D(\block[7][101] ), .S0(n1030), .S1(n996), .Y(n747) );
  MX2XL U1577 ( .A(n750), .B(n751), .S0(n977), .Y(blockdata[5]) );
  MX2XL U1578 ( .A(n754), .B(n755), .S0(n969), .Y(blockdata[103]) );
  MX4X1 U1579 ( .A(\block[0][103] ), .B(\block[1][103] ), .C(\block[2][103] ), 
        .D(\block[3][103] ), .S0(n1029), .S1(n996), .Y(n754) );
  MX4X1 U1580 ( .A(\block[4][103] ), .B(\block[5][103] ), .C(\block[6][103] ), 
        .D(\block[7][103] ), .S0(n1029), .S1(n996), .Y(n755) );
  MX2XL U1581 ( .A(n756), .B(n757), .S0(n977), .Y(blockdata[7]) );
  MX4X1 U1582 ( .A(\block[0][7] ), .B(\block[1][7] ), .C(\block[2][7] ), .D(
        \block[3][7] ), .S0(n1042), .S1(n1010), .Y(n756) );
  MX4X1 U1583 ( .A(\block[4][7] ), .B(\block[5][7] ), .C(\block[6][7] ), .D(
        \block[7][7] ), .S0(n1042), .S1(n1010), .Y(n757) );
  MXI2XL U1584 ( .A(n882), .B(n883), .S0(n975), .Y(blockdata[32]) );
  MXI4XL U1585 ( .A(\block[0][32] ), .B(\block[1][32] ), .C(\block[2][32] ), 
        .D(\block[3][32] ), .S0(n1038), .S1(n1007), .Y(n882) );
  MXI4XL U1586 ( .A(\block[4][32] ), .B(\block[5][32] ), .C(\block[6][32] ), 
        .D(\block[7][32] ), .S0(n1038), .S1(n1007), .Y(n883) );
  MXI2XL U1587 ( .A(n816), .B(n817), .S0(n969), .Y(blockdata[102]) );
  MXI4X1 U1588 ( .A(\block[0][102] ), .B(\block[1][102] ), .C(\block[2][102] ), 
        .D(\block[3][102] ), .S0(n1030), .S1(n996), .Y(n816) );
  MXI4X1 U1589 ( .A(\block[4][102] ), .B(\block[5][102] ), .C(\block[6][102] ), 
        .D(\block[7][102] ), .S0(n1030), .S1(n996), .Y(n817) );
  MXI4X1 U1590 ( .A(\block[0][6] ), .B(\block[1][6] ), .C(\block[2][6] ), .D(
        \block[3][6] ), .S0(n1042), .S1(n1010), .Y(n912) );
  MXI4X1 U1591 ( .A(\block[4][6] ), .B(\block[5][6] ), .C(\block[6][6] ), .D(
        \block[7][6] ), .S0(n1042), .S1(n1010), .Y(n913) );
  CLKMX2X2 U1592 ( .A(n758), .B(n759), .S0(n974), .Y(blockdata[44]) );
  CLKMX2X2 U1593 ( .A(n760), .B(n761), .S0(n971), .Y(blockdata[73]) );
  CLKMX2X2 U1594 ( .A(n762), .B(n763), .S0(n973), .Y(blockdata[45]) );
  CLKMX2X2 U1595 ( .A(n764), .B(n765), .S0(n976), .Y(blockdata[9]) );
  CLKMX2X2 U1596 ( .A(n766), .B(n767), .S0(n974), .Y(blockdata[43]) );
  CLKMX2X2 U1597 ( .A(n768), .B(n769), .S0(n971), .Y(blockdata[76]) );
  CLKMX2X2 U1598 ( .A(n770), .B(n771), .S0(n976), .Y(blockdata[10]) );
  CLKMX2X2 U1599 ( .A(n772), .B(n773), .S0(n971), .Y(blockdata[77]) );
  CLKMX2X2 U1600 ( .A(n774), .B(n775), .S0(n973), .Y(blockdata[47]) );
  CLKMX2X2 U1601 ( .A(n776), .B(n777), .S0(n968), .Y(blockdata[106]) );
  CLKMX2X2 U1602 ( .A(n778), .B(n779), .S0(n971), .Y(blockdata[75]) );
  CLKMX2X2 U1603 ( .A(n782), .B(n783), .S0(n971), .Y(blockdata[79]) );
  CLKMX2X2 U1604 ( .A(n784), .B(n785), .S0(n968), .Y(blockdata[110]) );
  CLKMX2X2 U1605 ( .A(n786), .B(n787), .S0(n968), .Y(blockdata[107]) );
  MX4X1 U1606 ( .A(\block[0][111] ), .B(\block[1][111] ), .C(\block[2][111] ), 
        .D(\block[3][111] ), .S0(n1028), .S1(n994), .Y(n788) );
  MX4X1 U1607 ( .A(\block[4][111] ), .B(\block[5][111] ), .C(\block[6][111] ), 
        .D(\block[7][111] ), .S0(n1028), .S1(n994), .Y(n789) );
  MXI2X1 U1608 ( .A(n1739), .B(n1537), .S0(n570), .Y(n1723) );
  MXI2X1 U1609 ( .A(n1738), .B(n1537), .S0(n564), .Y(n1722) );
  MXI2X1 U1610 ( .A(n1737), .B(n1537), .S0(n572), .Y(n1721) );
  MXI2X1 U1611 ( .A(n1736), .B(n1537), .S0(n566), .Y(n1720) );
  MXI2XL U1612 ( .A(n1747), .B(n1538), .S0(n570), .Y(n1731) );
  MXI2XL U1613 ( .A(n1746), .B(n1538), .S0(n564), .Y(n1730) );
  MXI2XL U1614 ( .A(n1745), .B(n1538), .S0(n572), .Y(n1729) );
  MXI2XL U1615 ( .A(n1744), .B(n1538), .S0(n566), .Y(n1728) );
  MXI2XL U1616 ( .A(n1743), .B(n1538), .S0(n573), .Y(n1727) );
  MXI2XL U1617 ( .A(n1742), .B(n1538), .S0(n567), .Y(n1726) );
  MXI2XL U1618 ( .A(n1741), .B(n1538), .S0(n571), .Y(n1725) );
  MXI2XL U1619 ( .A(n1740), .B(n1538), .S0(n565), .Y(n1724) );
  AO21XL U1620 ( .A0(mem_ready), .A1(n1540), .B0(valid), .Y(n1471) );
  NAND3BXL U1621 ( .AN(n1303), .B(proc_write), .C(n1049), .Y(n1473) );
  CLKINVX1 U1622 ( .A(proc_wdata[0]), .Y(n1469) );
  CLKINVX1 U1623 ( .A(proc_wdata[1]), .Y(n1467) );
  CLKINVX1 U1624 ( .A(proc_wdata[2]), .Y(n1465) );
  CLKINVX1 U1625 ( .A(proc_wdata[3]), .Y(n1463) );
  CLKINVX1 U1626 ( .A(proc_wdata[4]), .Y(n1461) );
  CLKINVX1 U1627 ( .A(proc_wdata[5]), .Y(n1459) );
  CLKINVX1 U1628 ( .A(proc_wdata[6]), .Y(n1457) );
  CLKINVX1 U1629 ( .A(proc_wdata[7]), .Y(n1455) );
  CLKINVX1 U1630 ( .A(proc_wdata[8]), .Y(n1453) );
  CLKINVX1 U1631 ( .A(proc_wdata[9]), .Y(n1451) );
  CLKINVX1 U1632 ( .A(proc_wdata[10]), .Y(n1449) );
  CLKINVX1 U1633 ( .A(proc_wdata[11]), .Y(n1447) );
  CLKINVX1 U1634 ( .A(proc_wdata[12]), .Y(n1445) );
  CLKINVX1 U1635 ( .A(proc_wdata[13]), .Y(n1443) );
  CLKINVX1 U1636 ( .A(proc_wdata[14]), .Y(n1441) );
  CLKINVX1 U1637 ( .A(proc_wdata[15]), .Y(n1439) );
  CLKINVX1 U1638 ( .A(proc_wdata[16]), .Y(n1437) );
  CLKINVX1 U1639 ( .A(proc_wdata[17]), .Y(n1435) );
  CLKINVX1 U1640 ( .A(proc_wdata[18]), .Y(n1433) );
  CLKINVX1 U1641 ( .A(proc_wdata[19]), .Y(n1431) );
  CLKINVX1 U1642 ( .A(proc_wdata[20]), .Y(n1429) );
  CLKINVX1 U1643 ( .A(proc_wdata[21]), .Y(n1427) );
  CLKINVX1 U1644 ( .A(proc_wdata[22]), .Y(n1425) );
  CLKINVX1 U1645 ( .A(proc_wdata[23]), .Y(n1423) );
  CLKINVX1 U1646 ( .A(proc_wdata[24]), .Y(n1421) );
  CLKINVX1 U1647 ( .A(proc_wdata[25]), .Y(n1419) );
  CLKINVX1 U1648 ( .A(proc_wdata[26]), .Y(n1417) );
  CLKINVX1 U1649 ( .A(proc_wdata[27]), .Y(n1415) );
  CLKINVX1 U1650 ( .A(proc_wdata[28]), .Y(n1413) );
  CLKINVX1 U1651 ( .A(proc_wdata[29]), .Y(n1411) );
  CLKINVX1 U1652 ( .A(proc_wdata[30]), .Y(n1409) );
  CLKINVX1 U1653 ( .A(proc_wdata[31]), .Y(n1407) );
  CLKINVX1 U1654 ( .A(proc_write), .Y(n1546) );
  MXI2X4 U1655 ( .A(n790), .B(n791), .S0(n967), .Y(blockdata[127]) );
  MXI2X4 U1656 ( .A(n792), .B(n793), .S0(n967), .Y(blockdata[124]) );
  MXI2X4 U1657 ( .A(n824), .B(n825), .S0(n969), .Y(blockdata[95]) );
  MXI2X4 U1658 ( .A(n826), .B(n827), .S0(n970), .Y(blockdata[92]) );
  MXI2X4 U1659 ( .A(n858), .B(n859), .S0(n972), .Y(blockdata[63]) );
  MXI2X4 U1660 ( .A(n860), .B(n861), .S0(n972), .Y(blockdata[60]) );
  MXI2X4 U1661 ( .A(n884), .B(n885), .S0(n975), .Y(blockdata[31]) );
  MXI2X4 U1662 ( .A(n886), .B(n887), .S0(n975), .Y(blockdata[28]) );
  MXI2X4 U1663 ( .A(n924), .B(n925), .S0(n977), .Y(valid) );
  MXI2X4 U1664 ( .A(n928), .B(n929), .S0(n978), .Y(tag[22]) );
  MXI2X4 U1665 ( .A(n932), .B(n933), .S0(n978), .Y(tag[18]) );
  MXI2X4 U1666 ( .A(n934), .B(n935), .S0(n978), .Y(tag[17]) );
  MXI2X4 U1667 ( .A(n938), .B(n939), .S0(n978), .Y(tag[15]) );
  MXI2X4 U1668 ( .A(n940), .B(n941), .S0(n978), .Y(tag[14]) );
  MXI2X4 U1669 ( .A(n942), .B(n943), .S0(n978), .Y(tag[13]) );
  MXI2X4 U1670 ( .A(n944), .B(n945), .S0(n978), .Y(tag[12]) );
  MXI2X4 U1671 ( .A(n946), .B(n947), .S0(n979), .Y(tag[11]) );
  MXI2X4 U1672 ( .A(n948), .B(n949), .S0(n979), .Y(tag[10]) );
  MXI2X4 U1673 ( .A(n950), .B(n951), .S0(n979), .Y(tag[8]) );
  MXI2X4 U1674 ( .A(n952), .B(n953), .S0(n979), .Y(tag[7]) );
  MXI2X4 U1675 ( .A(n954), .B(n955), .S0(n979), .Y(tag[5]) );
  MXI2X4 U1676 ( .A(n956), .B(n957), .S0(n979), .Y(tag[3]) );
  MXI2X4 U1677 ( .A(n960), .B(n961), .S0(n979), .Y(tag[1]) );
  MXI4X4 U1678 ( .A(\blocktag[4][17] ), .B(\blocktag[5][17] ), .C(
        \blocktag[6][17] ), .D(\blocktag[7][17] ), .S0(n1045), .S1(n980), .Y(
        n935) );
  MXI4X4 U1679 ( .A(\blocktag[0][17] ), .B(\blocktag[1][17] ), .C(
        \blocktag[2][17] ), .D(\blocktag[3][17] ), .S0(n1045), .S1(n985), .Y(
        n934) );
  MXI4X4 U1680 ( .A(\blocktag[4][14] ), .B(\blocktag[5][14] ), .C(
        \blocktag[6][14] ), .D(\blocktag[7][14] ), .S0(n1045), .S1(n980), .Y(
        n941) );
  MXI4X4 U1681 ( .A(\blocktag[0][14] ), .B(\blocktag[1][14] ), .C(
        \blocktag[2][14] ), .D(\blocktag[3][14] ), .S0(n1045), .S1(n983), .Y(
        n940) );
  MXI4X4 U1682 ( .A(\blocktag[4][13] ), .B(\blocktag[5][13] ), .C(
        \blocktag[6][13] ), .D(\blocktag[7][13] ), .S0(n1045), .S1(n982), .Y(
        n943) );
  MXI4X4 U1683 ( .A(\blocktag[0][13] ), .B(\blocktag[1][13] ), .C(
        \blocktag[2][13] ), .D(\blocktag[3][13] ), .S0(n1045), .S1(n1011), .Y(
        n942) );
  MXI4X4 U1684 ( .A(\blocktag[4][11] ), .B(\blocktag[5][11] ), .C(
        \blocktag[6][11] ), .D(\blocktag[7][11] ), .S0(n1046), .S1(n1012), .Y(
        n947) );
  MXI4X4 U1685 ( .A(\blocktag[0][11] ), .B(\blocktag[1][11] ), .C(
        \blocktag[2][11] ), .D(\blocktag[3][11] ), .S0(n1046), .S1(n1012), .Y(
        n946) );
  MXI4X4 U1686 ( .A(\blocktag[4][10] ), .B(\blocktag[5][10] ), .C(
        \blocktag[6][10] ), .D(\blocktag[7][10] ), .S0(n1046), .S1(n1012), .Y(
        n949) );
  MXI4X4 U1687 ( .A(\blocktag[0][10] ), .B(\blocktag[1][10] ), .C(
        \blocktag[2][10] ), .D(\blocktag[3][10] ), .S0(n1046), .S1(n1012), .Y(
        n948) );
  XNOR2X4 U1688 ( .A(proc_addr[8]), .B(tag[3]), .Y(n1263) );
  XNOR2X4 U1689 ( .A(proc_addr[10]), .B(tag[5]), .Y(n1262) );
  CLKINVX3 U1690 ( .A(tag[12]), .Y(n1509) );
  XOR2X4 U1691 ( .A(n1509), .B(proc_addr[17]), .Y(n1272) );
  CLKINVX3 U1692 ( .A(tag[14]), .Y(n1503) );
  XOR2X4 U1693 ( .A(n1503), .B(proc_addr[19]), .Y(n1271) );
  CLKINVX3 U1694 ( .A(tag[11]), .Y(n1512) );
  XOR2X4 U1695 ( .A(n1512), .B(proc_addr[16]), .Y(n1269) );
  CLKINVX3 U1696 ( .A(tag[8]), .Y(n1519) );
  XOR2X4 U1697 ( .A(n1519), .B(proc_addr[13]), .Y(n1273) );
  NAND2X4 U1698 ( .A(n1274), .B(n1273), .Y(n1275) );
  CLKINVX3 U1699 ( .A(tag[17]), .Y(n1497) );
  XOR2X4 U1700 ( .A(n1497), .B(proc_addr[22]), .Y(n1280) );
  CLKINVX3 U1701 ( .A(tag[10]), .Y(n1515) );
  XOR2X4 U1702 ( .A(n1533), .B(proc_addr[6]), .Y(n1277) );
  CLKINVX3 U1703 ( .A(tag[13]), .Y(n1506) );
  XOR2X4 U1704 ( .A(n1506), .B(proc_addr[18]), .Y(n1281) );
  XOR2X4 U1705 ( .A(n1488), .B(proc_addr[25]), .Y(n1290) );
  NAND2X4 U1706 ( .A(n1290), .B(n1289), .Y(n1291) );
  NAND2X2 U1707 ( .A(n1049), .B(n1546), .Y(n1540) );
  CLKINVX3 U1708 ( .A(n1301), .Y(n1337) );
  CLKINVX3 U1709 ( .A(blockdata[127]), .Y(n1712) );
  CLKINVX3 U1710 ( .A(blockdata[124]), .Y(n1695) );
  OAI221X2 U1711 ( .A0(n1050), .A1(n1660), .B0(n1427), .B1(n1052), .C0(n1314), 
        .Y(block_next[117]) );
  OAI221X2 U1712 ( .A0(n1050), .A1(n1655), .B0(n1429), .B1(n1052), .C0(n1315), 
        .Y(block_next[116]) );
  OAI221X2 U1713 ( .A0(n1051), .A1(n1650), .B0(n1431), .B1(n1053), .C0(n1316), 
        .Y(block_next[115]) );
  OAI221X2 U1714 ( .A0(n1051), .A1(n1645), .B0(n1433), .B1(n1053), .C0(n1317), 
        .Y(block_next[114]) );
  OAI221X2 U1715 ( .A0(n1051), .A1(n1640), .B0(n1435), .B1(n1053), .C0(n1318), 
        .Y(block_next[113]) );
  OAI221X2 U1716 ( .A0(n1051), .A1(n1635), .B0(n1437), .B1(n1053), .C0(n1319), 
        .Y(block_next[112]) );
  OAI221X2 U1717 ( .A0(n1051), .A1(n1630), .B0(n1439), .B1(n1053), .C0(n1320), 
        .Y(block_next[111]) );
  OAI221X2 U1718 ( .A0(n1051), .A1(n1625), .B0(n1441), .B1(n1053), .C0(n1321), 
        .Y(block_next[110]) );
  OAI221X2 U1719 ( .A0(n1051), .A1(n1620), .B0(n1443), .B1(n1053), .C0(n1322), 
        .Y(block_next[109]) );
  OAI221X2 U1720 ( .A0(n1051), .A1(n1615), .B0(n1445), .B1(n1053), .C0(n1323), 
        .Y(block_next[108]) );
  OAI221X2 U1721 ( .A0(n1051), .A1(n1610), .B0(n1447), .B1(n1053), .C0(n1324), 
        .Y(block_next[107]) );
  OAI221X2 U1722 ( .A0(n1051), .A1(n1605), .B0(n1449), .B1(n1053), .C0(n1325), 
        .Y(block_next[106]) );
  OAI221X2 U1723 ( .A0(n1051), .A1(n1600), .B0(n1451), .B1(n1053), .C0(n1326), 
        .Y(block_next[105]) );
  OAI221X2 U1724 ( .A0(n1050), .A1(n1585), .B0(n1457), .B1(n1053), .C0(n1329), 
        .Y(block_next[102]) );
  OAI221X2 U1725 ( .A0(n1051), .A1(n1575), .B0(n1461), .B1(n1052), .C0(n1331), 
        .Y(block_next[100]) );
  OAI221X2 U1726 ( .A0(n1050), .A1(n1570), .B0(n1463), .B1(n1053), .C0(n1332), 
        .Y(block_next[99]) );
  OAI221X2 U1727 ( .A0(n1050), .A1(n1565), .B0(n1465), .B1(n1052), .C0(n1333), 
        .Y(block_next[98]) );
  OAI221X2 U1728 ( .A0(n1050), .A1(n1560), .B0(n1467), .B1(n1052), .C0(n1334), 
        .Y(block_next[97]) );
  OAI221X2 U1729 ( .A0(n1050), .A1(n1555), .B0(n1469), .B1(n1052), .C0(n1335), 
        .Y(block_next[96]) );
  CLKINVX3 U1730 ( .A(n1338), .Y(n1371) );
  CLKINVX3 U1731 ( .A(blockdata[95]), .Y(n1709) );
  OAI221X2 U1732 ( .A0(n1054), .A1(n1709), .B0(n1407), .B1(n1057), .C0(n1339), 
        .Y(block_next[95]) );
  OAI221X2 U1733 ( .A0(n1054), .A1(n1703), .B0(n1409), .B1(n1057), .C0(n1340), 
        .Y(block_next[94]) );
  OAI221X2 U1734 ( .A0(n1054), .A1(n1698), .B0(n1411), .B1(n1057), .C0(n1341), 
        .Y(block_next[93]) );
  CLKINVX3 U1735 ( .A(blockdata[92]), .Y(n1693) );
  OAI221X2 U1736 ( .A0(n1054), .A1(n1693), .B0(n1413), .B1(n1057), .C0(n1342), 
        .Y(block_next[92]) );
  OAI221X2 U1737 ( .A0(n1054), .A1(n1553), .B0(n1469), .B1(n1056), .C0(n1370), 
        .Y(block_next[64]) );
  CLKINVX3 U1738 ( .A(blockdata[63]), .Y(n1707) );
  OAI221X2 U1739 ( .A0(n1058), .A1(n1707), .B0(n1407), .B1(n1060), .C0(n1373), 
        .Y(block_next[63]) );
  CLKINVX3 U1740 ( .A(blockdata[60]), .Y(n1692) );
  OAI221X2 U1741 ( .A0(n1058), .A1(n1692), .B0(n1413), .B1(n1060), .C0(n1376), 
        .Y(block_next[60]) );
  OAI221X2 U1742 ( .A0(n1058), .A1(n1587), .B0(n1455), .B1(n1061), .C0(n1397), 
        .Y(block_next[39]) );
  OAI221X2 U1743 ( .A0(n1059), .A1(n1582), .B0(n1457), .B1(n1060), .C0(n1398), 
        .Y(block_next[38]) );
  OAI221X2 U1744 ( .A0(n1058), .A1(n1577), .B0(n1459), .B1(n1060), .C0(n1399), 
        .Y(block_next[37]) );
  OAI221X2 U1745 ( .A0(n1059), .A1(n1572), .B0(n1461), .B1(n1060), .C0(n1400), 
        .Y(block_next[36]) );
  OAI221X2 U1746 ( .A0(n1058), .A1(n1567), .B0(n1463), .B1(n1060), .C0(n1401), 
        .Y(block_next[35]) );
  OAI221X2 U1747 ( .A0(n1059), .A1(n1557), .B0(n1467), .B1(n1060), .C0(n1403), 
        .Y(block_next[33]) );
  OAI221X2 U1748 ( .A0(n1059), .A1(n1552), .B0(n1469), .B1(n1060), .C0(n1404), 
        .Y(block_next[32]) );
  CLKINVX3 U1749 ( .A(blockdata[31]), .Y(n1714) );
  OAI221X2 U1750 ( .A0(n1065), .A1(n1407), .B0(n1063), .B1(n1714), .C0(n1406), 
        .Y(block_next[31]) );
  OAI221X2 U1751 ( .A0(n1065), .A1(n1409), .B0(n1063), .B1(n1706), .C0(n1408), 
        .Y(block_next[30]) );
  OAI221X2 U1752 ( .A0(n1065), .A1(n1411), .B0(n1063), .B1(n1701), .C0(n1410), 
        .Y(block_next[29]) );
  CLKINVX3 U1753 ( .A(blockdata[28]), .Y(n1696) );
  OAI221X2 U1754 ( .A0(n1065), .A1(n1413), .B0(n1063), .B1(n1696), .C0(n1412), 
        .Y(block_next[28]) );
  OAI221X2 U1755 ( .A0(n1065), .A1(n1415), .B0(n1063), .B1(n1691), .C0(n1414), 
        .Y(block_next[27]) );
  OAI221X2 U1756 ( .A0(n1066), .A1(n1469), .B0(n1064), .B1(n1556), .C0(n1468), 
        .Y(block_next[0]) );
  CLKINVX3 U1757 ( .A(n1471), .Y(n1537) );
  CLKINVX3 U1758 ( .A(mem_ready), .Y(n1539) );
  CLKINVX3 U1759 ( .A(n1477), .Y(blocktag_next[24]) );
  CLKINVX3 U1760 ( .A(n1480), .Y(blocktag_next[23]) );
  CLKINVX3 U1761 ( .A(n1483), .Y(blocktag_next[22]) );
  CLKINVX3 U1762 ( .A(n1486), .Y(blocktag_next[21]) );
  CLKINVX3 U1763 ( .A(n1489), .Y(blocktag_next[20]) );
  CLKINVX3 U1764 ( .A(n1492), .Y(blocktag_next[19]) );
  CLKINVX3 U1765 ( .A(n1495), .Y(blocktag_next[18]) );
  CLKINVX3 U1766 ( .A(n1498), .Y(blocktag_next[17]) );
  CLKINVX3 U1767 ( .A(n1499), .Y(blocktag_next[16]) );
  CLKINVX3 U1768 ( .A(n1501), .Y(blocktag_next[15]) );
  CLKINVX3 U1769 ( .A(n1504), .Y(blocktag_next[14]) );
  CLKINVX3 U1770 ( .A(n1507), .Y(blocktag_next[13]) );
  CLKINVX3 U1771 ( .A(n1510), .Y(blocktag_next[12]) );
  CLKINVX3 U1772 ( .A(n1513), .Y(blocktag_next[11]) );
  CLKINVX3 U1773 ( .A(n1516), .Y(blocktag_next[10]) );
  CLKINVX3 U1774 ( .A(n1517), .Y(blocktag_next[9]) );
  CLKINVX3 U1775 ( .A(n1520), .Y(blocktag_next[8]) );
  CLKINVX3 U1776 ( .A(n1523), .Y(blocktag_next[6]) );
  CLKINVX3 U1777 ( .A(n1526), .Y(blocktag_next[5]) );
  CLKINVX3 U1778 ( .A(n1527), .Y(blocktag_next[4]) );
  CLKINVX3 U1779 ( .A(n1531), .Y(blocktag_next[2]) );
  CLKINVX3 U1780 ( .A(n1534), .Y(blocktag_next[1]) );
  CLKAND2X4 U1781 ( .A(n1256), .B(blockdata[5]), .Y(n1851) );
  CLKAND2X4 U1782 ( .A(n1255), .B(blockdata[7]), .Y(n1850) );
  CLKAND2X4 U1783 ( .A(n1255), .B(blockdata[9]), .Y(n1848) );
  CLKAND2X4 U1784 ( .A(n1255), .B(blockdata[10]), .Y(n1847) );
  CLKAND2X4 U1785 ( .A(n1255), .B(blockdata[11]), .Y(n1846) );
  CLKAND2X4 U1786 ( .A(n1255), .B(blockdata[12]), .Y(n1845) );
  CLKAND2X4 U1787 ( .A(n1255), .B(blockdata[13]), .Y(n1844) );
  CLKAND2X4 U1788 ( .A(n1255), .B(blockdata[15]), .Y(n1843) );
  CLKAND2X4 U1789 ( .A(n1255), .B(blockdata[26]), .Y(n1832) );
  CLKAND2X4 U1790 ( .A(n1255), .B(blockdata[27]), .Y(n1831) );
  CLKAND2X4 U1791 ( .A(n1255), .B(blockdata[29]), .Y(n1830) );
  CLKAND2X4 U1792 ( .A(n1255), .B(blockdata[30]), .Y(n1829) );
  CLKAND2X4 U1793 ( .A(n1255), .B(blockdata[33]), .Y(n1827) );
  CLKAND2X4 U1794 ( .A(n1255), .B(blockdata[34]), .Y(n1826) );
  CLKAND2X4 U1795 ( .A(n1255), .B(blockdata[35]), .Y(n1825) );
  CLKAND2X4 U1796 ( .A(n1255), .B(blockdata[36]), .Y(n1824) );
  CLKAND2X4 U1797 ( .A(n1254), .B(blockdata[37]), .Y(n1823) );
  CLKAND2X4 U1798 ( .A(n1255), .B(blockdata[38]), .Y(n1822) );
  CLKAND2X4 U1799 ( .A(n1255), .B(blockdata[39]), .Y(n1821) );
  CLKAND2X4 U1800 ( .A(n1255), .B(blockdata[40]), .Y(n1820) );
  CLKAND2X4 U1801 ( .A(n1255), .B(blockdata[41]), .Y(n1819) );
  CLKAND2X4 U1802 ( .A(n1255), .B(blockdata[42]), .Y(n1818) );
  CLKAND2X4 U1803 ( .A(n1255), .B(blockdata[43]), .Y(n1817) );
  CLKAND2X4 U1804 ( .A(n1255), .B(blockdata[44]), .Y(n1816) );
  CLKAND2X4 U1805 ( .A(n1255), .B(blockdata[45]), .Y(n1815) );
  CLKAND2X4 U1806 ( .A(n1254), .B(blockdata[47]), .Y(n1814) );
  CLKAND2X4 U1807 ( .A(n1254), .B(blockdata[58]), .Y(n1803) );
  CLKAND2X4 U1808 ( .A(n1254), .B(blockdata[59]), .Y(n1802) );
  CLKAND2X4 U1809 ( .A(n1254), .B(blockdata[61]), .Y(n1801) );
  CLKAND2X4 U1810 ( .A(n1254), .B(blockdata[62]), .Y(n1800) );
  CLKAND2X4 U1811 ( .A(n1254), .B(blockdata[69]), .Y(n1794) );
  CLKAND2X4 U1812 ( .A(n1254), .B(blockdata[70]), .Y(n1793) );
  CLKAND2X4 U1813 ( .A(n1254), .B(blockdata[71]), .Y(n1792) );
  CLKAND2X4 U1814 ( .A(n1254), .B(blockdata[72]), .Y(n1791) );
  CLKAND2X4 U1815 ( .A(n1254), .B(blockdata[73]), .Y(n1790) );
  CLKAND2X4 U1816 ( .A(n1254), .B(blockdata[74]), .Y(n1789) );
  CLKAND2X4 U1817 ( .A(n1254), .B(blockdata[75]), .Y(n1788) );
  CLKAND2X4 U1818 ( .A(n1254), .B(blockdata[76]), .Y(n1787) );
  CLKAND2X4 U1819 ( .A(n1254), .B(blockdata[77]), .Y(n1786) );
  CLKAND2X4 U1820 ( .A(n1254), .B(blockdata[78]), .Y(n1785) );
  CLKAND2X4 U1821 ( .A(n1254), .B(blockdata[79]), .Y(n1784) );
  CLKAND2X4 U1822 ( .A(n1544), .B(n1248), .Y(n1779) );
  NAND2X2 U1823 ( .A(n692), .B(n1548), .Y(n1713) );
  OAI221X2 U1824 ( .A0(n1094), .A1(n1566), .B0(n1091), .B1(n1565), .C0(n1564), 
        .Y(proc_rdata[2]) );
  OAI221X2 U1825 ( .A0(n1094), .A1(n1591), .B0(n1091), .B1(n1590), .C0(n1589), 
        .Y(proc_rdata[7]) );
  OA22X4 U1826 ( .A0(n1089), .A1(n1693), .B0(n1085), .B1(n1692), .Y(n1694) );
  OAI221X2 U1827 ( .A0(n1096), .A1(n1696), .B0(n1092), .B1(n1695), .C0(n1694), 
        .Y(proc_rdata[28]) );
  OA22X4 U1828 ( .A0(n1089), .A1(n1709), .B0(n1085), .B1(n1707), .Y(n1711) );
  OAI221X2 U1829 ( .A0(n1096), .A1(n1714), .B0(n1092), .B1(n1712), .C0(n1711), 
        .Y(proc_rdata[31]) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, ICACHE_ren, ICACHE_stall, DCACHE_ren, DCACHE_stall,
         n2, n4, n11, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31, n33,
         n35, n37, n39, n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61,
         n63, n65, n67, n69, n71, n73, n75, n77, n81, n83, n85, n87, n89, n91,
         n93, n95, n97, n99, n101, n103, n105, n107, n109, n111, n113, n115,
         n117, n119, n121, n123, n125, n127, n129, n131, n133, n135, n137,
         n139, n141, n143, n145, n147, n149, n151, n154, n156, n158, n160,
         n162, n164, n166, n168, n170, n172, n174, n176, n178, n180, n182,
         n184, n186, n188, n190, n192, n194, n196, n198, n200, n202, n204,
         n206, n208, n210, n212, n214, n216, n218, n220, n222, n224, n228,
         n232, n236, n240, n244, n248, n252, n254, n256, n258, n260, n262,
         n277, n279, n281, n283, n285, n287, n289, n295, n296, n297, n299,
         n301, n302;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .clk(clk), .rst_n(n301), .ICACHE_ren(ICACHE_ren), 
        .ICACHE_addr(ICACHE_addr), .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(
        ICACHE_rdata), .DCACHE_ren(DCACHE_ren), .DCACHE_wen(DCACHE_wen), 
        .DCACHE_addr({DCACHE_addr[29:5], n468, n469, n470, DCACHE_addr[1:0]}), 
        .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(DCACHE_stall), 
        .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n302), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr({DCACHE_addr[29:4], n299, 
        DCACHE_addr[2:0]}), .proc_wdata(DCACHE_wdata), .proc_stall(
        DCACHE_stall), .proc_rdata(DCACHE_rdata), .mem_read(n303), .mem_write(
        n304), .mem_addr({mem_addr_D[31:18], n305, n306, mem_addr_D[15], n307, 
        mem_addr_D[13], n308, n309, mem_addr_D[10], n310, n311, mem_addr_D[7], 
        n312, n313, n314}), .mem_rdata(mem_rdata_D), .mem_wdata({
        mem_wdata_D[127:121], n315, n316, n317, n318, n319, n320, n321, n322, 
        n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
        n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
        n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
        n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
        n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
        n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
        n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
        n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
        mem_wdata_D[6:0]}), .mem_ready(mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n302), .proc_read(ICACHE_ren), 
        .proc_write(1'b0), .proc_addr({ICACHE_addr[29:5], n297, n296, n295, 
        ICACHE_addr[1:0]}), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(ICACHE_rdata), 
        .mem_read(n429), .mem_write(n430), .mem_addr({mem_addr_I[31:5], n431}), 
        .mem_rdata(mem_rdata_I), .mem_wdata({mem_wdata_I[127], n432, n433, 
        mem_wdata_I[124:122], n434, n435, n436, n437, n438, n439, n440, n441, 
        n442, n443, mem_wdata_I[111], n444, n445, n446, n447, n448, n449, n450, 
        n451, n452, n453, n454, n455, n456, n457, n458, mem_wdata_I[95], n459, 
        mem_wdata_I[93:90], n460, n461, n462, n463, n464, n465, n466, 
        mem_wdata_I[82:1], n467}), .mem_ready(mem_ready_I) );
  INVX3 U2 ( .A(n461), .Y(n11) );
  INVX3 U3 ( .A(n460), .Y(n13) );
  INVX3 U4 ( .A(n459), .Y(n15) );
  INVX3 U5 ( .A(n458), .Y(n17) );
  INVX3 U6 ( .A(n457), .Y(n19) );
  INVX3 U7 ( .A(n456), .Y(n21) );
  INVX3 U8 ( .A(n455), .Y(n23) );
  INVX3 U9 ( .A(n454), .Y(n25) );
  INVX3 U10 ( .A(n453), .Y(n27) );
  INVX3 U11 ( .A(n452), .Y(n29) );
  INVX3 U12 ( .A(n451), .Y(n31) );
  INVX3 U13 ( .A(n450), .Y(n33) );
  INVX3 U14 ( .A(n449), .Y(n35) );
  INVX3 U15 ( .A(n448), .Y(n39) );
  INVX3 U16 ( .A(n447), .Y(n41) );
  INVX3 U17 ( .A(n446), .Y(n43) );
  INVX3 U18 ( .A(n445), .Y(n45) );
  INVX3 U19 ( .A(n444), .Y(n47) );
  INVX3 U20 ( .A(n443), .Y(n49) );
  INVX3 U21 ( .A(n442), .Y(n51) );
  INVX3 U22 ( .A(n441), .Y(n53) );
  INVX3 U23 ( .A(n440), .Y(n55) );
  INVX3 U24 ( .A(n439), .Y(n57) );
  INVX3 U25 ( .A(n438), .Y(n59) );
  INVX3 U26 ( .A(n437), .Y(n61) );
  INVX3 U27 ( .A(n436), .Y(n63) );
  INVX3 U28 ( .A(n435), .Y(n65) );
  BUFX20 U29 ( .A(n428), .Y(mem_wdata_D[7]) );
  CLKBUFX12 U30 ( .A(n352), .Y(mem_wdata_D[83]) );
  INVX3 U31 ( .A(n351), .Y(n158) );
  INVX3 U32 ( .A(n350), .Y(n164) );
  INVX3 U33 ( .A(n349), .Y(n170) );
  INVX3 U34 ( .A(n348), .Y(n176) );
  INVX3 U35 ( .A(n347), .Y(n182) );
  INVX3 U36 ( .A(n346), .Y(n188) );
  INVX3 U37 ( .A(n345), .Y(n194) );
  INVX3 U38 ( .A(n344), .Y(n200) );
  INVX3 U39 ( .A(n343), .Y(n206) );
  INVX3 U40 ( .A(n342), .Y(n212) );
  INVX3 U41 ( .A(n341), .Y(n218) );
  INVX3 U42 ( .A(n340), .Y(n224) );
  INVX3 U43 ( .A(n339), .Y(n228) );
  INVX3 U44 ( .A(n338), .Y(n232) );
  INVX3 U45 ( .A(n337), .Y(n236) );
  INVX3 U46 ( .A(n336), .Y(n240) );
  INVX3 U47 ( .A(n335), .Y(n244) );
  INVX3 U48 ( .A(n334), .Y(n248) );
  INVX3 U49 ( .A(n333), .Y(n252) );
  INVX3 U50 ( .A(n332), .Y(n254) );
  INVX3 U51 ( .A(n331), .Y(n256) );
  INVX3 U52 ( .A(n330), .Y(n258) );
  INVX3 U53 ( .A(n329), .Y(n260) );
  INVX3 U54 ( .A(n328), .Y(n262) );
  CLKBUFX12 U55 ( .A(n327), .Y(mem_wdata_D[108]) );
  CLKBUFX12 U56 ( .A(n326), .Y(mem_wdata_D[109]) );
  CLKBUFX12 U57 ( .A(n325), .Y(mem_wdata_D[110]) );
  CLKBUFX12 U58 ( .A(n324), .Y(mem_wdata_D[111]) );
  CLKBUFX12 U59 ( .A(n323), .Y(mem_wdata_D[112]) );
  CLKBUFX12 U60 ( .A(n322), .Y(mem_wdata_D[113]) );
  CLKBUFX12 U61 ( .A(n321), .Y(mem_wdata_D[114]) );
  CLKBUFX12 U62 ( .A(n320), .Y(mem_wdata_D[115]) );
  CLKBUFX12 U63 ( .A(n319), .Y(mem_wdata_D[116]) );
  CLKBUFX12 U64 ( .A(n318), .Y(mem_wdata_D[117]) );
  CLKBUFX12 U65 ( .A(n317), .Y(mem_wdata_D[118]) );
  CLKBUFX12 U66 ( .A(n316), .Y(mem_wdata_D[119]) );
  CLKBUFX12 U67 ( .A(n315), .Y(mem_wdata_D[120]) );
  BUFX20 U68 ( .A(n468), .Y(DCACHE_addr[4]) );
  INVXL U69 ( .A(n299), .Y(n2) );
  INVX12 U70 ( .A(n2), .Y(DCACHE_addr[3]) );
  BUFX20 U71 ( .A(n469), .Y(n299) );
  BUFX20 U72 ( .A(ICACHE_addr[2]), .Y(n295) );
  BUFX12 U73 ( .A(ICACHE_addr[3]), .Y(n296) );
  INVX4 U74 ( .A(n314), .Y(n4) );
  CLKINVX20 U75 ( .A(n4), .Y(mem_addr_D[4]) );
  BUFX20 U76 ( .A(n466), .Y(mem_wdata_I[83]) );
  BUFX20 U77 ( .A(n465), .Y(mem_wdata_I[84]) );
  BUFX20 U78 ( .A(n464), .Y(mem_wdata_I[85]) );
  BUFX20 U79 ( .A(n463), .Y(mem_wdata_I[86]) );
  BUFX20 U80 ( .A(n462), .Y(mem_wdata_I[87]) );
  INVX20 U81 ( .A(n11), .Y(mem_wdata_I[88]) );
  INVX20 U82 ( .A(n13), .Y(mem_wdata_I[89]) );
  INVX20 U83 ( .A(n15), .Y(mem_wdata_I[94]) );
  INVX20 U84 ( .A(n17), .Y(mem_wdata_I[96]) );
  INVX20 U85 ( .A(n19), .Y(mem_wdata_I[97]) );
  INVX20 U86 ( .A(n21), .Y(mem_wdata_I[98]) );
  INVX20 U87 ( .A(n23), .Y(mem_wdata_I[99]) );
  INVX20 U88 ( .A(n25), .Y(mem_wdata_I[100]) );
  INVX20 U89 ( .A(n27), .Y(mem_wdata_I[101]) );
  INVX20 U90 ( .A(n29), .Y(mem_wdata_I[102]) );
  INVX20 U91 ( .A(n31), .Y(mem_wdata_I[103]) );
  INVX20 U92 ( .A(n33), .Y(mem_wdata_I[104]) );
  INVX20 U93 ( .A(n35), .Y(mem_wdata_I[105]) );
  INVX4 U94 ( .A(n431), .Y(n37) );
  INVX20 U95 ( .A(n37), .Y(mem_addr_I[4]) );
  INVX20 U96 ( .A(n39), .Y(mem_wdata_I[106]) );
  INVX20 U97 ( .A(n41), .Y(mem_wdata_I[107]) );
  INVX20 U98 ( .A(n43), .Y(mem_wdata_I[108]) );
  INVX20 U99 ( .A(n45), .Y(mem_wdata_I[109]) );
  INVX20 U100 ( .A(n47), .Y(mem_wdata_I[110]) );
  INVX20 U101 ( .A(n49), .Y(mem_wdata_I[112]) );
  INVX20 U102 ( .A(n51), .Y(mem_wdata_I[113]) );
  INVX20 U103 ( .A(n53), .Y(mem_wdata_I[114]) );
  INVX20 U104 ( .A(n55), .Y(mem_wdata_I[115]) );
  INVX20 U105 ( .A(n57), .Y(mem_wdata_I[116]) );
  INVX20 U106 ( .A(n59), .Y(mem_wdata_I[117]) );
  INVX20 U107 ( .A(n61), .Y(mem_wdata_I[118]) );
  INVX20 U108 ( .A(n63), .Y(mem_wdata_I[119]) );
  INVX20 U109 ( .A(n65), .Y(mem_wdata_I[120]) );
  CLKINVX6 U110 ( .A(n467), .Y(n67) );
  INVX20 U111 ( .A(n67), .Y(mem_wdata_I[0]) );
  CLKINVX6 U112 ( .A(n434), .Y(n69) );
  INVX20 U113 ( .A(n69), .Y(mem_wdata_I[121]) );
  CLKINVX6 U114 ( .A(n433), .Y(n71) );
  INVX20 U115 ( .A(n71), .Y(mem_wdata_I[125]) );
  CLKINVX6 U116 ( .A(n432), .Y(n73) );
  INVX20 U117 ( .A(n73), .Y(mem_wdata_I[126]) );
  INVX4 U118 ( .A(n313), .Y(n75) );
  CLKINVX20 U119 ( .A(n75), .Y(mem_addr_D[5]) );
  INVX4 U120 ( .A(n312), .Y(n77) );
  CLKINVX20 U121 ( .A(n77), .Y(mem_addr_D[6]) );
  CLKBUFX20 U122 ( .A(n398), .Y(mem_wdata_D[37]) );
  INVX4 U123 ( .A(n427), .Y(n81) );
  INVX20 U124 ( .A(n81), .Y(mem_wdata_D[8]) );
  INVX4 U125 ( .A(n389), .Y(n83) );
  INVX20 U126 ( .A(n83), .Y(mem_wdata_D[46]) );
  INVX4 U127 ( .A(n426), .Y(n85) );
  INVX20 U128 ( .A(n85), .Y(mem_wdata_D[9]) );
  INVX4 U129 ( .A(n388), .Y(n87) );
  INVX20 U130 ( .A(n87), .Y(mem_wdata_D[47]) );
  INVX4 U131 ( .A(n425), .Y(n89) );
  INVX20 U132 ( .A(n89), .Y(mem_wdata_D[10]) );
  INVX4 U133 ( .A(n387), .Y(n91) );
  INVX20 U134 ( .A(n91), .Y(mem_wdata_D[48]) );
  INVX4 U135 ( .A(n424), .Y(n93) );
  INVX20 U136 ( .A(n93), .Y(mem_wdata_D[11]) );
  INVX4 U137 ( .A(n386), .Y(n95) );
  INVX20 U138 ( .A(n95), .Y(mem_wdata_D[49]) );
  INVX4 U139 ( .A(n423), .Y(n97) );
  INVX20 U140 ( .A(n97), .Y(mem_wdata_D[12]) );
  INVX4 U141 ( .A(n385), .Y(n99) );
  INVX20 U142 ( .A(n99), .Y(mem_wdata_D[50]) );
  INVX4 U143 ( .A(n422), .Y(n101) );
  INVX20 U144 ( .A(n101), .Y(mem_wdata_D[13]) );
  INVX4 U145 ( .A(n384), .Y(n103) );
  INVX20 U146 ( .A(n103), .Y(mem_wdata_D[51]) );
  INVX4 U147 ( .A(n421), .Y(n105) );
  INVX20 U148 ( .A(n105), .Y(mem_wdata_D[14]) );
  INVX4 U149 ( .A(n383), .Y(n107) );
  INVX20 U150 ( .A(n107), .Y(mem_wdata_D[52]) );
  INVX4 U151 ( .A(n420), .Y(n109) );
  INVX20 U152 ( .A(n109), .Y(mem_wdata_D[15]) );
  INVX4 U153 ( .A(n382), .Y(n111) );
  INVX20 U154 ( .A(n111), .Y(mem_wdata_D[53]) );
  INVX4 U155 ( .A(n419), .Y(n113) );
  INVX20 U156 ( .A(n113), .Y(mem_wdata_D[16]) );
  INVX4 U157 ( .A(n381), .Y(n115) );
  INVX20 U158 ( .A(n115), .Y(mem_wdata_D[54]) );
  INVX4 U159 ( .A(n418), .Y(n117) );
  INVX20 U160 ( .A(n117), .Y(mem_wdata_D[17]) );
  INVX4 U161 ( .A(n380), .Y(n119) );
  INVX20 U162 ( .A(n119), .Y(mem_wdata_D[55]) );
  INVX4 U163 ( .A(n417), .Y(n121) );
  INVX20 U164 ( .A(n121), .Y(mem_wdata_D[18]) );
  INVX4 U165 ( .A(n379), .Y(n123) );
  INVX20 U166 ( .A(n123), .Y(mem_wdata_D[56]) );
  INVX4 U167 ( .A(n416), .Y(n125) );
  INVX20 U168 ( .A(n125), .Y(mem_wdata_D[19]) );
  INVX4 U169 ( .A(n378), .Y(n127) );
  INVX20 U170 ( .A(n127), .Y(mem_wdata_D[57]) );
  INVX4 U171 ( .A(n415), .Y(n129) );
  INVX20 U172 ( .A(n129), .Y(mem_wdata_D[20]) );
  INVX4 U173 ( .A(n377), .Y(n131) );
  INVX20 U174 ( .A(n131), .Y(mem_wdata_D[58]) );
  INVX4 U175 ( .A(n414), .Y(n133) );
  INVX20 U176 ( .A(n133), .Y(mem_wdata_D[21]) );
  INVX4 U177 ( .A(n376), .Y(n135) );
  INVX20 U178 ( .A(n135), .Y(mem_wdata_D[59]) );
  INVX4 U179 ( .A(n413), .Y(n137) );
  INVX20 U180 ( .A(n137), .Y(mem_wdata_D[22]) );
  INVX4 U181 ( .A(n375), .Y(n139) );
  INVX20 U182 ( .A(n139), .Y(mem_wdata_D[60]) );
  INVX4 U183 ( .A(n412), .Y(n141) );
  INVX20 U184 ( .A(n141), .Y(mem_wdata_D[23]) );
  INVX4 U185 ( .A(n374), .Y(n143) );
  INVX20 U186 ( .A(n143), .Y(mem_wdata_D[61]) );
  INVX4 U187 ( .A(n411), .Y(n145) );
  INVX20 U188 ( .A(n145), .Y(mem_wdata_D[24]) );
  INVX4 U189 ( .A(n373), .Y(n147) );
  INVX20 U190 ( .A(n147), .Y(mem_wdata_D[62]) );
  INVX4 U191 ( .A(n410), .Y(n149) );
  INVX20 U192 ( .A(n149), .Y(mem_wdata_D[25]) );
  INVX4 U193 ( .A(n372), .Y(n151) );
  INVX20 U194 ( .A(n151), .Y(mem_wdata_D[63]) );
  INVX4 U195 ( .A(n409), .Y(n154) );
  INVX20 U196 ( .A(n154), .Y(mem_wdata_D[26]) );
  INVX4 U197 ( .A(n371), .Y(n156) );
  INVX20 U198 ( .A(n156), .Y(mem_wdata_D[64]) );
  INVX20 U199 ( .A(n158), .Y(mem_wdata_D[84]) );
  INVX4 U200 ( .A(n408), .Y(n160) );
  INVX20 U201 ( .A(n160), .Y(mem_wdata_D[27]) );
  INVX4 U202 ( .A(n370), .Y(n162) );
  INVX20 U203 ( .A(n162), .Y(mem_wdata_D[65]) );
  INVX20 U204 ( .A(n164), .Y(mem_wdata_D[85]) );
  INVX4 U205 ( .A(n407), .Y(n166) );
  INVX20 U206 ( .A(n166), .Y(mem_wdata_D[28]) );
  INVX4 U207 ( .A(n369), .Y(n168) );
  INVX20 U208 ( .A(n168), .Y(mem_wdata_D[66]) );
  INVX20 U209 ( .A(n170), .Y(mem_wdata_D[86]) );
  INVX4 U210 ( .A(n406), .Y(n172) );
  INVX20 U211 ( .A(n172), .Y(mem_wdata_D[29]) );
  INVX4 U212 ( .A(n368), .Y(n174) );
  INVX20 U213 ( .A(n174), .Y(mem_wdata_D[67]) );
  INVX20 U214 ( .A(n176), .Y(mem_wdata_D[87]) );
  INVX4 U215 ( .A(n405), .Y(n178) );
  INVX20 U216 ( .A(n178), .Y(mem_wdata_D[30]) );
  INVX4 U217 ( .A(n367), .Y(n180) );
  INVX20 U218 ( .A(n180), .Y(mem_wdata_D[68]) );
  INVX20 U219 ( .A(n182), .Y(mem_wdata_D[88]) );
  INVX4 U220 ( .A(n404), .Y(n184) );
  INVX20 U221 ( .A(n184), .Y(mem_wdata_D[31]) );
  INVX4 U222 ( .A(n366), .Y(n186) );
  INVX20 U223 ( .A(n186), .Y(mem_wdata_D[69]) );
  INVX20 U224 ( .A(n188), .Y(mem_wdata_D[89]) );
  INVX4 U225 ( .A(n403), .Y(n190) );
  INVX20 U226 ( .A(n190), .Y(mem_wdata_D[32]) );
  INVX4 U227 ( .A(n365), .Y(n192) );
  INVX20 U228 ( .A(n192), .Y(mem_wdata_D[70]) );
  INVX20 U229 ( .A(n194), .Y(mem_wdata_D[90]) );
  INVX4 U230 ( .A(n402), .Y(n196) );
  INVX20 U231 ( .A(n196), .Y(mem_wdata_D[33]) );
  INVX4 U232 ( .A(n364), .Y(n198) );
  INVX20 U233 ( .A(n198), .Y(mem_wdata_D[71]) );
  INVX20 U234 ( .A(n200), .Y(mem_wdata_D[91]) );
  INVX4 U235 ( .A(n401), .Y(n202) );
  INVX20 U236 ( .A(n202), .Y(mem_wdata_D[34]) );
  INVX4 U237 ( .A(n363), .Y(n204) );
  INVX20 U238 ( .A(n204), .Y(mem_wdata_D[72]) );
  INVX20 U239 ( .A(n206), .Y(mem_wdata_D[92]) );
  INVX4 U240 ( .A(n400), .Y(n208) );
  INVX20 U241 ( .A(n208), .Y(mem_wdata_D[35]) );
  INVX4 U242 ( .A(n362), .Y(n210) );
  INVX20 U243 ( .A(n210), .Y(mem_wdata_D[73]) );
  INVX20 U244 ( .A(n212), .Y(mem_wdata_D[93]) );
  INVX4 U245 ( .A(n399), .Y(n214) );
  INVX20 U246 ( .A(n214), .Y(mem_wdata_D[36]) );
  INVX4 U247 ( .A(n361), .Y(n216) );
  INVX20 U248 ( .A(n216), .Y(mem_wdata_D[74]) );
  INVX20 U249 ( .A(n218), .Y(mem_wdata_D[94]) );
  INVX4 U250 ( .A(n397), .Y(n220) );
  INVX20 U251 ( .A(n220), .Y(mem_wdata_D[38]) );
  INVX4 U252 ( .A(n360), .Y(n222) );
  INVX20 U253 ( .A(n222), .Y(mem_wdata_D[75]) );
  INVX20 U254 ( .A(n224), .Y(mem_wdata_D[95]) );
  BUFX20 U255 ( .A(n396), .Y(mem_wdata_D[39]) );
  BUFX20 U256 ( .A(n359), .Y(mem_wdata_D[76]) );
  INVX20 U257 ( .A(n228), .Y(mem_wdata_D[96]) );
  BUFX20 U258 ( .A(n395), .Y(mem_wdata_D[40]) );
  BUFX20 U259 ( .A(n358), .Y(mem_wdata_D[77]) );
  INVX20 U260 ( .A(n232), .Y(mem_wdata_D[97]) );
  BUFX20 U261 ( .A(n394), .Y(mem_wdata_D[41]) );
  BUFX20 U262 ( .A(n357), .Y(mem_wdata_D[78]) );
  INVX20 U263 ( .A(n236), .Y(mem_wdata_D[98]) );
  BUFX20 U264 ( .A(n393), .Y(mem_wdata_D[42]) );
  BUFX20 U265 ( .A(n356), .Y(mem_wdata_D[79]) );
  INVX20 U266 ( .A(n240), .Y(mem_wdata_D[99]) );
  BUFX20 U267 ( .A(n392), .Y(mem_wdata_D[43]) );
  BUFX20 U268 ( .A(n355), .Y(mem_wdata_D[80]) );
  INVX20 U269 ( .A(n244), .Y(mem_wdata_D[100]) );
  BUFX20 U270 ( .A(n391), .Y(mem_wdata_D[44]) );
  BUFX20 U271 ( .A(n354), .Y(mem_wdata_D[81]) );
  INVX20 U272 ( .A(n248), .Y(mem_wdata_D[101]) );
  BUFX20 U273 ( .A(n390), .Y(mem_wdata_D[45]) );
  BUFX20 U274 ( .A(n353), .Y(mem_wdata_D[82]) );
  INVX20 U275 ( .A(n252), .Y(mem_wdata_D[102]) );
  INVX20 U276 ( .A(n254), .Y(mem_wdata_D[103]) );
  INVX20 U277 ( .A(n256), .Y(mem_wdata_D[104]) );
  INVX20 U278 ( .A(n258), .Y(mem_wdata_D[105]) );
  INVX20 U279 ( .A(n260), .Y(mem_wdata_D[106]) );
  INVX20 U280 ( .A(n262), .Y(mem_wdata_D[107]) );
  CLKBUFX20 U281 ( .A(n470), .Y(DCACHE_addr[2]) );
  INVXL U282 ( .A(n301), .Y(n302) );
  CLKINVX3 U283 ( .A(n311), .Y(n277) );
  CLKINVX3 U284 ( .A(n307), .Y(n285) );
  CLKINVX3 U285 ( .A(n310), .Y(n279) );
  CLKINVX3 U286 ( .A(n309), .Y(n281) );
  CLKINVX3 U287 ( .A(n306), .Y(n287) );
  BUFX8 U288 ( .A(ICACHE_addr[4]), .Y(n297) );
  BUFX8 U289 ( .A(rst_n), .Y(n301) );
  BUFX12 U290 ( .A(n304), .Y(mem_write_D) );
  BUFX12 U291 ( .A(n430), .Y(mem_write_I) );
  BUFX12 U292 ( .A(n303), .Y(mem_read_D) );
  BUFX12 U293 ( .A(n429), .Y(mem_read_I) );
  INVX12 U294 ( .A(n285), .Y(mem_addr_D[14]) );
  INVX12 U295 ( .A(n279), .Y(mem_addr_D[9]) );
  INVX12 U296 ( .A(n281), .Y(mem_addr_D[11]) );
  INVX12 U297 ( .A(n287), .Y(mem_addr_D[16]) );
  INVX12 U298 ( .A(n283), .Y(mem_addr_D[12]) );
  CLKINVX1 U299 ( .A(n308), .Y(n283) );
  INVX12 U300 ( .A(n289), .Y(mem_addr_D[17]) );
  CLKINVX1 U301 ( .A(n305), .Y(n289) );
  INVX12 U302 ( .A(n277), .Y(mem_addr_D[8]) );
endmodule

